*****************************************************************************
* CDL Netlist:
* Cell Name: ram
* Netlisted on: Dec 21 13:51:54 2006
*****************************************************************************


*****************************************************************************
* Global Net Declarations
*****************************************************************************
*.GLOBAL gnd vdd

.OPTION SCALE=1E-6

*****************************************************************************
* PIN Control Statement
*****************************************************************************
*.PIN gnd vdd


*****************************************************************************
* BIPOLAR Declarations
*****************************************************************************


*.LDD

*****************************************************************************
* Parameter Statement
*****************************************************************************
.PARAM


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*         0                                                                    *
* Block: colmux                                                               *
* Last Time Saved: Dec 12 11:40:47 2006                                       *
*******************************************************************************
.subckt colmux DB DB_ bl<15> bl<14> bl<13> bl<12> bl<11> bl<10> bl<9> bl<8>
+bl<7> bl<6> bl<5> bl<4> bl<3> bl<2> bl<1> bl<0> bl_<15> bl_<14> bl_<13>
+bl_<12> bl_<11> bl_<10> bl_<9> bl_<8> bl_<7> bl_<6> bl_<5> bl_<4> bl_<3>
+bl_<2> bl_<1> bl_<0> ysel<15> ysel<14> ysel<13> ysel<12> ysel<11> ysel<10>
+ysel<9> ysel<8> ysel<7> ysel<6> ysel<5> ysel<4> ysel<3> ysel<2> ysel<1>
+ysel<0>
*.NOPIN gnd vdd
MN0_15 bl<15> ysel<15> DB gnd n18ll w=1.5 l=0.18
MN0_14 bl<14> ysel<14> DB gnd n18ll w=1.5 l=0.18
MN0_13 bl<13> ysel<13> DB gnd n18ll w=1.5 l=0.18
MN0_12 bl<12> ysel<12> DB gnd n18ll w=1.5 l=0.18
MN0_11 bl<11> ysel<11> DB gnd n18ll w=1.5 l=0.18
MN0_10 bl<10> ysel<10> DB gnd n18ll w=1.5 l=0.18
MN0_9 bl<9> ysel<9> DB gnd n18ll w=1.5 l=0.18
MN0_8 bl<8> ysel<8> DB gnd n18ll w=1.5 l=0.18
MN0_7 bl<7> ysel<7> DB gnd n18ll w=1.5 l=0.18
MN0_6 bl<6> ysel<6> DB gnd n18ll w=1.5 l=0.18
MN0_5 bl<5> ysel<5> DB gnd n18ll w=1.5 l=0.18
MN0_4 bl<4> ysel<4> DB gnd n18ll w=1.5 l=0.18
MN0_3 bl<3> ysel<3> DB gnd n18ll w=1.5 l=0.18
MN0_2 bl<2> ysel<2> DB gnd n18ll w=1.5 l=0.18
MN0_1 bl<1> ysel<1> DB gnd n18ll w=1.5 l=0.18
MN0_0 bl<0> ysel<0> DB gnd n18ll w=1.5 l=0.18
MN1_15 bl_<15> ysel<15> DB_ gnd n18ll w=1.5 l=0.18
MN1_14 bl_<14> ysel<14> DB_ gnd n18ll w=1.5 l=0.18
MN1_13 bl_<13> ysel<13> DB_ gnd n18ll w=1.5 l=0.18
MN1_12 bl_<12> ysel<12> DB_ gnd n18ll w=1.5 l=0.18
MN1_11 bl_<11> ysel<11> DB_ gnd n18ll w=1.5 l=0.18
MN1_10 bl_<10> ysel<10> DB_ gnd n18ll w=1.5 l=0.18
MN1_9 bl_<9> ysel<9> DB_ gnd n18ll w=1.5 l=0.18
MN1_8 bl_<8> ysel<8> DB_ gnd n18ll w=1.5 l=0.18
MN1_7 bl_<7> ysel<7> DB_ gnd n18ll w=1.5 l=0.18
MN1_6 bl_<6> ysel<6> DB_ gnd n18ll w=1.5 l=0.18
MN1_5 bl_<5> ysel<5> DB_ gnd n18ll w=1.5 l=0.18
MN1_4 bl_<4> ysel<4> DB_ gnd n18ll w=1.5 l=0.18
MN1_3 bl_<3> ysel<3> DB_ gnd n18ll w=1.5 l=0.18
MN1_2 bl_<2> ysel<2> DB_ gnd n18ll w=1.5 l=0.18
MN1_1 bl_<1> ysel<1> DB_ gnd n18ll w=1.5 l=0.18
MN1_0 bl_<0> ysel<0> DB_ gnd n18ll w=1.5 l=0.18
.ends colmux


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                  1                                                           *
* Block: inv                                                                  *
* Last Time Saved: Aug 18 08:37:34 2004                                       *
*******************************************************************************
.subckt inv Y A ln=0.54 wn=2.7 lp=0.54 wp=5.4
MP0 Y A vdd vdd p18ll w=wp l=lp
MN0 Y A gnd gnd n18ll w=wn l=ln
.ends inv


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                       2                                                      *
* Block: nand2                                                                *
* Last Time Saved: Aug 18 08:34:53 2004                                       *
*******************************************************************************
.subckt nand2 Y A B lp=0.54 wp=5.4 ln=0.54 wn=2.7
MN0 net13 B gnd gnd n18ll w=wn l=ln
MN1 Y A net13 gnd n18ll w=wn l=ln
MP0 Y B vdd vdd p18ll w=wp l=lp
MP1 Y A vdd vdd p18ll w=wp l=lp
.ends nand2


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                            3                                                 *
* Block: preck_gen                                                            *
* Last Time Saved: Dec 12 11:40:19 2006                                       *
*******************************************************************************
.subckt preck_gen PRECK sck_bar
XI3 net5 net17 inv ln=0.18 wn=0.4 lp=0.18 wp=1
XI4 PRECK net5 inv ln=0.18 wn=1.5 lp=0.18 wp=4
XI93 net018 sck_bar inv ln=1.0 wn=0.5 lp=1.0 wp=1.25
XI92 net012 net018 inv ln=1.0 wn=0.5 lp=1.0 wp=1.25
XI90 net7 net014 inv ln=1.0 wn=0.5 lp=1.0 wp=1.25
XI91 net014 net012 inv ln=1.0 wn=0.5 lp=1.0 wp=1.25
XI2 net17 sck_bar net7 nand2 lp=0.18 wp=0.6 ln=0.18 wn=0.4
.ends preck_gen


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                        4                                                     *
* Block: rdwr_drive                                                           *
* Last Time Saved: Dec 12 11:40:57 2006                                       *
*******************************************************************************
.subckt rdwr_drive dout BL BL_ preck rd_en wr_en wrdata wrdata_
MN8 vdd net8 BL_ vdd p18ll w=6 l=0.18
MP0 BL net23 vdd vdd p18ll w=6 l=0.18
MP4 BL_ preck vdd vdd p18ll w=2.0 l=0.18
MP1 BL preck vdd vdd p18ll w=2.0 l=0.18
MP5 BL_ preck BL vdd p18ll w=0.5 l=0.18
MN7 vdd net090 dout vdd p18ll w=6 l=0.18
XI53 net063 rd_en data_out_ nand2 lp=0.18 wp=1 ln=0.18 wn=0.8
XI34 net26 wrdata wr_en nand2 lp=0.18 wp=1 ln=0.18 wn=0.8
XI33 net8 wr_en wrdata_ nand2 lp=0.18 wp=1 ln=0.18 wn=0.8
XI32 net20 wr_en wrdata_ nand2 lp=0.18 wp=1 ln=0.18 wn=0.8
XI18 net23 wrdata wr_en nand2 lp=0.18 wp=1 ln=0.18 wn=0.8
XI52 net090 data_out rd_en nand2 lp=0.18 wp=1 ln=0.18 wn=0.8
MP3 gnd net089 BL_ gnd n18ll w=2 l=0.18
MN5 BL net0103 gnd gnd n18ll w=2 l=0.18
MN4 data_out_ net32 gnd gnd n18ll w=1 l=0.18
MN0 data_out net52 gnd gnd n18ll w=1 l=0.18
MN9 gnd net0112 dout gnd n18ll w=2 l=0.18
XI49 net0112 net063 inv ln=0.18 wn=0.3 lp=0.18 wp=0.6
XI46 net089 net26 inv ln=0.18 wn=0.3 lp=0.18 wp=0.6
XI42 data_out_ data_out inv ln=0.18 wn=0.3 lp=0.18 wp=0.6
XI45 net0103 net20 inv ln=0.18 wn=0.3 lp=0.18 wp=0.6
XI41 net32 BL_ inv ln=0.18 wn=0.4 lp=0.18 wp=1
XI6 net52 BL inv ln=0.18 wn=0.4 lp=0.18 wp=1
XI43 data_out data_out_ inv ln=0.18 wn=0.3 lp=0.18 wp=0.6
.ends rdwr_drive


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                          5                                                   *
* Block: precharge                                                            *
* Last Time Saved: Dec 12 11:40:27 2006                                       *
*******************************************************************************
.subckt precharge bl bl_ precharge
*.NOPIN gnd
MP2 bl_ precharge bl vdd p18ll w=0.5 l=0.18
MP1 bl_ precharge vdd vdd p18ll w=2.0 l=0.18
MP0 bl precharge vdd vdd p18ll w=2.0 l=0.18
.ends precharge


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                            6                                                 *
* Block: memcell                                                              *
* Last Time Saved: Dec 12 09:51:41 2006                                       *
*******************************************************************************
.subckt memcell BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7>
+BL<6> BL<5> BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12>
+BL_<11> BL_<10> BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1>
+BL_<0> WL
MN0_15 BL<15> WL d<15> gnd n18ll w=0.24 l=0.22
MN0_14 BL<14> WL d<14> gnd n18ll w=0.24 l=0.22
MN0_13 BL<13> WL d<13> gnd n18ll w=0.24 l=0.22
MN0_12 BL<12> WL d<12> gnd n18ll w=0.24 l=0.22
MN0_11 BL<11> WL d<11> gnd n18ll w=0.24 l=0.22
MN0_10 BL<10> WL d<10> gnd n18ll w=0.24 l=0.22
MN0_9 BL<9> WL d<9> gnd n18ll w=0.24 l=0.22
MN0_8 BL<8> WL d<8> gnd n18ll w=0.24 l=0.22
MN0_7 BL<7> WL d<7> gnd n18ll w=0.24 l=0.22
MN0_6 BL<6> WL d<6> gnd n18ll w=0.24 l=0.22
MN0_5 BL<5> WL d<5> gnd n18ll w=0.24 l=0.22
MN0_4 BL<4> WL d<4> gnd n18ll w=0.24 l=0.22
MN0_3 BL<3> WL d<3> gnd n18ll w=0.24 l=0.22
MN0_2 BL<2> WL d<2> gnd n18ll w=0.24 l=0.22
MN0_1 BL<1> WL d<1> gnd n18ll w=0.24 l=0.22
MN0_0 BL<0> WL d<0> gnd n18ll w=0.24 l=0.22
MN1_15 d_<15> WL BL_<15> gnd n18ll w=0.24 l=0.22
MN1_14 d_<14> WL BL_<14> gnd n18ll w=0.24 l=0.22
MN1_13 d_<13> WL BL_<13> gnd n18ll w=0.24 l=0.22
MN1_12 d_<12> WL BL_<12> gnd n18ll w=0.24 l=0.22
MN1_11 d_<11> WL BL_<11> gnd n18ll w=0.24 l=0.22
MN1_10 d_<10> WL BL_<10> gnd n18ll w=0.24 l=0.22
MN1_9 d_<9> WL BL_<9> gnd n18ll w=0.24 l=0.22
MN1_8 d_<8> WL BL_<8> gnd n18ll w=0.24 l=0.22
MN1_7 d_<7> WL BL_<7> gnd n18ll w=0.24 l=0.22
MN1_6 d_<6> WL BL_<6> gnd n18ll w=0.24 l=0.22
MN1_5 d_<5> WL BL_<5> gnd n18ll w=0.24 l=0.22
MN1_4 d_<4> WL BL_<4> gnd n18ll w=0.24 l=0.22
MN1_3 d_<3> WL BL_<3> gnd n18ll w=0.24 l=0.22
MN1_2 d_<2> WL BL_<2> gnd n18ll w=0.24 l=0.22
MN1_1 d_<1> WL BL_<1> gnd n18ll w=0.24 l=0.22
MN1_0 d_<0> WL BL_<0> gnd n18ll w=0.24 l=0.22
XI0_15 d<15> d_<15> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI0_14 d<14> d_<14> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI0_13 d<13> d_<13> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI0_12 d<12> d_<12> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI0_11 d<11> d_<11> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI0_10 d<10> d_<10> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI0_9 d<9> d_<9> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI0_8 d<8> d_<8> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI0_7 d<7> d_<7> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI0_6 d<6> d_<6> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI0_5 d<5> d_<5> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI0_4 d<4> d_<4> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI0_3 d<3> d_<3> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI0_2 d<2> d_<2> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI0_1 d<1> d_<1> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI0_0 d<0> d_<0> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI1_15 d_<15> d<15> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI1_14 d_<14> d<14> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI1_13 d_<13> d<13> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI1_12 d_<12> d<12> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI1_11 d_<11> d<11> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI1_10 d_<10> d<10> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI1_9 d_<9> d<9> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI1_8 d_<8> d<8> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI1_7 d_<7> d<7> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI1_6 d_<6> d<6> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI1_5 d_<5> d<5> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI1_4 d_<4> d<4> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI1_3 d_<3> d<3> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI1_2 d_<2> d<2> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI1_1 d_<1> d<1> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
XI1_0 d_<0> d<0> inv ln=0.18 wn=0.35 lp=0.18 wp=0.20
.ends memcell


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                             7                                                *
* Block: memarray_64x16                                                       *
* Last Time Saved: Dec 12 11:40:37 2006                                       *
*******************************************************************************
.subckt memarray_64x16 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8>
+BL<7> BL<6> BL<5> BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13>
+BL_<12> BL_<11> BL_<10> BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3>
+BL_<2> BL_<1> BL_<0> WL<63> WL<62> WL<61> WL<60> WL<59> WL<58> WL<57> WL<56>
+WL<55> WL<54> WL<53> WL<52> WL<51> WL<50> WL<49> WL<48> WL<47> WL<46> WL<45>
+WL<44> WL<43> WL<42> WL<41> WL<40> WL<39> WL<38> WL<37> WL<36> WL<35> WL<34>
+WL<33> WL<32> WL<31> WL<30> WL<29> WL<28> WL<27> WL<26> WL<25> WL<24> WL<23>
+WL<22> WL<21> WL<20> WL<19> WL<18> WL<17> WL<16> WL<15> WL<14> WL<13> WL<12>
+WL<11> WL<10> WL<9> WL<8> WL<7> WL<6> WL<5> WL<4> WL<3> WL<2> WL<1> WL<0>
MN0_15 gnd gnd BL<15> gnd n18ll w=0.24 l=0.22 m=2
MN0_14 gnd gnd BL<14> gnd n18ll w=0.24 l=0.22 m=2
MN0_13 gnd gnd BL<13> gnd n18ll w=0.24 l=0.22 m=2
MN0_12 gnd gnd BL<12> gnd n18ll w=0.24 l=0.22 m=2
MN0_11 gnd gnd BL<11> gnd n18ll w=0.24 l=0.22 m=2
MN0_10 gnd gnd BL<10> gnd n18ll w=0.24 l=0.22 m=2
MN0_9 gnd gnd BL<9> gnd n18ll w=0.24 l=0.22 m=2
MN0_8 gnd gnd BL<8> gnd n18ll w=0.24 l=0.22 m=2
MN0_7 gnd gnd BL<7> gnd n18ll w=0.24 l=0.22 m=2
MN0_6 gnd gnd BL<6> gnd n18ll w=0.24 l=0.22 m=2
MN0_5 gnd gnd BL<5> gnd n18ll w=0.24 l=0.22 m=2
MN0_4 gnd gnd BL<4> gnd n18ll w=0.24 l=0.22 m=2
MN0_3 gnd gnd BL<3> gnd n18ll w=0.24 l=0.22 m=2
MN0_2 gnd gnd BL<2> gnd n18ll w=0.24 l=0.22 m=2
MN0_1 gnd gnd BL<1> gnd n18ll w=0.24 l=0.22 m=2
MN0_0 gnd gnd BL<0> gnd n18ll w=0.24 l=0.22 m=2
MN1_15 gnd gnd BL_<15> gnd n18ll w=0.24 l=0.22 m=2
MN1_14 gnd gnd BL_<14> gnd n18ll w=0.24 l=0.22 m=2
MN1_13 gnd gnd BL_<13> gnd n18ll w=0.24 l=0.22 m=2
MN1_12 gnd gnd BL_<12> gnd n18ll w=0.24 l=0.22 m=2
MN1_11 gnd gnd BL_<11> gnd n18ll w=0.24 l=0.22 m=2
MN1_10 gnd gnd BL_<10> gnd n18ll w=0.24 l=0.22 m=2
MN1_9 gnd gnd BL_<9> gnd n18ll w=0.24 l=0.22 m=2
MN1_8 gnd gnd BL_<8> gnd n18ll w=0.24 l=0.22 m=2
MN1_7 gnd gnd BL_<7> gnd n18ll w=0.24 l=0.22 m=2
MN1_6 gnd gnd BL_<6> gnd n18ll w=0.24 l=0.22 m=2
MN1_5 gnd gnd BL_<5> gnd n18ll w=0.24 l=0.22 m=2
MN1_4 gnd gnd BL_<4> gnd n18ll w=0.24 l=0.22 m=2
MN1_3 gnd gnd BL_<3> gnd n18ll w=0.24 l=0.22 m=2
MN1_2 gnd gnd BL_<2> gnd n18ll w=0.24 l=0.22 m=2
MN1_1 gnd gnd BL_<1> gnd n18ll w=0.24 l=0.22 m=2
MN1_0 gnd gnd BL_<0> gnd n18ll w=0.24 l=0.22 m=2
XI0_63 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<63>
+memcell
XI0_62 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<62>
+memcell
XI0_61 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<61>
+memcell
XI0_60 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<60>
+memcell
XI0_59 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<59>
+memcell
XI0_58 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<58>
+memcell
XI0_57 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<57>
+memcell
XI0_56 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<56>
+memcell
XI0_55 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<55>
+memcell
XI0_54 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<54>
+memcell
XI0_53 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<53>
+memcell
XI0_52 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<52>
+memcell
XI0_51 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<51>
+memcell
XI0_50 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<50>
+memcell
XI0_49 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<49>
+memcell
XI0_48 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<48>
+memcell
XI0_47 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<47>
+memcell
XI0_46 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<46>
+memcell
XI0_45 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<45>
+memcell
XI0_44 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<44>
+memcell
XI0_43 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<43>
+memcell
XI0_42 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<42>
+memcell
XI0_41 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<41>
+memcell
XI0_40 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<40>
+memcell
XI0_39 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<39>
+memcell
XI0_38 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<38>
+memcell
XI0_37 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<37>
+memcell
XI0_36 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<36>
+memcell
XI0_35 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<35>
+memcell
XI0_34 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<34>
+memcell
XI0_33 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<33>
+memcell
XI0_32 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<32>
+memcell
XI0_31 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<31>
+memcell
XI0_30 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<30>
+memcell
XI0_29 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<29>
+memcell
XI0_28 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<28>
+memcell
XI0_27 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<27>
+memcell
XI0_26 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<26>
+memcell
XI0_25 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<25>
+memcell
XI0_24 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<24>
+memcell
XI0_23 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<23>
+memcell
XI0_22 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<22>
+memcell
XI0_21 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<21>
+memcell
XI0_20 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<20>
+memcell
XI0_19 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<19>
+memcell
XI0_18 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<18>
+memcell
XI0_17 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<17>
+memcell
XI0_16 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<16>
+memcell
XI0_15 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<15>
+memcell
XI0_14 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<14>
+memcell
XI0_13 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<13>
+memcell
XI0_12 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<12>
+memcell
XI0_11 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<11>
+memcell
XI0_10 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<10>
+memcell
XI0_9 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<9>
+memcell
XI0_8 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<8>
+memcell
XI0_7 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<7>
+memcell
XI0_6 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<6>
+memcell
XI0_5 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<5>
+memcell
XI0_4 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<4>
+memcell
XI0_3 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<3>
+memcell
XI0_2 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<2>
+memcell
XI0_1 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<1>
+memcell
XI0_0 BL<15> BL<14> BL<13> BL<12> BL<11> BL<10> BL<9> BL<8> BL<7> BL<6> BL<5>
+BL<4> BL<3> BL<2> BL<1> BL<0> BL_<15> BL_<14> BL_<13> BL_<12> BL_<11> BL_<10>
+BL_<9> BL_<8> BL_<7> BL_<6> BL_<5> BL_<4> BL_<3> BL_<2> BL_<1> BL_<0> WL<0>
+memcell
.ends memarray_64x16


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                          8                                                   *
* Block: memblock                                                             *
* Last Time Saved: Dec 12 11:40:10 2006                                       *
*******************************************************************************
.subckt memblock dout rd_en sck_bar wr_en wrdata wrdata_ xsel<63> xsel<62>
+xsel<61> xsel<60> xsel<59> xsel<58> xsel<57> xsel<56> xsel<55> xsel<54>
+xsel<53> xsel<52> xsel<51> xsel<50> xsel<49> xsel<48> xsel<47> xsel<46>
+xsel<45> xsel<44> xsel<43> xsel<42> xsel<41> xsel<40> xsel<39> xsel<38>
+xsel<37> xsel<36> xsel<35> xsel<34> xsel<33> xsel<32> xsel<31> xsel<30>
+xsel<29> xsel<28> xsel<27> xsel<26> xsel<25> xsel<24> xsel<23> xsel<22>
+xsel<21> xsel<20> xsel<19> xsel<18> xsel<17> xsel<16> xsel<15> xsel<14>
+xsel<13> xsel<12> xsel<11> xsel<10> xsel<9> xsel<8> xsel<7> xsel<6> xsel<5>
+xsel<4> xsel<3> xsel<2> xsel<1> xsel<0> ysel<15> ysel<14> ysel<13> ysel<12>
+ysel<11> ysel<10> ysel<9> ysel<8> ysel<7> ysel<6> ysel<5> ysel<4> ysel<3>
+ysel<2> ysel<1> ysel<0>
XI2 net9 net12 net21<0> net21<1> net21<2> net21<3> net21<4> net21<5> net21<6>
+net21<7> net21<8> net21<9> net21<10> net21<11> net21<12> net21<13> net21<14>
+net21<15> net20<0> net20<1> net20<2> net20<3> net20<4> net20<5> net20<6>
+net20<7> net20<8> net20<9> net20<10> net20<11> net20<12> net20<13> net20<14>
+net20<15> ysel<15> ysel<14> ysel<13> ysel<12> ysel<11> ysel<10> ysel<9>
+ysel<8> ysel<7> ysel<6> ysel<5> ysel<4> ysel<3> ysel<2> ysel<1> ysel<0> colmux
XI3 preck sck_bar preck_gen
XI4 dout net9 net12 preck rd_en wr_en wrdata wrdata_ rdwr_drive
XI1_15 net21<0> net20<0> preck precharge
XI1_14 net21<1> net20<1> preck precharge
XI1_13 net21<2> net20<2> preck precharge
XI1_12 net21<3> net20<3> preck precharge
XI1_11 net21<4> net20<4> preck precharge
XI1_10 net21<5> net20<5> preck precharge
XI1_9 net21<6> net20<6> preck precharge
XI1_8 net21<7> net20<7> preck precharge
XI1_7 net21<8> net20<8> preck precharge
XI1_6 net21<9> net20<9> preck precharge
XI1_5 net21<10> net20<10> preck precharge
XI1_4 net21<11> net20<11> preck precharge
XI1_3 net21<12> net20<12> preck precharge
XI1_2 net21<13> net20<13> preck precharge
XI1_1 net21<14> net20<14> preck precharge
XI1_0 net21<15> net20<15> preck precharge
XI0 net21<0> net21<1> net21<2> net21<3> net21<4> net21<5> net21<6> net21<7>
+net21<8> net21<9> net21<10> net21<11> net21<12> net21<13> net21<14> net21<15>
+net20<0> net20<1> net20<2> net20<3> net20<4> net20<5> net20<6> net20<7>
+net20<8> net20<9> net20<10> net20<11> net20<12> net20<13> net20<14> net20<15>
+xsel<63> xsel<62> xsel<61> xsel<60> xsel<59> xsel<58> xsel<57> xsel<56>
+xsel<55> xsel<54> xsel<53> xsel<52> xsel<51> xsel<50> xsel<49> xsel<48>
+xsel<47> xsel<46> xsel<45> xsel<44> xsel<43> xsel<42> xsel<41> xsel<40>
+xsel<39> xsel<38> xsel<37> xsel<36> xsel<35> xsel<34> xsel<33> xsel<32>
+xsel<31> xsel<30> xsel<29> xsel<28> xsel<27> xsel<26> xsel<25> xsel<24>
+xsel<23> xsel<22> xsel<21> xsel<20> xsel<19> xsel<18> xsel<17> xsel<16>
+xsel<15> xsel<14> xsel<13> xsel<12> xsel<11> xsel<10> xsel<9> xsel<8> xsel<7>
+xsel<6> xsel<5> xsel<4> xsel<3> xsel<2> xsel<1> xsel<0> memarray_64x16
.ends memblock


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                                 9                                            *
* Block: Latch                                                                *
* Last Time Saved: Dec 12 09:40:01 2006                                       *
*******************************************************************************
.subckt Latch Q QN CLK D
XI8 QN net095 inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI6 Q net090 inv wn=1 wp=3 ln=0.18 lp=0.18 maxSheets=1
XI7 net044 D inv wn=0.3 wp=0.6 ln=0.18 lp=0.18 maxSheets=1
MN14 net30 vdd net81 gnd n18ll w=0.5 l=0.6
MN5 net090 net095 net81 gnd n18ll w=1.2 l=0.18
MN10 net81 D net78 gnd n18ll w=1.2 l=0.18
MN12 net30 net044 net78 gnd n18ll w=1.2 l=0.18
MN11 net095 net090 net30 gnd n18ll w=1.2 l=0.18
MN13 net78 CLK gnd gnd n18ll w=1.2 l=0.18
MP25 net090 CLK vdd vdd p18ll w=0.5 l=0.18
MP27 net095 CLK vdd vdd p18ll w=0.5 l=0.18
MP24 net090 net095 vdd vdd p18ll w=1.0 l=0.18
MP26 net095 net090 vdd vdd p18ll w=1.0 l=0.18
.ends Latch


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                          10                                                   *
* Block: sck_bar_gen                                                          *
* Last Time Saved: Dec 12 09:40:11 2006                                       *
*******************************************************************************
.subckt sck_bar_gen sck_bar CS ck_extern
XI0 sck net022 ck_extern CS Latch sheetSize=Asize maxSheets=1
XI24 sck_bar net030 inv maxSheets=1 ln=0.25 wp=3 wn=1.2 lp=0.25
XI17 sck_bar net036 inv maxSheets=1 lp=0.25 wn=1.2 wp=3 ln=0.25
XI23 sck_bar net030 inv maxSheets=1 lp=0.25 ln=0.25 wn=1.2 wp=3
XI21 net030 net038 inv maxSheets=1 lp=0.25 ln=0.25 wp=1.5 wn=0.6
XI20 net036 net038 inv maxSheets=1 ln=0.25 lp=0.25 wp=1.5 wn=0.6
XI22 sck_bar net036 inv maxSheets=1 lp=0.25 wn=1.2 wp=3 ln=0.25
XI13 net038 sck inv maxSheets=1 wn=0.6 wp=1.5 lp=0.25 ln=0.25
.ends sck_bar_gen


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                          11                                                   *
* Block: DFF                                                                  *
* Last Time Saved: Dec 15 13:40:04 2006                                       *
*******************************************************************************
.subckt DFF Q QN CK D
MN17 gnd net24 Q gnd n18ll w=0.6 l=0.18
MN16 gnd s QN gnd n18ll w=0.6 l=0.18
MN15 gnd net24 s gnd n18ll w=0.32 l=0.18
MN13 gnd m net15 gnd n18ll w=0.74 l=0.18
MN14 net20 s gnd gnd n18ll w=0.3 l=0.18
MN12 net20 cn net24 gnd n18ll w=0.3 l=0.18
MN10 net15 c net24 gnd n18ll w=0.74 l=0.18
MN8 net26 m gnd gnd n18ll w=0.3 l=0.18
MN7 gnd pm m gnd n18ll w=0.3 l=0.18
MN6 net26 c pm gnd n18ll w=0.3 l=0.18
MN3 gnd D net36 gnd n18ll w=0.3 l=0.18
MN2 net36 cn pm gnd n18ll w=0.3 l=0.18
MN0 gnd cn c gnd n18ll w=0.3 l=0.18
MN5 gnd CK cn gnd n18ll w=0.42 l=0.18
MP15 vdd s net60 vdd p18ll w=0.3 l=0.18
MP14 vdd net24 Q vdd p18ll w=0.9 l=0.18
MP13 vdd s QN vdd p18ll w=0.9 l=0.18
MP12 vdd net24 s vdd p18ll w=0.48 l=0.18
MP11 net66 m vdd vdd p18ll w=1.12 l=0.18
MP8 net66 cn net24 vdd p18ll w=1.12 l=0.18
MP7 net60 c net24 vdd p18ll w=0.3 l=0.18
MP5 vdd pm m vdd p18ll w=0.42 l=0.18
MP4 net75 m vdd vdd p18ll w=0.42 l=0.18
MP2 net75 cn pm vdd p18ll w=0.42 l=0.18
MP100 net77 c pm vdd p18ll w=0.42 l=0.18
MP1 vdd D net77 vdd p18ll w=0.42 l=0.18
MP0 vdd cn c vdd p18ll w=0.44 l=0.18
MP24 vdd CK cn vdd p18ll w=0.64 l=0.18
.ends DFF


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                          12                                                   *
* Block: ck_gen                                                               *
* Last Time Saved: Dec 12 09:43:35 2006                                       *
*******************************************************************************
.subckt ck_gen CK sck_bar
XI3 net16 net25 inv wn=0.4 wp=1 ln=0.25 lp=0.25 maxSheets=1
XI4 CK net16 inv wn=1 wp=3 ln=0.25 lp=0.25 maxSheets=1
XI2 net25 sck_bar inv maxSheets=1 ln=0.25 lp=0.25 wp=0.6 wn=0.3
.ends ck_gen


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                           13                                                  *
* Block: signals_gen                                                          *
* Last Time Saved: Dec 18 09:31:40 2006                                       *
*******************************************************************************
.subckt signals_gen addr<9> addr<8> addr<7> addr<6> addr<5> addr<4> addr<3>
+addr<2> addr<1> addr<0> addr_<9> addr_<8> addr_<7> addr_<6> addr_<5> addr_<4>
+addr_<3> addr_<2> addr_<1> addr_<0> rd_en wr_en wrdata<7> wrdata<6> wrdata<5>
+wrdata<4> wrdata<3> wrdata<2> wrdata<1> wrdata<0> wrdata_<7> wrdata_<6>
+wrdata_<5> wrdata_<4> wrdata_<3> wrdata_<2> wrdata_<1> wrdata_<0> A<9> A<8>
+A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> DIN<7> DIN<6> DIN<5> DIN<4> DIN<3>
+DIN<2> DIN<1> DIN<0> RD WR sck_bar
XI90_7 net023<0> net028<0> inv maxSheets=1 wn=0.22 lp=0.18 ln=0.18 wp=0.6
XI90_6 net023<1> net028<1> inv maxSheets=1 wn=0.22 lp=0.18 ln=0.18 wp=0.6
XI90_5 net023<2> net028<2> inv maxSheets=1 wn=0.22 lp=0.18 ln=0.18 wp=0.6
XI90_4 net023<3> net028<3> inv maxSheets=1 wn=0.22 lp=0.18 ln=0.18 wp=0.6
XI90_3 net023<4> net028<4> inv maxSheets=1 wn=0.22 lp=0.18 ln=0.18 wp=0.6
XI90_2 net023<5> net028<5> inv maxSheets=1 wn=0.22 lp=0.18 ln=0.18 wp=0.6
XI90_1 net023<6> net028<6> inv maxSheets=1 wn=0.22 lp=0.18 ln=0.18 wp=0.6
XI90_0 net023<7> net028<7> inv maxSheets=1 wn=0.22 lp=0.18 ln=0.18 wp=0.6
XI7_7 wrdata<7> net023<0> inv maxSheets=1 wn=1 lp=0.18 ln=0.18 wp=3
XI7_6 wrdata<6> net023<1> inv maxSheets=1 wn=1 lp=0.18 ln=0.18 wp=3
XI7_5 wrdata<5> net023<2> inv maxSheets=1 wn=1 lp=0.18 ln=0.18 wp=3
XI7_4 wrdata<4> net023<3> inv maxSheets=1 wn=1 lp=0.18 ln=0.18 wp=3
XI7_3 wrdata<3> net023<4> inv maxSheets=1 wn=1 lp=0.18 ln=0.18 wp=3
XI7_2 wrdata<2> net023<5> inv maxSheets=1 wn=1 lp=0.18 ln=0.18 wp=3
XI7_1 wrdata<1> net023<6> inv maxSheets=1 wn=1 lp=0.18 ln=0.18 wp=3
XI7_0 wrdata<0> net023<7> inv maxSheets=1 wn=1 lp=0.18 ln=0.18 wp=3
XI10_7 net017<0> net025<0> inv maxSheets=1 wp=0.6 ln=0.18 lp=0.18 wn=0.22
XI10_6 net017<1> net025<1> inv maxSheets=1 wp=0.6 ln=0.18 lp=0.18 wn=0.22
XI10_5 net017<2> net025<2> inv maxSheets=1 wp=0.6 ln=0.18 lp=0.18 wn=0.22
XI10_4 net017<3> net025<3> inv maxSheets=1 wp=0.6 ln=0.18 lp=0.18 wn=0.22
XI10_3 net017<4> net025<4> inv maxSheets=1 wp=0.6 ln=0.18 lp=0.18 wn=0.22
XI10_2 net017<5> net025<5> inv maxSheets=1 wp=0.6 ln=0.18 lp=0.18 wn=0.22
XI10_1 net017<6> net025<6> inv maxSheets=1 wp=0.6 ln=0.18 lp=0.18 wn=0.22
XI10_0 net017<7> net025<7> inv maxSheets=1 wp=0.6 ln=0.18 lp=0.18 wn=0.22
XI11_7 wrdata_<7> net017<0> inv maxSheets=1 ln=0.18 lp=0.18 wn=1 wp=3
XI11_6 wrdata_<6> net017<1> inv maxSheets=1 ln=0.18 lp=0.18 wn=1 wp=3
XI11_5 wrdata_<5> net017<2> inv maxSheets=1 ln=0.18 lp=0.18 wn=1 wp=3
XI11_4 wrdata_<4> net017<3> inv maxSheets=1 ln=0.18 lp=0.18 wn=1 wp=3
XI11_3 wrdata_<3> net017<4> inv maxSheets=1 ln=0.18 lp=0.18 wn=1 wp=3
XI11_2 wrdata_<2> net017<5> inv maxSheets=1 ln=0.18 lp=0.18 wn=1 wp=3
XI11_1 wrdata_<1> net017<6> inv maxSheets=1 ln=0.18 lp=0.18 wn=1 wp=3
XI11_0 wrdata_<0> net017<7> inv maxSheets=1 ln=0.18 lp=0.18 wn=1 wp=3
XI4_7 net028<0> net025<0> ck DIN<7> DFF sheetSize=Bsize maxSheets=1
XI4_6 net028<1> net025<1> ck DIN<6> DFF sheetSize=Bsize maxSheets=1
XI4_5 net028<2> net025<2> ck DIN<5> DFF sheetSize=Bsize maxSheets=1
XI4_4 net028<3> net025<3> ck DIN<4> DFF sheetSize=Bsize maxSheets=1
XI4_3 net028<4> net025<4> ck DIN<3> DFF sheetSize=Bsize maxSheets=1
XI4_2 net028<5> net025<5> ck DIN<2> DFF sheetSize=Bsize maxSheets=1
XI4_1 net028<6> net025<6> ck DIN<1> DFF sheetSize=Bsize maxSheets=1
XI4_0 net028<7> net025<7> ck DIN<0> DFF sheetSize=Bsize maxSheets=1
XI6 ck sck_bar ck_gen sheetSize=Asize maxSheets=1
XI2 rd_en net23 ck RD Latch maxSheets=1
XI1 wr_en net27 ck WR Latch maxSheets=1
XI0_9 addr<9> addr_<9> ck A<9> Latch maxSheets=1
XI0_8 addr<8> addr_<8> ck A<8> Latch maxSheets=1
XI0_7 addr<7> addr_<7> ck A<7> Latch maxSheets=1
XI0_6 addr<6> addr_<6> ck A<6> Latch maxSheets=1
XI0_5 addr<5> addr_<5> ck A<5> Latch maxSheets=1
XI0_4 addr<4> addr_<4> ck A<4> Latch maxSheets=1
XI0_3 addr<3> addr_<3> ck A<3> Latch maxSheets=1
XI0_2 addr<2> addr_<2> ck A<2> Latch maxSheets=1
XI0_1 addr<1> addr_<1> ck A<1> Latch maxSheets=1
XI0_0 addr<0> addr_<0> ck A<0> Latch maxSheets=1
.ends signals_gen


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                            14                                                 *
* Block: nor2                                                                 *
* Last Time Saved: Aug 18 08:30:12 2004                                       *
*******************************************************************************
.subckt nor2 Y A B lp=0.54 wp=5.4 ln=0.54 wn=2.7
MN1 Y A gnd gnd n18ll w=wn l=ln
MN0 Y B gnd gnd n18ll w=wn l=ln
MP0 Y B net8 vdd p18ll w=wp l=lp
MP1 net8 A vdd vdd p18ll w=wp l=lp
.ends nor2


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                               15                                              *
* Block: nand3                                                                *
* Last Time Saved: Aug 18 08:34:35 2004                                       *
*******************************************************************************
.subckt nand3 Y A B C lp=0.54 wp=5.4 ln=0.54 wn=2.7
MN1 Y A net14 gnd n18ll w=wn l=ln
MN0 net14 B net15 gnd n18ll w=wn l=ln
MN2 net15 C gnd gnd n18ll w=wn l=ln
MP1 Y B vdd vdd p18ll w=wp l=lp
MP0 Y C vdd vdd p18ll w=wp l=lp
MP2 Y A vdd vdd p18ll w=wp l=lp
.ends nand3


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                                 16                                            *
* Block: xdec                                                                 *
* Last Time Saved: Dec 12 09:45:28 2006                                       *
*******************************************************************************
.subckt xdec xsel<63> xsel<62> xsel<61> xsel<60> xsel<59> xsel<58> xsel<57>
+xsel<56> xsel<55> xsel<54> xsel<53> xsel<52> xsel<51> xsel<50> xsel<49>
+xsel<48> xsel<47> xsel<46> xsel<45> xsel<44> xsel<43> xsel<42> xsel<41>
+xsel<40> xsel<39> xsel<38> xsel<37> xsel<36> xsel<35> xsel<34> xsel<33>
+xsel<32> xsel<31> xsel<30> xsel<29> xsel<28> xsel<27> xsel<26> xsel<25>
+xsel<24> xsel<23> xsel<22> xsel<21> xsel<20> xsel<19> xsel<18> xsel<17>
+xsel<16> xsel<15> xsel<14> xsel<13> xsel<12> xsel<11> xsel<10> xsel<9> xsel<8>
+xsel<7> xsel<6> xsel<5> xsel<4> xsel<3> xsel<2> xsel<1> xsel<0> A<5> A<4> A<3>
+A<2> A<1> A<0> A_<5> A_<4> A_<3> A_<2> A_<1> A_<0>
XI2_63 xsel<63> net020<0> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_62 xsel<62> net020<1> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_61 xsel<61> net020<2> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_60 xsel<60> net020<3> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_59 xsel<59> net020<4> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_58 xsel<58> net020<5> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_57 xsel<57> net020<6> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_56 xsel<56> net020<7> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_55 xsel<55> net020<8> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_54 xsel<54> net020<9> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_53 xsel<53> net020<10> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_52 xsel<52> net020<11> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_51 xsel<51> net020<12> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_50 xsel<50> net020<13> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_49 xsel<49> net020<14> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_48 xsel<48> net020<15> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_47 xsel<47> net020<16> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_46 xsel<46> net020<17> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_45 xsel<45> net020<18> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_44 xsel<44> net020<19> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_43 xsel<43> net020<20> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_42 xsel<42> net020<21> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_41 xsel<41> net020<22> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_40 xsel<40> net020<23> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_39 xsel<39> net020<24> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_38 xsel<38> net020<25> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_37 xsel<37> net020<26> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_36 xsel<36> net020<27> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_35 xsel<35> net020<28> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_34 xsel<34> net020<29> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_33 xsel<33> net020<30> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_32 xsel<32> net020<31> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_31 xsel<31> net020<32> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_30 xsel<30> net020<33> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_29 xsel<29> net020<34> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_28 xsel<28> net020<35> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_27 xsel<27> net020<36> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_26 xsel<26> net020<37> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_25 xsel<25> net020<38> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_24 xsel<24> net020<39> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_23 xsel<23> net020<40> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_22 xsel<22> net020<41> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_21 xsel<21> net020<42> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_20 xsel<20> net020<43> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_19 xsel<19> net020<44> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_18 xsel<18> net020<45> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_17 xsel<17> net020<46> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_16 xsel<16> net020<47> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_15 xsel<15> net020<48> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_14 xsel<14> net020<49> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_13 xsel<13> net020<50> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_12 xsel<12> net020<51> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_11 xsel<11> net020<52> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_10 xsel<10> net020<53> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_9 xsel<9> net020<54> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_8 xsel<8> net020<55> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_7 xsel<7> net020<56> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_6 xsel<6> net020<57> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_5 xsel<5> net020<58> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_4 xsel<4> net020<59> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_3 xsel<3> net020<60> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_2 xsel<2> net020<61> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_1 xsel<1> net020<62> inv ln=0.18 wn=3 lp=0.18 wp=9
XI2_0 xsel<0> net020<63> inv ln=0.18 wn=3 lp=0.18 wp=9
XI10_63 net020<0> net024<0> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_62 net020<1> net024<1> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_61 net020<2> net024<2> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_60 net020<3> net024<3> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_59 net020<4> net024<4> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_58 net020<5> net024<5> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_57 net020<6> net024<6> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_56 net020<7> net024<7> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_55 net020<8> net024<8> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_54 net020<9> net024<9> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_53 net020<10> net024<10> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_52 net020<11> net024<11> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_51 net020<12> net024<12> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_50 net020<13> net024<13> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_49 net020<14> net024<14> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_48 net020<15> net024<15> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_47 net020<16> net024<16> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_46 net020<17> net024<17> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_45 net020<18> net024<18> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_44 net020<19> net024<19> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_43 net020<20> net024<20> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_42 net020<21> net024<21> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_41 net020<22> net024<22> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_40 net020<23> net024<23> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_39 net020<24> net024<24> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_38 net020<25> net024<25> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_37 net020<26> net024<26> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_36 net020<27> net024<27> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_35 net020<28> net024<28> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_34 net020<29> net024<29> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_33 net020<30> net024<30> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_32 net020<31> net024<31> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_31 net020<32> net024<32> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_30 net020<33> net024<33> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_29 net020<34> net024<34> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_28 net020<35> net024<35> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_27 net020<36> net024<36> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_26 net020<37> net024<37> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_25 net020<38> net024<38> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_24 net020<39> net024<39> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_23 net020<40> net024<40> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_22 net020<41> net024<41> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_21 net020<42> net024<42> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_20 net020<43> net024<43> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_19 net020<44> net024<44> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_18 net020<45> net024<45> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_17 net020<46> net024<46> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_16 net020<47> net024<47> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_15 net020<48> net024<48> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_14 net020<49> net024<49> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_13 net020<50> net024<50> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_12 net020<51> net024<51> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_11 net020<52> net024<52> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_10 net020<53> net024<53> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_9 net020<54> net024<54> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_8 net020<55> net024<55> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_7 net020<56> net024<56> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_6 net020<57> net024<57> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_5 net020<58> net024<58> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_4 net020<59> net024<59> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_3 net020<60> net024<60> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_2 net020<61> net024<61> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_1 net020<62> net024<62> inv ln=0.18 wn=1 lp=0.18 wp=3
XI10_0 net020<63> net024<63> inv ln=0.18 wn=1 lp=0.18 wp=3
XI26_63 net024<0> net029<0> net026<0> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_62 net024<1> net029<1> net026<1> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_61 net024<2> net029<2> net026<2> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_60 net024<3> net029<3> net026<3> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_59 net024<4> net029<4> net026<4> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_58 net024<5> net029<5> net026<5> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_57 net024<6> net029<6> net026<6> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_56 net024<7> net029<7> net026<7> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_55 net024<8> net029<8> net026<8> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_54 net024<9> net029<9> net026<9> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_53 net024<10> net029<10> net026<10> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_52 net024<11> net029<11> net026<11> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_51 net024<12> net029<12> net026<12> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_50 net024<13> net029<13> net026<13> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_49 net024<14> net029<14> net026<14> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_48 net024<15> net029<15> net026<15> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_47 net024<16> net029<16> net026<16> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_46 net024<17> net029<17> net026<17> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_45 net024<18> net029<18> net026<18> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_44 net024<19> net029<19> net026<19> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_43 net024<20> net029<20> net026<20> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_42 net024<21> net029<21> net026<21> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_41 net024<22> net029<22> net026<22> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_40 net024<23> net029<23> net026<23> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_39 net024<24> net029<24> net026<24> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_38 net024<25> net029<25> net026<25> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_37 net024<26> net029<26> net026<26> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_36 net024<27> net029<27> net026<27> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_35 net024<28> net029<28> net026<28> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_34 net024<29> net029<29> net026<29> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_33 net024<30> net029<30> net026<30> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_32 net024<31> net029<31> net026<31> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_31 net024<32> net029<32> net026<32> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_30 net024<33> net029<33> net026<33> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_29 net024<34> net029<34> net026<34> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_28 net024<35> net029<35> net026<35> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_27 net024<36> net029<36> net026<36> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_26 net024<37> net029<37> net026<37> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_25 net024<38> net029<38> net026<38> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_24 net024<39> net029<39> net026<39> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_23 net024<40> net029<40> net026<40> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_22 net024<41> net029<41> net026<41> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_21 net024<42> net029<42> net026<42> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_20 net024<43> net029<43> net026<43> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_19 net024<44> net029<44> net026<44> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_18 net024<45> net029<45> net026<45> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_17 net024<46> net029<46> net026<46> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_16 net024<47> net029<47> net026<47> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_15 net024<48> net029<48> net026<48> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_14 net024<49> net029<49> net026<49> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_13 net024<50> net029<50> net026<50> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_12 net024<51> net029<51> net026<51> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_11 net024<52> net029<52> net026<52> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_10 net024<53> net029<53> net026<53> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_9 net024<54> net029<54> net026<54> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_8 net024<55> net029<55> net026<55> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_7 net024<56> net029<56> net026<56> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_6 net024<57> net029<57> net026<57> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_5 net024<58> net029<58> net026<58> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_4 net024<59> net029<59> net026<59> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_3 net024<60> net029<60> net026<60> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_2 net024<61> net029<61> net026<61> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_1 net024<62> net029<62> net026<62> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI26_0 net024<63> net029<63> net026<63> nor2 lp=0.18 wp=1.5 ln=0.18 wn=0.5
XI25_63 net029<0> A<0> A<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_62 net029<1> A_<0> A<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_61 net029<2> A<0> A_<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_60 net029<3> A_<0> A_<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_59 net029<4> A<0> A<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_58 net029<5> A_<0> A<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_57 net029<6> A<0> A_<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_56 net029<7> A_<0> A_<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_55 net029<8> A<0> A<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_54 net029<9> A_<0> A<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_53 net029<10> A<0> A_<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_52 net029<11> A_<0> A_<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_51 net029<12> A<0> A<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_50 net029<13> A_<0> A<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_49 net029<14> A<0> A_<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_48 net029<15> A_<0> A_<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_47 net029<16> A<0> A<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_46 net029<17> A_<0> A<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_45 net029<18> A<0> A_<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_44 net029<19> A_<0> A_<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_43 net029<20> A<0> A<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_42 net029<21> A_<0> A<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_41 net029<22> A<0> A_<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_40 net029<23> A_<0> A_<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_39 net029<24> A<0> A<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_38 net029<25> A_<0> A<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_37 net029<26> A<0> A_<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_36 net029<27> A_<0> A_<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_35 net029<28> A<0> A<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_34 net029<29> A_<0> A<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_33 net029<30> A<0> A_<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_32 net029<31> A_<0> A_<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_31 net029<32> A<0> A<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_30 net029<33> A_<0> A<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_29 net029<34> A<0> A_<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_28 net029<35> A_<0> A_<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_27 net029<36> A<0> A<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_26 net029<37> A_<0> A<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_25 net029<38> A<0> A_<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_24 net029<39> A_<0> A_<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_23 net029<40> A<0> A<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_22 net029<41> A_<0> A<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_21 net029<42> A<0> A_<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_20 net029<43> A_<0> A_<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_19 net029<44> A<0> A<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_18 net029<45> A_<0> A<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_17 net029<46> A<0> A_<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_16 net029<47> A_<0> A_<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_15 net029<48> A<0> A<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_14 net029<49> A_<0> A<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_13 net029<50> A<0> A_<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_12 net029<51> A_<0> A_<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_11 net029<52> A<0> A<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_10 net029<53> A_<0> A<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_9 net029<54> A<0> A_<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_8 net029<55> A_<0> A_<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_7 net029<56> A<0> A<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_6 net029<57> A_<0> A<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_5 net029<58> A<0> A_<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_4 net029<59> A_<0> A_<1> A<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_3 net029<60> A<0> A<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_2 net029<61> A_<0> A<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_1 net029<62> A<0> A_<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI25_0 net029<63> A_<0> A_<1> A_<2> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_63 net026<0> A<3> A<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_62 net026<1> A<3> A<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_61 net026<2> A<3> A<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_60 net026<3> A<3> A<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_59 net026<4> A<3> A<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_58 net026<5> A<3> A<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_57 net026<6> A<3> A<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_56 net026<7> A<3> A<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_55 net026<8> A_<3> A<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_54 net026<9> A_<3> A<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_53 net026<10> A_<3> A<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_52 net026<11> A_<3> A<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_51 net026<12> A_<3> A<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_50 net026<13> A_<3> A<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_49 net026<14> A_<3> A<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_48 net026<15> A_<3> A<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_47 net026<16> A<3> A_<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_46 net026<17> A<3> A_<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_45 net026<18> A<3> A_<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_44 net026<19> A<3> A_<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_43 net026<20> A<3> A_<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_42 net026<21> A<3> A_<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_41 net026<22> A<3> A_<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_40 net026<23> A<3> A_<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_39 net026<24> A_<3> A_<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_38 net026<25> A_<3> A_<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_37 net026<26> A_<3> A_<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_36 net026<27> A_<3> A_<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_35 net026<28> A_<3> A_<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_34 net026<29> A_<3> A_<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_33 net026<30> A_<3> A_<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_32 net026<31> A_<3> A_<4> A<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_31 net026<32> A<3> A<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_30 net026<33> A<3> A<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_29 net026<34> A<3> A<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_28 net026<35> A<3> A<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_27 net026<36> A<3> A<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_26 net026<37> A<3> A<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_25 net026<38> A<3> A<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_24 net026<39> A<3> A<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_23 net026<40> A_<3> A<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_22 net026<41> A_<3> A<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_21 net026<42> A_<3> A<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_20 net026<43> A_<3> A<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_19 net026<44> A_<3> A<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_18 net026<45> A_<3> A<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_17 net026<46> A_<3> A<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_16 net026<47> A_<3> A<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_15 net026<48> A<3> A_<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_14 net026<49> A<3> A_<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_13 net026<50> A<3> A_<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_12 net026<51> A<3> A_<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_11 net026<52> A<3> A_<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_10 net026<53> A<3> A_<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_9 net026<54> A<3> A_<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_8 net026<55> A<3> A_<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_7 net026<56> A_<3> A_<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_6 net026<57> A_<3> A_<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_5 net026<58> A_<3> A_<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_4 net026<59> A_<3> A_<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_3 net026<60> A_<3> A_<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_2 net026<61> A_<3> A_<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_1 net026<62> A_<3> A_<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
XI24_0 net026<63> A_<3> A_<4> A_<5> nand3 lp=0.18 wp=0.4 ln=0.18 wn=0.4
.ends xdec


*******************************************************************************
* Sub-Circuit Netlist:                                                        *
*                                 17                                            *
* Block: ydec                                                                 *
* Last Time Saved: Dec 12 09:44:20 2006                                       *
*******************************************************************************
.subckt ydec ysel<15> ysel<14> ysel<13> ysel<12> ysel<11> ysel<10> ysel<9>
+ysel<8> ysel<7> ysel<6> ysel<5> ysel<4> ysel<3> ysel<2> ysel<1> ysel<0> A<9>
+A<8> A<7> A<6> A_<9> A_<8> A_<7> A_<6>
XI3_15 net014<0> net018<0> net017<0> nor2 wp=1.5 lp=0.18 ln=0.18 maxSheets=1
+wn=0.5
XI3_14 net014<1> net018<1> net017<1> nor2 wp=1.5 lp=0.18 ln=0.18 maxSheets=1
+wn=0.5
XI3_13 net014<2> net018<2> net017<2> nor2 wp=1.5 lp=0.18 ln=0.18 maxSheets=1
+wn=0.5
XI3_12 net014<3> net018<3> net017<3> nor2 wp=1.5 lp=0.18 ln=0.18 maxSheets=1
+wn=0.5
XI3_11 net014<4> net018<4> net017<4> nor2 wp=1.5 lp=0.18 ln=0.18 maxSheets=1
+wn=0.5
XI3_10 net014<5> net018<5> net017<5> nor2 wp=1.5 lp=0.18 ln=0.18 maxSheets=1
+wn=0.5
XI3_9 net014<6> net018<6> net017<6> nor2 wp=1.5 lp=0.18 ln=0.18 maxSheets=1
+wn=0.5
XI3_8 net014<7> net018<7> net017<7> nor2 wp=1.5 lp=0.18 ln=0.18 maxSheets=1
+wn=0.5
XI3_7 net014<8> net018<8> net017<8> nor2 wp=1.5 lp=0.18 ln=0.18 maxSheets=1
+wn=0.5
XI3_6 net014<9> net018<9> net017<9> nor2 wp=1.5 lp=0.18 ln=0.18 maxSheets=1
+wn=0.5
XI3_5 net014<10> net018<10> net017<10> nor2 wp=1.5 lp=0.18 ln=0.18 maxSheets=1
+wn=0.5
XI3_4 net014<11> net018<11> net017<11> nor2 wp=1.5 lp=0.18 ln=0.18 maxSheets=1
+wn=0.5
XI3_3 net014<12> net018<12> net017<12> nor2 wp=1.5 lp=0.18 ln=0.18 maxSheets=1
+wn=0.5
XI3_2 net014<13> net018<13> net017<13> nor2 wp=1.5 lp=0.18 ln=0.18 maxSheets=1
+wn=0.5
XI3_1 net014<14> net018<14> net017<14> nor2 wp=1.5 lp=0.18 ln=0.18 maxSheets=1
+wn=0.5
XI3_0 net014<15> net018<15> net017<15> nor2 wp=2 lp=0.18 ln=0.18 maxSheets=1
+wn=0.5
XI1_15 net018<0> A<6> A<7> nand2 lp=0.18 ln=0.18 maxSheets=1 wp=0.5 wn=0.5
XI1_14 net018<1> A_<6> A<7> nand2 lp=0.18 ln=0.18 maxSheets=1 wp=0.5 wn=0.5
XI1_13 net018<2> A<6> A_<7> nand2 lp=0.18 ln=0.18 maxSheets=1 wp=0.5 wn=0.5
XI1_12 net018<3> A_<6> A_<7> nand2 lp=0.18 ln=0.18 maxSheets=1 wp=0.5 wn=0.5
XI1_11 net018<4> A<6> A<7> nand2 lp=0.18 ln=0.18 maxSheets=1 wp=0.5 wn=0.5
XI1_10 net018<5> A_<6> A<7> nand2 lp=0.18 ln=0.18 maxSheets=1 wp=0.5 wn=0.5
XI1_9 net018<6> A<6> A_<7> nand2 lp=0.18 ln=0.18 maxSheets=1 wp=0.5 wn=0.5
XI1_8 net018<7> A_<6> A_<7> nand2 lp=0.18 ln=0.18 maxSheets=1 wp=0.5 wn=0.5
XI1_7 net018<8> A<6> A<7> nand2 lp=0.18 ln=0.18 maxSheets=1 wp=0.5 wn=0.5
XI1_6 net018<9> A_<6> A<7> nand2 lp=0.18 ln=0.18 maxSheets=1 wp=0.5 wn=0.5
XI1_5 net018<10> A<6> A_<7> nand2 lp=0.18 ln=0.18 maxSheets=1 wp=0.5 wn=0.5
XI1_4 net018<11> A_<6> A_<7> nand2 lp=0.18 ln=0.18 maxSheets=1 wp=0.5 wn=0.5
XI1_3 net018<12> A<6> A<7> nand2 lp=0.18 ln=0.18 maxSheets=1 wp=0.5 wn=0.5
XI1_2 net018<13> A_<6> A<7> nand2 lp=0.18 ln=0.18 maxSheets=1 wp=0.5 wn=0.5
XI1_1 net018<14> A<6> A_<7> nand2 lp=0.18 ln=0.18 maxSheets=1 wp=0.5 wn=0.5
XI1_0 net018<15> A_<6> A_<7> nand2 lp=0.18 ln=0.18 maxSheets=1 wp=0.5 wn=0.5
XI2_15 net017<0> A<8> A<9> nand2 maxSheets=1 ln=0.18 lp=0.18 wp=0.5 wn=0.5
XI2_14 net017<1> A<8> A<9> nand2 maxSheets=1 ln=0.18 lp=0.18 wp=0.5 wn=0.5
XI2_13 net017<2> A<8> A<9> nand2 maxSheets=1 ln=0.18 lp=0.18 wp=0.5 wn=0.5
XI2_12 net017<3> A<8> A<9> nand2 maxSheets=1 ln=0.18 lp=0.18 wp=0.5 wn=0.5
XI2_11 net017<4> A_<8> A<9> nand2 maxSheets=1 ln=0.18 lp=0.18 wp=0.5 wn=0.5
XI2_10 net017<5> A_<8> A<9> nand2 maxSheets=1 ln=0.18 lp=0.18 wp=0.5 wn=0.5
XI2_9 net017<6> A_<8> A<9> nand2 maxSheets=1 ln=0.18 lp=0.18 wp=0.5 wn=0.5
XI2_8 net017<7> A_<8> A<9> nand2 maxSheets=1 ln=0.18 lp=0.18 wp=0.5 wn=0.5
XI2_7 net017<8> A<8> A_<9> nand2 maxSheets=1 ln=0.18 lp=0.18 wp=0.5 wn=0.5
XI2_6 net017<9> A<8> A_<9> nand2 maxSheets=1 ln=0.18 lp=0.18 wp=0.5 wn=0.5
XI2_5 net017<10> A<8> A_<9> nand2 maxSheets=1 ln=0.18 lp=0.18 wp=0.5 wn=0.5
XI2_4 net017<11> A<8> A_<9> nand2 maxSheets=1 ln=0.18 lp=0.18 wp=0.5 wn=0.5
XI2_3 net017<12> A_<8> A_<9> nand2 maxSheets=1 ln=0.18 lp=0.18 wp=0.5 wn=0.5
XI2_2 net017<13> A_<8> A_<9> nand2 maxSheets=1 ln=0.18 lp=0.18 wp=0.5 wn=0.5
XI2_1 net017<14> A_<8> A_<9> nand2 maxSheets=1 ln=0.18 lp=0.18 wp=0.5 wn=0.5
XI2_0 net017<15> A_<8> A_<9> nand2 maxSheets=1 ln=0.18 lp=0.18 wp=0.5 wn=0.5
XI4_15 net021<0> net014<0> inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI4_14 net021<1> net014<1> inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI4_13 net021<2> net014<2> inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI4_12 net021<3> net014<3> inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI4_11 net021<4> net014<4> inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI4_10 net021<5> net014<5> inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI4_9 net021<6> net014<6> inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI4_8 net021<7> net014<7> inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI4_7 net021<8> net014<8> inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI4_6 net021<9> net014<9> inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI4_5 net021<10> net014<10> inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI4_4 net021<11> net014<11> inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI4_3 net021<12> net014<12> inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI4_2 net021<13> net014<13> inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI4_1 net021<14> net014<14> inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI4_0 net021<15> net014<15> inv lp=0.18 ln=0.18 wp=3 wn=1 maxSheets=1
XI7_15 ysel<15> net021<0> inv lp=0.18 ln=0.18 wp=9 wn=3 maxSheets=1
XI7_14 ysel<14> net021<1> inv lp=0.18 ln=0.18 wp=9 wn=3 maxSheets=1
XI7_13 ysel<13> net021<2> inv lp=0.18 ln=0.18 wp=9 wn=3 maxSheets=1
XI7_12 ysel<12> net021<3> inv lp=0.18 ln=0.18 wp=9 wn=3 maxSheets=1
XI7_11 ysel<11> net021<4> inv lp=0.18 ln=0.18 wp=9 wn=3 maxSheets=1
XI7_10 ysel<10> net021<5> inv lp=0.18 ln=0.18 wp=9 wn=3 maxSheets=1
XI7_9 ysel<9> net021<6> inv lp=0.18 ln=0.18 wp=9 wn=3 maxSheets=1
XI7_8 ysel<8> net021<7> inv lp=0.18 ln=0.18 wp=9 wn=3 maxSheets=1
XI7_7 ysel<7> net021<8> inv lp=0.18 ln=0.18 wp=9 wn=3 maxSheets=1
XI7_6 ysel<6> net021<9> inv lp=0.18 ln=0.18 wp=9 wn=3 maxSheets=1
XI7_5 ysel<5> net021<10> inv lp=0.18 ln=0.18 wp=9 wn=3 maxSheets=1
XI7_4 ysel<4> net021<11> inv lp=0.18 ln=0.18 wp=9 wn=3 maxSheets=1
XI7_3 ysel<3> net021<12> inv lp=0.18 ln=0.18 wp=9 wn=3 maxSheets=1
XI7_2 ysel<2> net021<13> inv lp=0.18 ln=0.18 wp=9 wn=3 maxSheets=1
XI7_1 ysel<1> net021<14> inv lp=0.18 ln=0.18 wp=9 wn=3 maxSheets=1
XI7_0 ysel<0> net021<15> inv lp=0.18 ln=0.18 wp=9 wn=3 maxSheets=1
.ends ydec


*******************************************************************************
* Main Circuit Netlist:                                                       *
*                            18                                                 *
* Block: RAM_1kx8                                                             *
* Last Time Saved: Dec 19 09:16:36 2006                                       *
*******************************************************************************
.subckt ram DOUT<7> DOUT<6> DOUT<5> DOUT<4> DOUT<3> DOUT<2> DOUT<1>
+DOUT<0> A<9> A<8> A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> CLK CS DIN<7> DIN<6>
+DIN<5> DIN<4> DIN<3> DIN<2> DIN<1> DIN<0> RD WR
XI11_7 DOUT<7> rd_en sck_bar wr_en wrdata<7> wrdata_<7> xsel<63> xsel<62>
+xsel<61> xsel<60> xsel<59> xsel<58> xsel<57> xsel<56> xsel<55> xsel<54>
+xsel<53> xsel<52> xsel<51> xsel<50> xsel<49> xsel<48> xsel<47> xsel<46>
+xsel<45> xsel<44> xsel<43> xsel<42> xsel<41> xsel<40> xsel<39> xsel<38>
+xsel<37> xsel<36> xsel<35> xsel<34> xsel<33> xsel<32> xsel<31> xsel<30>
+xsel<29> xsel<28> xsel<27> xsel<26> xsel<25> xsel<24> xsel<23> xsel<22>
+xsel<21> xsel<20> xsel<19> xsel<18> xsel<17> xsel<16> xsel<15> xsel<14>
+xsel<13> xsel<12> xsel<11> xsel<10> xsel<9> xsel<8> xsel<7> xsel<6> xsel<5>
+xsel<4> xsel<3> xsel<2> xsel<1> xsel<0> ysel<15> ysel<14> ysel<13> ysel<12>
+ysel<11> ysel<10> ysel<9> ysel<8> ysel<7> ysel<6> ysel<5> ysel<4> ysel<3>
+ysel<2> ysel<1> ysel<0> memblock maxSheets=1 sheetSize=Bsize
XI11_6 DOUT<6> rd_en sck_bar wr_en wrdata<6> wrdata_<6> xsel<63> xsel<62>
+xsel<61> xsel<60> xsel<59> xsel<58> xsel<57> xsel<56> xsel<55> xsel<54>
+xsel<53> xsel<52> xsel<51> xsel<50> xsel<49> xsel<48> xsel<47> xsel<46>
+xsel<45> xsel<44> xsel<43> xsel<42> xsel<41> xsel<40> xsel<39> xsel<38>
+xsel<37> xsel<36> xsel<35> xsel<34> xsel<33> xsel<32> xsel<31> xsel<30>
+xsel<29> xsel<28> xsel<27> xsel<26> xsel<25> xsel<24> xsel<23> xsel<22>
+xsel<21> xsel<20> xsel<19> xsel<18> xsel<17> xsel<16> xsel<15> xsel<14>
+xsel<13> xsel<12> xsel<11> xsel<10> xsel<9> xsel<8> xsel<7> xsel<6> xsel<5>
+xsel<4> xsel<3> xsel<2> xsel<1> xsel<0> ysel<15> ysel<14> ysel<13> ysel<12>
+ysel<11> ysel<10> ysel<9> ysel<8> ysel<7> ysel<6> ysel<5> ysel<4> ysel<3>
+ysel<2> ysel<1> ysel<0> memblock maxSheets=1 sheetSize=Bsize
XI11_5 DOUT<5> rd_en sck_bar wr_en wrdata<5> wrdata_<5> xsel<63> xsel<62>
+xsel<61> xsel<60> xsel<59> xsel<58> xsel<57> xsel<56> xsel<55> xsel<54>
+xsel<53> xsel<52> xsel<51> xsel<50> xsel<49> xsel<48> xsel<47> xsel<46>
+xsel<45> xsel<44> xsel<43> xsel<42> xsel<41> xsel<40> xsel<39> xsel<38>
+xsel<37> xsel<36> xsel<35> xsel<34> xsel<33> xsel<32> xsel<31> xsel<30>
+xsel<29> xsel<28> xsel<27> xsel<26> xsel<25> xsel<24> xsel<23> xsel<22>
+xsel<21> xsel<20> xsel<19> xsel<18> xsel<17> xsel<16> xsel<15> xsel<14>
+xsel<13> xsel<12> xsel<11> xsel<10> xsel<9> xsel<8> xsel<7> xsel<6> xsel<5>
+xsel<4> xsel<3> xsel<2> xsel<1> xsel<0> ysel<15> ysel<14> ysel<13> ysel<12>
+ysel<11> ysel<10> ysel<9> ysel<8> ysel<7> ysel<6> ysel<5> ysel<4> ysel<3>
+ysel<2> ysel<1> ysel<0> memblock maxSheets=1 sheetSize=Bsize
XI11_4 DOUT<4> rd_en sck_bar wr_en wrdata<4> wrdata_<4> xsel<63> xsel<62>
+xsel<61> xsel<60> xsel<59> xsel<58> xsel<57> xsel<56> xsel<55> xsel<54>
+xsel<53> xsel<52> xsel<51> xsel<50> xsel<49> xsel<48> xsel<47> xsel<46>
+xsel<45> xsel<44> xsel<43> xsel<42> xsel<41> xsel<40> xsel<39> xsel<38>
+xsel<37> xsel<36> xsel<35> xsel<34> xsel<33> xsel<32> xsel<31> xsel<30>
+xsel<29> xsel<28> xsel<27> xsel<26> xsel<25> xsel<24> xsel<23> xsel<22>
+xsel<21> xsel<20> xsel<19> xsel<18> xsel<17> xsel<16> xsel<15> xsel<14>
+xsel<13> xsel<12> xsel<11> xsel<10> xsel<9> xsel<8> xsel<7> xsel<6> xsel<5>
+xsel<4> xsel<3> xsel<2> xsel<1> xsel<0> ysel<15> ysel<14> ysel<13> ysel<12>
+ysel<11> ysel<10> ysel<9> ysel<8> ysel<7> ysel<6> ysel<5> ysel<4> ysel<3>
+ysel<2> ysel<1> ysel<0> memblock maxSheets=1 sheetSize=Bsize
XI11_3 DOUT<3> rd_en sck_bar wr_en wrdata<3> wrdata_<3> xsel<63> xsel<62>
+xsel<61> xsel<60> xsel<59> xsel<58> xsel<57> xsel<56> xsel<55> xsel<54>
+xsel<53> xsel<52> xsel<51> xsel<50> xsel<49> xsel<48> xsel<47> xsel<46>
+xsel<45> xsel<44> xsel<43> xsel<42> xsel<41> xsel<40> xsel<39> xsel<38>
+xsel<37> xsel<36> xsel<35> xsel<34> xsel<33> xsel<32> xsel<31> xsel<30>
+xsel<29> xsel<28> xsel<27> xsel<26> xsel<25> xsel<24> xsel<23> xsel<22>
+xsel<21> xsel<20> xsel<19> xsel<18> xsel<17> xsel<16> xsel<15> xsel<14>
+xsel<13> xsel<12> xsel<11> xsel<10> xsel<9> xsel<8> xsel<7> xsel<6> xsel<5>
+xsel<4> xsel<3> xsel<2> xsel<1> xsel<0> ysel<15> ysel<14> ysel<13> ysel<12>
+ysel<11> ysel<10> ysel<9> ysel<8> ysel<7> ysel<6> ysel<5> ysel<4> ysel<3>
+ysel<2> ysel<1> ysel<0> memblock maxSheets=1 sheetSize=Bsize
XI11_2 DOUT<2> rd_en sck_bar wr_en wrdata<2> wrdata_<2> xsel<63> xsel<62>
+xsel<61> xsel<60> xsel<59> xsel<58> xsel<57> xsel<56> xsel<55> xsel<54>
+xsel<53> xsel<52> xsel<51> xsel<50> xsel<49> xsel<48> xsel<47> xsel<46>
+xsel<45> xsel<44> xsel<43> xsel<42> xsel<41> xsel<40> xsel<39> xsel<38>
+xsel<37> xsel<36> xsel<35> xsel<34> xsel<33> xsel<32> xsel<31> xsel<30>
+xsel<29> xsel<28> xsel<27> xsel<26> xsel<25> xsel<24> xsel<23> xsel<22>
+xsel<21> xsel<20> xsel<19> xsel<18> xsel<17> xsel<16> xsel<15> xsel<14>
+xsel<13> xsel<12> xsel<11> xsel<10> xsel<9> xsel<8> xsel<7> xsel<6> xsel<5>
+xsel<4> xsel<3> xsel<2> xsel<1> xsel<0> ysel<15> ysel<14> ysel<13> ysel<12>
+ysel<11> ysel<10> ysel<9> ysel<8> ysel<7> ysel<6> ysel<5> ysel<4> ysel<3>
+ysel<2> ysel<1> ysel<0> memblock maxSheets=1 sheetSize=Bsize
XI11_1 DOUT<1> rd_en sck_bar wr_en wrdata<1> wrdata_<1> xsel<63> xsel<62>
+xsel<61> xsel<60> xsel<59> xsel<58> xsel<57> xsel<56> xsel<55> xsel<54>
+xsel<53> xsel<52> xsel<51> xsel<50> xsel<49> xsel<48> xsel<47> xsel<46>
+xsel<45> xsel<44> xsel<43> xsel<42> xsel<41> xsel<40> xsel<39> xsel<38>
+xsel<37> xsel<36> xsel<35> xsel<34> xsel<33> xsel<32> xsel<31> xsel<30>
+xsel<29> xsel<28> xsel<27> xsel<26> xsel<25> xsel<24> xsel<23> xsel<22>
+xsel<21> xsel<20> xsel<19> xsel<18> xsel<17> xsel<16> xsel<15> xsel<14>
+xsel<13> xsel<12> xsel<11> xsel<10> xsel<9> xsel<8> xsel<7> xsel<6> xsel<5>
+xsel<4> xsel<3> xsel<2> xsel<1> xsel<0> ysel<15> ysel<14> ysel<13> ysel<12>
+ysel<11> ysel<10> ysel<9> ysel<8> ysel<7> ysel<6> ysel<5> ysel<4> ysel<3>
+ysel<2> ysel<1> ysel<0> memblock maxSheets=1 sheetSize=Bsize
XI11_0 DOUT<0> rd_en sck_bar wr_en wrdata<0> wrdata_<0> xsel<63> xsel<62>
+xsel<61> xsel<60> xsel<59> xsel<58> xsel<57> xsel<56> xsel<55> xsel<54>
+xsel<53> xsel<52> xsel<51> xsel<50> xsel<49> xsel<48> xsel<47> xsel<46>
+xsel<45> xsel<44> xsel<43> xsel<42> xsel<41> xsel<40> xsel<39> xsel<38>
+xsel<37> xsel<36> xsel<35> xsel<34> xsel<33> xsel<32> xsel<31> xsel<30>
+xsel<29> xsel<28> xsel<27> xsel<26> xsel<25> xsel<24> xsel<23> xsel<22>
+xsel<21> xsel<20> xsel<19> xsel<18> xsel<17> xsel<16> xsel<15> xsel<14>
+xsel<13> xsel<12> xsel<11> xsel<10> xsel<9> xsel<8> xsel<7> xsel<6> xsel<5>
+xsel<4> xsel<3> xsel<2> xsel<1> xsel<0> ysel<15> ysel<14> ysel<13> ysel<12>
+ysel<11> ysel<10> ysel<9> ysel<8> ysel<7> ysel<6> ysel<5> ysel<4> ysel<3>
+ysel<2> ysel<1> ysel<0> memblock maxSheets=1 sheetSize=Bsize
XI10 sck_bar CS CLK sck_bar_gen maxSheets=1 sheetSize=Asize
XI5 addr<9> addr<8> addr<7> addr<6> addr<5> addr<4> addr<3> addr<2> addr<1>
+addr<0> addr_<9> addr_<8> addr_<7> addr_<6> addr_<5> addr_<4> addr_<3>
+addr_<2> addr_<1> addr_<0> rd_en wr_en wrdata<7> wrdata<6> wrdata<5> wrdata<4>
+wrdata<3> wrdata<2> wrdata<1> wrdata<0> wrdata_<7> wrdata_<6> wrdata_<5>
+wrdata_<4> wrdata_<3> wrdata_<2> wrdata_<1> wrdata_<0> A<9> A<8> A<7> A<6>
+A<5> A<4> A<3> A<2> A<1> A<0> DIN<7> DIN<6> DIN<5> DIN<4> DIN<3> DIN<2> DIN<1>
+DIN<0> RD WR sck_bar signals_gen maxSheets=1 sheetSize=Asize
XI2 xsel<63> xsel<62> xsel<61> xsel<60> xsel<59> xsel<58> xsel<57> xsel<56>
+xsel<55> xsel<54> xsel<53> xsel<52> xsel<51> xsel<50> xsel<49> xsel<48>
+xsel<47> xsel<46> xsel<45> xsel<44> xsel<43> xsel<42> xsel<41> xsel<40>
+xsel<39> xsel<38> xsel<37> xsel<36> xsel<35> xsel<34> xsel<33> xsel<32>
+xsel<31> xsel<30> xsel<29> xsel<28> xsel<27> xsel<26> xsel<25> xsel<24>
+xsel<23> xsel<22> xsel<21> xsel<20> xsel<19> xsel<18> xsel<17> xsel<16>
+xsel<15> xsel<14> xsel<13> xsel<12> xsel<11> xsel<10> xsel<9> xsel<8> xsel<7>
+xsel<6> xsel<5> xsel<4> xsel<3> xsel<2> xsel<1> xsel<0> addr<5> addr<4>
+addr<3> addr<2> addr<1> addr<0> addr_<5> addr_<4> addr_<3> addr_<2> addr_<1>
+addr_<0> xdec maxSheets=1 sheetSize=Asize
XI6 ysel<15> ysel<14> ysel<13> ysel<12> ysel<11> ysel<10> ysel<9> ysel<8>
+ysel<7> ysel<6> ysel<5> ysel<4> ysel<3> ysel<2> ysel<1> ysel<0> addr<9>
+addr<8> addr<7> addr<6> addr_<9> addr_<8> addr_<7>  ydec maxSheets=1
+sheetSize=Asize
.ends ram 

*******************************************************************************
* Main Circuit Netlist:                                                       *
*                           19                                                  *
* Block: QDFFRBN                                                            *
* Last Time Saved: Dec 19 09:16:36 2006                                       *
*******************************************************************************


.SUBCKT QDFFRBN Q  D  CK  RB  VDD  VSS  
MMI_96 G1 CK1 G2 VDD P_18_G2 l=1.8e-07 w=4.4e-07
MMI_164 RL CK1 MPW VDD P_18_G2 l=1.8e-07 w=4.4e-07
MMI_165 G2 CKB G4 VDD P_18_G2 l=1.8e-07 w=4.4e-07
MMI_166 G3 CKB RL VDD P_18_G2 l=1.8e-07 w=1.04e-06
MMI_160 RL CKB MPW VSS N_18_G2 l=1.8e-07 w=4.4e-07
MMI_89 G1 CKB G2 VSS N_18_G2 l=1.8e-07 w=4.4e-07
MMI_161 G3 CK1 RL VSS N_18_G2 l=1.8e-07 w=7.6e-07
MMI_162 G2 CK1 G4 VSS N_18_G2 l=1.8e-07 w=4.4e-07
XG9 RB G3 G4 DECAP_NAND2_G9
XG10 RB RL QB1 DECAP_NAND2_G10
XG11 D G1 DECAP_INV_G11
XG12 CK CKB DECAP_INV_G12
XG13 CKB CK1 DECAP_INV_G12
XG14 G2 G3 DECAP_INV_G13
XG15 QB1 MPW DECAP_INV_G12
XG16 QB1 Q DECAP_INV_G14
.ENDS


*******************************************************************************
* Main Circuit Netlist:                                                       *
*                            20                                                 *
* Block: DBZRSBN                                                          *
* Last Time Saved: Dec 19 09:16:36 2006                                       *
*******************************************************************************
.SUBCKT DBZRSBN Q  QB  D  TD  CKB  SEL  RB  SB  VDD  VSS  
MMI_151 G1 D N_9 VDD P_18_G2 l=1.8e-07 w=1.83e-06
MMI171 G1 SELB N_7 VDD P_18_G2 l=1.8e-07 w=4.4e-07
MMI172 N_7 TD VDD VDD P_18_G2 l=1.8e-07 w=4.4e-07
MMI_152 N_9 SEL VDD VDD P_18_G2 l=1.8e-07 w=1.03e-06
MMI_96 G1 CK1 G2 VDD P_18_G2 l=1.8e-07 w=4.4e-07
MMI_164 RL CK1 MPW VDD P_18_G2 l=1.8e-07 w=4.4e-07
MMI_165 G2 CKB1 G4 VDD P_18_G2 l=1.8e-07 w=4.4e-07
MMI_166 G3 CKB1 RL VDD P_18_G2 l=1.8e-07 w=1.04e-06
MMI_156 G1 D N_10 VSS N_18_G2 l=1.8e-07 w=1e-06
MMI_155 N_10 SELB VSS VSS N_18_G2 l=1.8e-07 w=8.5e-07
MMI173 N_8 TD VSS VSS N_18_G2 l=1.8e-07 w=4.4e-07
MMI174 G1 SEL N_8 VSS N_18_G2 l=1.8e-07 w=4.4e-07
MMI_160 RL CKB1 MPW VSS N_18_G2 l=1.8e-07 w=4.4e-07
MMI_89 G1 CKB1 G2 VSS N_18_G2 l=1.8e-07 w=4.4e-07
MMI_161 G3 CK1 RL VSS N_18_G2 l=1.8e-07 w=7.6e-07
MMI_162 G2 CK1 G4 VSS N_18_G2 l=1.8e-07 w=4.4e-07
XG17 SB G2 G3 DECAP_NAND2_G15
XG18 RB G3 G4 DECAP_NAND2_G16
XG19 RB RL QB1 DECAP_NAND2_G17
XG20 SB QB1 MPW DECAP_NAND2_G18
XG21 SEL SELB DECAP_INV_G19
XG22 CKB CK1 DECAP_INV_G19
XG23 CK1 CKB1 DECAP_INV_G19
XG24 QB1 Q DECAP_INV_G20
XG25 MPW QB DECAP_INV_G20
.ENDS

*******************************************************************************
* Main Circuit Netlist:                                                       *
*                            21                                                 *
* Block: HC8_SfrSp_DW01_dec_0                                                          *
* Last Time Saved: Dec 19 09:16:36 2006                                       *
*******************************************************************************

.SUBCKT HC8_SfrSp_DW01_dec_0 A[7]  A[6]  A[5]  A[4]  A[3]  A[2]  A[1]  A[0]  SUM[7]  SUM[6]  SUM[5]  SUM[4]  SUM[3]  SUM[2]  SUM[1]  SUM[0]  VDD  VSS  
XU1_B_3 carry_4_ A[3] carry_3_ VDD VSS OR2
XU1_B_4 carry_5_ A[4] carry_4_ VDD VSS OR2
XU1_B_5 carry_6_ A[5] carry_5_ VDD VSS OR2
XU1_B_2 carry_3_ A[2] carry_2_ VDD VSS OR2
XU1_B_1 carry_2_ A[1] A[0] VDD VSS OR2
XU1_A_3 SUM[3] A[3] carry_3_ VDD VSS XNR2
XU1_A_4 SUM[4] A[4] carry_4_ VDD VSS XNR2
XU1_A_5 SUM[5] A[5] carry_5_ VDD VSS XNR2
XU1_A_6 SUM[6] A[6] carry_6_ VDD VSS XNR2
XU1_A_1 SUM[1] A[1] A[0] VDD VSS XNR2
XU1_A_2 SUM[2] A[2] carry_2_ VDD VSS XNR2
XU6 SUM[7] A[7] n5 VDD VSS XOR2
XU7 n5 A[6] carry_6_ VDD VSS NR2
XU8 SUM[0] A[0] VDD VSS INV1
.ENDS

*******************************************************************************
* Main Circuit Netlist:                                                       *
*                            22                                                 *
* Block: HC8_SfrSp                                                          *
* Last Time Saved: Dec 19 09:16:36 2006                                       *
*******************************************************************************

.SUBCKT HC8_SfrSp SysRst_n  SysClk  SfrAddr[7]  SfrAddr[6]  SfrAddr[5]  SfrAddr[4]  SfrAddr[3]  SfrAddr[2]  SfrAddr[1]  SfrAddr[0]  SfrDataIn[7]  SfrDataIn[6]  SfrDataIn[5]  SfrDataIn[4]  SfrDataIn[3]  SfrDataIn[2]  SfrDataIn[1]  SfrDataIn[0]  SfrWr  SpInc  SpDec  SpDataOut[7]  SpDataOut[6]  SpDataOut[5]  SpDataOut[4]  SpDataOut[3]  SpDataOut[2]  SpDataOut[1]  SpDataOut[0]  SysClk__L3_N55  VDD  VSS  
XSpDataOut_reg_0_ SpDataOut[0] XSpDataOut_reg_0_/QB n58 SysClk__L3_N55 n2 VDD VSS DFFSBN
XSpDataOut_reg_1_ SpDataOut[1] XSpDataOut_reg_1_/QB n56 SysClk n2 VDD VSS DFFSBN
XSpDataOut_reg_2_ SpDataOut[2] XSpDataOut_reg_2_/QB n55 SysClk n2 VDD VSS DFFSBN
XU3 n51 SpDataOut[6] n40 SfrDataIn[6] n41 n21 n42 n12 n1 VDD VSS AO2222
XU4 n52 SpDataOut[5] n40 SfrDataIn[5] n41 n20 n42 n37 n1 VDD VSS AO2222
XU5 n53 SpDataOut[4] n40 SfrDataIn[4] n41 n19 n42 n11 n1 VDD VSS AO2222
XU6 n54 SpDataOut[3] n40 SfrDataIn[3] n41 n18 n42 n10 n1 VDD VSS AO2222
XU7 n55 SpDataOut[2] n40 SfrDataIn[2] n41 n17 n42 n9 n1 VDD VSS AO2222
XU8 n56 SpDataOut[1] n40 SfrDataIn[1] n41 n16 n42 n8 n1 VDD VSS AO2222
XU9 n57 SpDataOut[7] n40 SfrDataIn[7] n41 n22 n42 n13 n1 VDD VSS AO2222
XU10 n58 SpDataOut[0] n40 SfrDataIn[0] n41 n15 n42 n7 n1 VDD VSS AO2222
XU15 n44 n45 n46 n47 VDD VSS AN3
XU16 n47 SfrWr SfrAddr[7] SfrAddr[0] SfrAddr[1] VDD VSS AN4B1
XU12 n43 SpDec VDD VSS INV2
Xsub_593 SpDataOut[7] SpDataOut[6] SpDataOut[5] SpDataOut[4] SpDataOut[3] SpDataOut[2] SpDataOut[1] SpDataOut[0] n22 n21 n20 n19 n18 n17 n16 n15 VDD VSS HC8_SfrSp_DW01_dec_0
Xadd_591 SpDataOut[7] SpDataOut[6] SpDataOut[5] SpDataOut[4] SpDataOut[3] SpDataOut[2] SpDataOut[1] SpDataOut[0] n13 n12 n37 n11 n10 n9 n8 n7 VDD VSS HC8_SfrSp_DW01_inc_0
XSpDataOut_reg_7_ SpDataOut[7] n57 SysClk__L3_N55 n2 VDD VSS QDFFRBN
XSpDataOut_reg_6_ SpDataOut[6] n51 SysClk__L3_N55 n2 VDD VSS QDFFRBN
XSpDataOut_reg_5_ SpDataOut[5] n52 SysClk__L3_N55 n2 VDD VSS QDFFRBN
XSpDataOut_reg_3_ SpDataOut[3] n54 SysClk__L3_N55 n2 VDD VSS QDFFRBN
XSpDataOut_reg_4_ SpDataOut[4] n53 SysClk__L3_N55 n2 VDD VSS QDFFRBN
XU11 n42 n43 n1 VDD VSS NR2
XU13 n41 SpDec n1 n40 VDD VSS NR3
XU14 n1 SpInc VDD VSS BUF1
XU17 n2 SysRst_n VDD VSS BUF1
XU18 n40 SpDec SpInc n44 VDD VSS NR3
XU19 n46 SfrAddr[4] SfrAddr[6] SfrAddr[5] VDD VSS NR3
XU20 n45 SfrAddr[3] SfrAddr[2] VDD VSS NR2
.ENDS

*******************************************************************************
* Main Circuit Netlist:                                                       *
*                            23                                                 *
* Block: CIU192_Core                                                          *
* Last Time Saved: Dec 19 09:16:36 2006                                       *
*******************************************************************************

.SUBCKT CIU192_Core EXTCORE_Rst_n  EXTCORE_Clk  EXTCORE_Data  COREEXT_Data  VPP  VNN  EXTCORE_TpIn  EXTCORE_TpClk  EXTCORE_PORBypass_n  EXTCORE_PORIn_n  EXTCORE_FDBypass_n  EXTCORE_VDBypass_n  COREEXT_TpOut  COREEXT_POROut  COREEXT_FDH  COREEXT_FDL  COREEXT_FDOUT  COREEXT_VDREG  COREEXT_VD15  COREEXT_VD33  COREEXT_VD36  COREEXT_OSCOut  VBG06  VBG11  VDD  VCC  VSS  VDD  VCC  VSS  
XU8_BG VBG06 VBG11 IB IB1A IB2A IB1B IB2B ESFRCPU_IntVect_7_ VCC VSS STCEF018BG0615
XU9_REG IB1B IB2B IB1A IB2A VBG06 ESFRVR_Psb VDD VCC VSS STCEF018REG18_10
XU10_POR COREEXT_POROut VDD VSS STCEF018POR
XU11_VD VDD COREEXT_VDREG VBG11 IB1 IB2 IB7 ESFRVD_Pd COREEXT_VD36 COREEXT_VD33 XU11_VD/VD18 COREEXT_VD15 VDD VSS VCC VSS STCEF018VD1833_1536
XU12_FD EXTCORE_Clk VBG11 IB ESFRFD_Pd RSTFD_RS COREEXT_FDOUT COREEXT_FDH COREEXT_FDL IB1 IB2 IB7 VDD VSS VCC VSS STCEF018FD7K9M
XU_OscClk_1 net_OscClk CKMUESFR_OscClk_20M VDD VSS BUF4
XU_OscClk_2 COREEXT_OSCOut net_OscClk VDD VSS BUF8
XU1_CPU n3 SysClk__L3_N1 CPURAM_Addr[7] CPURAM_Addr[6] CPURAM_Addr[5] CPURAM_Addr[4] CPURAM_Addr[3] CPURAM_Addr[2] CPURAM_Addr[1] CPURAM_Addr[0] CPURAM_Cs_n CPURAM_Rd_n CPURAM_Wr_n CPURAM_Data[7] CPURAM_Data[6] CPURAM_Data[5] CPURAM_Data[4] CPURAM_Data[3] CPURAM_Data[2] CPURAM_Data[1] CPURAM_Data[0] RAMCPU_Data[7] RAMCPU_Data[6] RAMCPU_Data[5] RAMCPU_Data[4] RAMCPU_Data[3] RAMCPU_Data[2] RAMCPU_Data[1] RAMCPU_Data[0] CPUEMEM_Addr[15] CPUEMEM_Addr[14] CPUEMEM_Addr[13] CPUEMEM_Addr[12] CPUEMEM_Addr[11] CPUEMEM_Addr[10] CPUEMEM_Addr[9] CPUEMEM_Addr[8] CPUEMEM_Addr[7] CPUEMEM_Addr[6] CPUEMEM_Addr[5] CPUEMEM_Addr[4] CPUEMEM_Addr[3] CPUEMEM_Addr[2] CPUEMEM_Addr[1] CPUEMEM_Addr[0] CPUEMEM_Data[7] CPUEMEM_Data[6] CPUEMEM_Data[5] CPUEMEM_Data[4] CPUEMEM_Data[3] CPUEMEM_Data[2] CPUEMEM_Data[1] CPUEMEM_Data[0] CPUEMEM_PsCs_n CPUEMEM_PsRd_n CPUEMEM_PsWr_n CPUXRAM_Cs_n CPUXRAM_Rd_n CPUXRAM_Wr_n SYNOPSYS_UNCONNECTED_1 TSTCPU_ProgData[7] TSTCPU_ProgData[6] TSTCPU_ProgData[5] TSTCPU_ProgData[4] TSTCPU_ProgData[3] TSTCPU_ProgData[2] TSTCPU_ProgData[1] TSTCPU_ProgData[0] XRAMCPU_Data[7] XRAMCPU_Data[6] XRAMCPU_Data[5] XRAMCPU_Data[4] XRAMCPU_Data[3] XRAMCPU_Data[2] XRAMCPU_Data[1] XRAMCPU_Data[0] ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ net2 CPUESFR_BusAddr[7] CPUESFR_BusAddr[6] CPUESFR_BusAddr[5] CPUESFR_BusAddr[4] CPUESFR_BusAddr[3] CPUESFR_BusAddr[2] CPUESFR_BusAddr[1] CPUESFR_BusAddr[0] CPUESFR_BusData[7] CPUESFR_BusData[6] CPUESFR_BusData[5] CPUESFR_BusData[4] CPUESFR_BusData[3] CPUESFR_BusData[2] CPUESFR_BusData[1] CPUESFR_BusData[0] CPUESFR_BusWr ESFRCPU_BusData[7] ESFRCPU_BusData[6] ESFRCPU_BusData[5] ESFRCPU_BusData[4] ESFRCPU_BusData[3] ESFRCPU_BusData[2] ESFRCPU_BusData[1] ESFRCPU_BusData[0] ESFRCPU_IntReq ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect[5] ESFRCPU_IntVect[4] ESFRCPU_IntVect[3] ESFRCPU_IntVect_7_ ESFRCPU_IntVect[1] ESFRCPU_IntVect[0] CPUESFR_IntAck_r CPUESFR_Reti ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ SYNOPSYS_UNCONNECTED_2 SYNOPSYS_UNCONNECTED_3 ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ CPUEXT_IrData[23] CPUEXT_IrData[22] CPUEXT_IrData[21] CPUEXT_IrData[20] CPUEXT_IrData[19] CPUEXT_IrData[18] CPUEXT_IrData[17] CPUEXT_IrData[16] CPUEXT_IrData[15] CPUEXT_IrData[14] CPUEXT_IrData[13] CPUEXT_IrData[12] CPUEXT_IrData[11] CPUEXT_IrData[10] CPUEXT_IrData[9] CPUEXT_IrData[8] CPUEXT_IrData[7] CPUEXT_IrData[6] CPUEXT_IrData[5] CPUEXT_IrData[4] CPUEXT_IrData[3] CPUEXT_IrData[2] CPUEXT_IrData[1] CPUEXT_IrData[0] SYNOPSYS_UNCONNECTED_4 SYNOPSYS_UNCONNECTED_5 SYNOPSYS_UNCONNECTED_6 SYNOPSYS_UNCONNECTED_7 SYNOPSYS_UNCONNECTED_8 SYNOPSYS_UNCONNECTED_9 SYNOPSYS_UNCONNECTED_10 SYNOPSYS_UNCONNECTED_11 SYNOPSYS_UNCONNECTED_12 SYNOPSYS_UNCONNECTED_13 SYNOPSYS_UNCONNECTED_14 SYNOPSYS_UNCONNECTED_15 SYNOPSYS_UNCONNECTED_16 SYNOPSYS_UNCONNECTED_17 SYNOPSYS_UNCONNECTED_18 SYNOPSYS_UNCONNECTED_19 CPUTST_AccData[7] CPUTST_AccData[6] CPUTST_AccData[5] CPUTST_AccData[4] CPUTST_AccData[3] CPUTST_AccData[2] CPUTST_AccData[1] CPUTST_AccData[0] SYNOPSYS_UNCONNECTED_20 SYNOPSYS_UNCONNECTED_21 SYNOPSYS_UNCONNECTED_22 SYNOPSYS_UNCONNECTED_23 SYNOPSYS_UNCONNECTED_24 SYNOPSYS_UNCONNECTED_25 SYNOPSYS_UNCONNECTED_26 SYNOPSYS_UNCONNECTED_27 SYNOPSYS_UNCONNECTED_28 SYNOPSYS_UNCONNECTED_29 SYNOPSYS_UNCONNECTED_30 SYNOPSYS_UNCONNECTED_31 SYNOPSYS_UNCONNECTED_32 SYNOPSYS_UNCONNECTED_33 SYNOPSYS_UNCONNECTED_34 SYNOPSYS_UNCONNECTED_35 SYNOPSYS_UNCONNECTED_36 SYNOPSYS_UNCONNECTED_37 SYNOPSYS_UNCONNECTED_38 SYNOPSYS_UNCONNECTED_39 SYNOPSYS_UNCONNECTED_40 SYNOPSYS_UNCONNECTED_41 SYNOPSYS_UNCONNECTED_42 SYNOPSYS_UNCONNECTED_43 SYNOPSYS_UNCONNECTED_44 SYNOPSYS_UNCONNECTED_45 SYNOPSYS_UNCONNECTED_46 SYNOPSYS_UNCONNECTED_47 SYNOPSYS_UNCONNECTED_48 SYNOPSYS_UNCONNECTED_49 SYNOPSYS_UNCONNECTED_50 SYNOPSYS_UNCONNECTED_51 SYNOPSYS_UNCONNECTED_52 SYNOPSYS_UNCONNECTED_53 SYNOPSYS_UNCONNECTED_54 SYNOPSYS_UNCONNECTED_55 SYNOPSYS_UNCONNECTED_56 SYNOPSYS_UNCONNECTED_57 SYNOPSYS_UNCONNECTED_58 SYNOPSYS_UNCONNECTED_59 CPUEXT_CurState[1] CPUEXT_CurState[0] SysClk__L3_N10 SysClk__L3_N12 SysClk__L3_N16 SysClk__L3_N17 SysClk__L3_N19 SysClk__L3_N2 SysClk__L3_N21 SysClk__L3_N23 SysClk__L3_N25 SysClk__L3_N26 SysClk__L3_N29 SysClk__L3_N3 SysClk__L3_N30 SysClk__L3_N31 SysClk__L3_N33 SysClk__L3_N34 SysClk__L3_N37 SysClk__L3_N38 SysClk__L3_N39 SysClk__L3_N4 SysClk__L3_N40 SysClk__L3_N45 SysClk__L3_N46 SysClk__L3_N48 SysClk__L3_N49 SysClk__L3_N53 SysClk__L3_N54 SysClk__L3_N55 SysClk__L3_N56 SysClk__L3_N59 SysClk__L3_N6 SysClk__L3_N7 SysClk__L3_N70 SysClk__L3_N73 SysClk__L3_N74 SysClk__L3_N76 VDD VSS HC8_CPU
XU2_RAM n4 SysClk__L3_N0 CPURAM_Addr[7] CPURAM_Addr[6] CPURAM_Addr[5] CPURAM_Addr[4] CPURAM_Addr[3] CPURAM_Addr[2] CPURAM_Addr[1] CPURAM_Addr[0] CPURAM_Cs_n CPURAM_Rd_n CPURAM_Wr_n CPURAM_Data[7] CPURAM_Data[6] CPURAM_Data[5] CPURAM_Data[4] CPURAM_Data[3] CPURAM_Data[2] CPURAM_Data[1] CPURAM_Data[0] RAMCPU_Data[7] RAMCPU_Data[6] RAMCPU_Data[5] RAMCPU_Data[4] RAMCPU_Data[3] RAMCPU_Data[2] RAMCPU_Data[1] RAMCPU_Data[0] CPUEMEM_Addr[15] CPUEMEM_Addr[14] CPUEMEM_Addr[13] CPUEMEM_Addr[12] CPUEMEM_Addr[11] CPUEMEM_Addr[10] CPUEMEM_Addr[9] CPUEMEM_Addr[8] CPUEMEM_Addr[7] CPUEMEM_Addr[6] CPUEMEM_Addr[5] CPUEMEM_Addr[4] CPUEMEM_Addr[3] CPUEMEM_Addr[2] CPUEMEM_Addr[1] CPUEMEM_Addr[0] CPUEMEM_Data[7] CPUEMEM_Data[6] CPUEMEM_Data[5] CPUEMEM_Data[4] CPUEMEM_Data[3] CPUEMEM_Data[2] CPUEMEM_Data[1] CPUEMEM_Data[0] CPUXRAM_Cs_n CPUXRAM_Rd_n CPUXRAM_Wr_n XRAMCPU_Data[7] XRAMCPU_Data[6] XRAMCPU_Data[5] XRAMCPU_Data[4] XRAMCPU_Data[3] XRAMCPU_Data[2] XRAMCPU_Data[1] XRAMCPU_Data[0] ESFRMEM_StandbyEn SysClk__L3_N1 SysClk__L3_N10 SysClk__L3_N21 SysClk__L3_N23 SysClk__L3_N26 SysClk__L3_N31 SysClk__L3_N33 SysClk__L3_N34 SysClk__L3_N9 VDD VSS CIU192_RAM
XU3_FLS n4 SysClk__L3_N4 CPUEMEM_Addr[15] CPUEMEM_Addr[14] CPUEMEM_Addr[13] CPUEMEM_Addr[12] CPUEMEM_Addr[11] CPUEMEM_Addr[10] CPUEMEM_Addr[9] CPUEMEM_Addr[8] CPUEMEM_Addr[7] CPUEMEM_Addr[6] CPUEMEM_Addr[5] CPUEMEM_Addr[4] CPUEMEM_Addr[3] CPUEMEM_Addr[2] CPUEMEM_Addr[1] CPUEMEM_Addr[0] CPUEMEM_Data[7] CPUEMEM_Data[6] CPUEMEM_Data[5] CPUEMEM_Data[4] CPUEMEM_Data[3] CPUEMEM_Data[2] CPUEMEM_Data[1] CPUEMEM_Data[0] CPUEMEM_PsCs_n CPUEMEM_PsRd_n CPUEMEM_PsWr_n CPUEXT_IrData[23] CPUEXT_IrData[22] CPUEXT_IrData[21] CPUEXT_IrData[20] CPUEXT_IrData[19] CPUEXT_IrData[18] CPUEXT_IrData[17] CPUEXT_IrData[16] CPUEXT_IrData[15] CPUEXT_IrData[14] CPUEXT_IrData[13] CPUEXT_IrData[12] CPUEXT_IrData[11] CPUEXT_IrData[10] CPUEXT_IrData[9] CPUEXT_IrData[8] CPUEXT_IrData[7] CPUEXT_IrData[6] CPUEXT_IrData[5] CPUEXT_IrData[4] CPUEXT_IrData[3] CPUEXT_IrData[2] CPUEXT_IrData[1] CPUEXT_IrData[0] CPUEXT_CurState[1] CPUEXT_CurState[0] ESFRMEM_StandbyEn ESFRFLS_NvrSel ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRCPU_IntVect_7_ ESFRFLS_Bsr[2] ESFRFLS_Bsr[1] ESFRFLS_Bsr[0] ESFRFLS_OSCEN CKMUESFR_SciClk__L2_N1 FLSCKMU_HoldEn FLSCKMU_OscClk_20M RSTFLS_SysRstFin RSTFLS_Rst_n FLSTST_Data[15] FLSTST_Data[14] FLSTST_Data[13] FLSTST_Data[12] FLSTST_Data[11] FLSTST_Data[10] FLSTST_Data[9] FLSTST_Data[8] FLSTST_Data[7] FLSTST_Data[6] FLSTST_Data[5] FLSTST_Data[4] FLSTST_Data[3] FLSTST_Data[2] FLSTST_Data[1] FLSTST_Data[0] FLSTST_TBIT TSTFLS_Data[15] TSTFLS_Data[14] TSTFLS_Data[13] TSTFLS_Data[12] TSTFLS_Data[11] TSTFLS_Data[10] TSTFLS_Data[9] TSTFLS_Data[8] TSTFLS_Data[7] TSTFLS_Data[6] TSTFLS_Data[5] TSTFLS_Data[4] TSTFLS_Data[3] TSTFLS_Data[2] TSTFLS_Data[1] TSTFLS_Data[0] TSTFLS_Addr[17] TSTFLS_Addr[16] TSTFLS_Addr[15] TSTFLS_Addr[14] TSTFLS_Addr[13] TSTFLS_Addr[12] TSTFLS_Addr[11] TSTFLS_Addr[10] TSTFLS_Addr[9] TSTFLS_Addr[8] TSTFLS_Addr[7] TSTFLS_Addr[6] TSTFLS_Addr[5] TSTFLS_Addr[4] TSTFLS_Addr[3] TSTFLS_Addr[2] TSTFLS_Addr[1] TSTFLS_Addr[0] TSTFLS_IFREN TSTFLS_FlsRstb TSTFLS_BYTE TSTFLS_CS TSTFLS_OE TSTFLS_NVSTR TSTFLS_PROG TSTFLS_SERA TSTFLS_MASE TSTFLS_TME TSTFLS_TMR TSTFLS_FlsTestEn FLSTST_ProgData[7] FLSTST_ProgData[6] FLSTST_ProgData[5] FLSTST_ProgData[4] FLSTST_ProgData[3] FLSTST_ProgData[2] FLSTST_ProgData[1] FLSTST_ProgData[0] VPP VNN VDD VSS SysClk__L3_N5 SysClk__L3_N8 VDD VSS CIU192_FLS
XU4_CKMU EXTCORE_Clk RSTCKMU_RstFin n4 CKMURST_Clk ESFRCKMU_StandbyEn ESFRCKMU_Ckcon[0] SYNOPSYS_UNCONNECTED_60 CKMUESFR_SciClk CKMUESFR_OscClk_20M TSTCKMU_FuncTestEn CKMUTST_Clk FLSCKMU_OscClk_20M FLSCKMU_HoldEn SysClk CKMUESFR_OscClk_20M__L3_N0 VDD VSS CIU192_CKMU
XU5_RST n2 EXTCORE_PORBypass_n EXTCORE_PORIn_n EXTCORE_FDBypass_n EXTCORE_VDBypass_n CKMURST_Clk__L7_N0 RSTCKMU_RstFin n1 COREEXT_VD15 COREEXT_VD33 COREEXT_VD36 COREEXT_VDREG COREEXT_FDL COREEXT_FDH RSTFD_RS RSTFLS_Rst_n RSTFLS_SysRstFin ESFRFD_Pd ESFRVD_Pd RSTESFR_Fdout RSTESFR_Vdout RSTTST_PorRst_n SysRst_n CKMURST_Clk__L7_N1 CKMURST_Clk__L7_N2 CKMURST_Clk__L7_N3 VDD VSS CIU192_RST
XU6_ESFR n3 SysClk CPUESFR_BusAddr[7] CPUESFR_BusAddr[6] CPUESFR_BusAddr[5] CPUESFR_BusAddr[4] CPUESFR_BusAddr[3] CPUESFR_BusAddr[2] CPUESFR_BusAddr[1] CPUESFR_BusAddr[0] CPUESFR_BusData[7] CPUESFR_BusData[6] CPUESFR_BusData[5] CPUESFR_BusData[4] CPUESFR_BusData[3] CPUESFR_BusData[2] CPUESFR_BusData[1] CPUESFR_BusData[0] CPUESFR_BusWr ESFRCPU_BusData[7] ESFRCPU_BusData[6] ESFRCPU_BusData[5] ESFRCPU_BusData[4] ESFRCPU_BusData[3] ESFRCPU_BusData[2] ESFRCPU_BusData[1] ESFRCPU_BusData[0] ESFRCPU_IntReq CPUESFR_IntAck_r CPUESFR_Reti SYNOPSYS_UNCONNECTED_61 SYNOPSYS_UNCONNECTED_62 ESFRCPU_IntVect[5] ESFRCPU_IntVect[4] ESFRCPU_IntVect[3] SYNOPSYS_UNCONNECTED_63 ESFRCPU_IntVect[1] ESFRCPU_IntVect[0] CPURAM_Cs_n n2 EXTCORE_Data CKMUESFR_SciClk__L2_N0 EXTCORE_Clk CKMUESFR_OscClk_20M__L13_N0 ESFRCKMU_StandbyEn SYNOPSYS_UNCONNECTED_64 SYNOPSYS_UNCONNECTED_65 SYNOPSYS_UNCONNECTED_66 SYNOPSYS_UNCONNECTED_67 SYNOPSYS_UNCONNECTED_68 SYNOPSYS_UNCONNECTED_69 SYNOPSYS_UNCONNECTED_70 ESFRCKMU_Ckcon[0] COREEXT_POROut RSTESFR_Vdout RSTESFR_Fdout ESFRFD_Pd ESFRVD_Pd ESFRVR_Psb ESFRFLS_OSCEN ESFRMEM_StandbyEn ESFRFLS_NvrSel SYNOPSYS_UNCONNECTED_71 SYNOPSYS_UNCONNECTED_72 SYNOPSYS_UNCONNECTED_73 SYNOPSYS_UNCONNECTED_74 SYNOPSYS_UNCONNECTED_75 SYNOPSYS_UNCONNECTED_76 SYNOPSYS_UNCONNECTED_77 ESFRFLS_Bsr[2] ESFRFLS_Bsr[1] ESFRFLS_Bsr[0] ESFRTST_SciData TSTESFR_ClrFTOE ESFRTST_FuncTstOutEn TSTESFR_VDTestEn TSTESFR_FDTestEn SysClk__L3_N11 SysClk__L3_N12 SysClk__L3_N13 SysClk__L3_N14 SysClk__L3_N15 SysClk__L3_N17 SysClk__L3_N18 SysClk__L3_N20 SysClk__L3_N22 SysClk__L3_N24 SysClk__L3_N27 SysClk__L3_N28 SysClk__L3_N32 SysClk__L3_N35 SysClk__L3_N36 SysClk__L3_N41 SysClk__L3_N42 SysClk__L3_N43 SysClk__L3_N44 SysClk__L3_N47 SysClk__L3_N49 SysClk__L3_N5 SysClk__L3_N50 SysClk__L3_N51 SysClk__L3_N52 SysClk__L3_N54 SysClk__L3_N57 SysClk__L3_N58 SysClk__L3_N60 SysClk__L3_N61 SysClk__L3_N62 SysClk__L3_N63 SysClk__L3_N64 SysClk__L3_N65 SysClk__L3_N66 SysClk__L3_N67 SysClk__L3_N68 SysClk__L3_N69 SysClk__L3_N71 SysClk__L3_N72 SysClk__L3_N74 SysClk__L3_N75 SysClk__L3_N76 SysClk__L3_N77 SysClk__L3_N78 SysClk__L3_N79 CKMUESFR_SciClk__L2_N2 CKMUESFR_SciClk__L2_N3 CKMUESFR_SciClk__L2_N4 CKMUESFR_SciClk__L2_N5 CKMUESFR_SciClk__L2_N6 VDD VSS CIU192_ESFR
XU7_TST EXTCORE_Data n2 COREEXT_Data EXTCORE_TpClk EXTCORE_TpIn COREEXT_TpOut RSTTST_PorRst_n CKMUTST_Clk TSTCKMU_FuncTestEn ESFRTST_SciData ESFRTST_FuncTstOutEn TSTESFR_ClrFTOE TSTESFR_VDTestEn TSTESFR_FDTestEn SysRst_n CPUTST_AccData[7] CPUTST_AccData[6] CPUTST_AccData[5] CPUTST_AccData[4] CPUTST_AccData[3] CPUTST_AccData[2] CPUTST_AccData[1] CPUTST_AccData[0] TSTCPU_ProgData[7] TSTCPU_ProgData[6] TSTCPU_ProgData[5] TSTCPU_ProgData[4] TSTCPU_ProgData[3] TSTCPU_ProgData[2] TSTCPU_ProgData[1] TSTCPU_ProgData[0] FLSTST_Data[15] FLSTST_Data[14] FLSTST_Data[13] FLSTST_Data[12] FLSTST_Data[11] FLSTST_Data[10] FLSTST_Data[9] FLSTST_Data[8] FLSTST_Data[7] FLSTST_Data[6] FLSTST_Data[5] FLSTST_Data[4] FLSTST_Data[3] FLSTST_Data[2] FLSTST_Data[1] FLSTST_Data[0] FLSTST_TBIT TSTFLS_Data[15] TSTFLS_Data[14] TSTFLS_Data[13] TSTFLS_Data[12] TSTFLS_Data[11] TSTFLS_Data[10] TSTFLS_Data[9] TSTFLS_Data[8] TSTFLS_Data[7] TSTFLS_Data[6] TSTFLS_Data[5] TSTFLS_Data[4] TSTFLS_Data[3] TSTFLS_Data[2] TSTFLS_Data[1] TSTFLS_Data[0] TSTFLS_Addr[17] TSTFLS_Addr[16] TSTFLS_Addr[15] TSTFLS_Addr[14] TSTFLS_Addr[13] TSTFLS_Addr[12] TSTFLS_Addr[11] TSTFLS_Addr[10] TSTFLS_Addr[9] TSTFLS_Addr[8] TSTFLS_Addr[7] TSTFLS_Addr[6] TSTFLS_Addr[5] TSTFLS_Addr[4] TSTFLS_Addr[3] TSTFLS_Addr[2] TSTFLS_Addr[1] TSTFLS_Addr[0] TSTFLS_IFREN TSTFLS_FlsRstb TSTFLS_BYTE TSTFLS_CS TSTFLS_OE TSTFLS_NVSTR TSTFLS_PROG TSTFLS_SERA TSTFLS_MASE TSTFLS_TME TSTFLS_TMR TSTFLS_FlsTestEn FLSTST_ProgData[7] FLSTST_ProgData[6] FLSTST_ProgData[5] FLSTST_ProgData[4] FLSTST_ProgData[3] FLSTST_ProgData[2] FLSTST_ProgData[1] FLSTST_ProgData[0] VDD VSS CIU192_TST
XU35_SPARECELL VDD VSS CIU192_SpareCell
XU1 n1 COREEXT_POROut VDD VSS BUF1
XU2 n3 SysRst_n VDD VSS BUF1
XU3 n2 EXTCORE_Rst_n VDD VSS BUF1
XU4 n4 SysRst_n VDD VSS BUF1
XU5 ESFRCPU_IntVect_7_ VDD VSS TIE0
XU6 net2 VDD VSS TIE1
XCKMUESFR_OscClk_20M__L13_I0 CKMUESFR_OscClk_20M__L13_N0 CKMUESFR_OscClk_20M__L12_N0 VDD VSS BUF4CK
XCKMUESFR_OscClk_20M__L12_I0 CKMUESFR_OscClk_20M__L12_N0 CKMUESFR_OscClk_20M__L11_N0 VDD VSS BUF4CK
XCKMUESFR_OscClk_20M__L11_I0 CKMUESFR_OscClk_20M__L11_N0 CKMUESFR_OscClk_20M__L10_N0 VDD VSS BUF4CK
XCKMUESFR_OscClk_20M__L10_I0 CKMUESFR_OscClk_20M__L10_N0 CKMUESFR_OscClk_20M__L9_N0 VDD VSS BUF4CK
XCKMUESFR_OscClk_20M__L9_I0 CKMUESFR_OscClk_20M__L9_N0 CKMUESFR_OscClk_20M__L8_N0 VDD VSS BUF4CK
XCKMUESFR_OscClk_20M__L8_I0 CKMUESFR_OscClk_20M__L8_N0 CKMUESFR_OscClk_20M__L7_N0 VDD VSS BUF4CK
XCKMUESFR_OscClk_20M__L7_I0 CKMUESFR_OscClk_20M__L7_N0 CKMUESFR_OscClk_20M__L6_N0 VDD VSS BUF4CK
XCKMUESFR_OscClk_20M__L6_I0 CKMUESFR_OscClk_20M__L6_N0 CKMUESFR_OscClk_20M__L5_N0 VDD VSS BUF2CK
XCKMUESFR_OscClk_20M__L5_I0 CKMUESFR_OscClk_20M__L5_N0 CKMUESFR_OscClk_20M__L4_N0 VDD VSS BUF2CK
XCKMUESFR_OscClk_20M__L4_I0 CKMUESFR_OscClk_20M__L4_N0 CKMUESFR_OscClk_20M__L3_N0 VDD VSS BUF6CK
XCKMUESFR_OscClk_20M__L3_I0 CKMUESFR_OscClk_20M__L3_N0 CKMUESFR_OscClk_20M__L2_N0 VDD VSS BUF3CK
XCKMUESFR_OscClk_20M__L2_I0 CKMUESFR_OscClk_20M__L2_N0 CKMUESFR_OscClk_20M__L1_N0 VDD VSS BUF12CK
XCKMUESFR_OscClk_20M__L1_I0 CKMUESFR_OscClk_20M__L1_N0 CKMUESFR_OscClk_20M VDD VSS BUF2CK
XCKMURST_Clk__L7_I3 CKMURST_Clk__L7_N3 CKMURST_Clk__L6_N0 VDD VSS BUF12CK
XCKMURST_Clk__L7_I2 CKMURST_Clk__L7_N2 CKMURST_Clk__L6_N0 VDD VSS BUF12CK
XCKMURST_Clk__L7_I1 CKMURST_Clk__L7_N1 CKMURST_Clk__L6_N0 VDD VSS BUF12CK
XCKMURST_Clk__L7_I0 CKMURST_Clk__L7_N0 CKMURST_Clk__L6_N0 VDD VSS BUF12CK
XCKMURST_Clk__L6_I0 CKMURST_Clk__L6_N0 CKMURST_Clk__L5_N0 VDD VSS BUF12CK
XCKMURST_Clk__L5_I0 CKMURST_Clk__L5_N0 CKMURST_Clk__L4_N0 VDD VSS BUF8CK
XCKMURST_Clk__L4_I0 CKMURST_Clk__L4_N0 CKMURST_Clk__L3_N0 VDD VSS BUF8CK
XCKMURST_Clk__L3_I0 CKMURST_Clk__L3_N0 CKMURST_Clk__L2_N0 VDD VSS BUF8CK
XCKMURST_Clk__L2_I0 CKMURST_Clk__L2_N0 CKMURST_Clk__L1_N0 VDD VSS BUF8CK
XCKMURST_Clk__L1_I0 CKMURST_Clk__L1_N0 CKMURST_Clk VDD VSS BUF12CK
XCKMUESFR_SciClk__L2_I6 CKMUESFR_SciClk__L2_N6 CKMUESFR_SciClk__L1_N0 VDD VSS BUF12CK
XCKMUESFR_SciClk__L2_I5 CKMUESFR_SciClk__L2_N5 CKMUESFR_SciClk__L1_N0 VDD VSS BUF12CK
XCKMUESFR_SciClk__L2_I4 CKMUESFR_SciClk__L2_N4 CKMUESFR_SciClk__L1_N0 VDD VSS BUF12CK
XCKMUESFR_SciClk__L2_I3 CKMUESFR_SciClk__L2_N3 CKMUESFR_SciClk__L1_N0 VDD VSS BUF12CK
XCKMUESFR_SciClk__L2_I2 CKMUESFR_SciClk__L2_N2 CKMUESFR_SciClk__L1_N0 VDD VSS BUF12CK
XCKMUESFR_SciClk__L2_I1 CKMUESFR_SciClk__L2_N1 CKMUESFR_SciClk__L1_N0 VDD VSS BUF12CK
XCKMUESFR_SciClk__L2_I0 CKMUESFR_SciClk__L2_N0 CKMUESFR_SciClk__L1_N0 VDD VSS BUF12CK
XCKMUESFR_SciClk__L1_I0 CKMUESFR_SciClk__L1_N0 CKMUESFR_SciClk VDD VSS BUF12CK
XSysClk__L3_I79 SysClk__L3_N79 SysClk__L2_N8 VDD VSS BUF12CK
XSysClk__L3_I78 SysClk__L3_N78 SysClk__L2_N8 VDD VSS BUF12CK
XSysClk__L3_I77 SysClk__L3_N77 SysClk__L2_N8 VDD VSS BUF12CK
XSysClk__L3_I76 SysClk__L3_N76 SysClk__L2_N8 VDD VSS BUF12CK
XSysClk__L3_I75 SysClk__L3_N75 SysClk__L2_N8 VDD VSS BUF12CK
XSysClk__L3_I74 SysClk__L3_N74 SysClk__L2_N8 VDD VSS BUF12CK
XSysClk__L3_I73 SysClk__L3_N73 SysClk__L2_N8 VDD VSS BUF12CK
XSysClk__L3_I72 SysClk__L3_N72 SysClk__L2_N8 VDD VSS BUF12CK
XSysClk__L3_I71 SysClk__L3_N71 SysClk__L2_N8 VDD VSS BUF12CK
XSysClk__L3_I70 SysClk__L3_N70 SysClk__L2_N8 VDD VSS BUF12CK
XSysClk__L3_I69 SysClk__L3_N69 SysClk__L2_N7 VDD VSS BUF12CK
XSysClk__L3_I68 SysClk__L3_N68 SysClk__L2_N7 VDD VSS BUF12CK
XSysClk__L3_I67 SysClk__L3_N67 SysClk__L2_N7 VDD VSS BUF12CK
XSysClk__L3_I66 SysClk__L3_N66 SysClk__L2_N7 VDD VSS BUF12CK
XSysClk__L3_I65 SysClk__L3_N65 SysClk__L2_N7 VDD VSS BUF12CK
XSysClk__L3_I64 SysClk__L3_N64 SysClk__L2_N7 VDD VSS BUF12CK
XSysClk__L3_I63 SysClk__L3_N63 SysClk__L2_N7 VDD VSS BUF12CK
XSysClk__L3_I62 SysClk__L3_N62 SysClk__L2_N7 VDD VSS BUF12CK
XSysClk__L3_I61 SysClk__L3_N61 SysClk__L2_N7 VDD VSS BUF12CK
XSysClk__L3_I60 SysClk__L3_N60 SysClk__L2_N7 VDD VSS BUF12CK
XSysClk__L3_I59 SysClk__L3_N59 SysClk__L2_N6 VDD VSS BUF12CK
XSysClk__L3_I58 SysClk__L3_N58 SysClk__L2_N6 VDD VSS BUF12CK
XSysClk__L3_I57 SysClk__L3_N57 SysClk__L2_N6 VDD VSS BUF12CK
XSysClk__L3_I56 SysClk__L3_N56 SysClk__L2_N6 VDD VSS BUF12CK
XSysClk__L3_I55 SysClk__L3_N55 SysClk__L2_N6 VDD VSS BUF12CK
XSysClk__L3_I54 SysClk__L3_N54 SysClk__L2_N6 VDD VSS BUF12CK
XSysClk__L3_I53 SysClk__L3_N53 SysClk__L2_N6 VDD VSS BUF6CK
XSysClk__L3_I52 SysClk__L3_N52 SysClk__L2_N6 VDD VSS BUF12CK
XSysClk__L3_I51 SysClk__L3_N51 SysClk__L2_N6 VDD VSS BUF12CK
XSysClk__L3_I50 SysClk__L3_N50 SysClk__L2_N6 VDD VSS BUF12CK
XSysClk__L3_I49 SysClk__L3_N49 SysClk__L2_N5 VDD VSS BUF12CK
XSysClk__L3_I48 SysClk__L3_N48 SysClk__L2_N5 VDD VSS BUF12CK
XSysClk__L3_I47 SysClk__L3_N47 SysClk__L2_N5 VDD VSS BUF12CK
XSysClk__L3_I46 SysClk__L3_N46 SysClk__L2_N5 VDD VSS BUF12CK
XSysClk__L3_I45 SysClk__L3_N45 SysClk__L2_N5 VDD VSS BUF12CK
XSysClk__L3_I44 SysClk__L3_N44 SysClk__L2_N5 VDD VSS BUF12CK
XSysClk__L3_I43 SysClk__L3_N43 SysClk__L2_N5 VDD VSS BUF12CK
XSysClk__L3_I42 SysClk__L3_N42 SysClk__L2_N5 VDD VSS BUF12CK
XSysClk__L3_I41 SysClk__L3_N41 SysClk__L2_N5 VDD VSS BUF12CK
XSysClk__L3_I40 SysClk__L3_N40 SysClk__L2_N5 VDD VSS BUF12CK
XSysClk__L3_I39 SysClk__L3_N39 SysClk__L2_N4 VDD VSS BUF12CK
XSysClk__L3_I38 SysClk__L3_N38 SysClk__L2_N4 VDD VSS BUF12CK
XSysClk__L3_I37 SysClk__L3_N37 SysClk__L2_N4 VDD VSS BUF12CK
XSysClk__L3_I36 SysClk__L3_N36 SysClk__L2_N4 VDD VSS BUF12CK
XSysClk__L3_I35 SysClk__L3_N35 SysClk__L2_N4 VDD VSS BUF12CK
XSysClk__L3_I34 SysClk__L3_N34 SysClk__L2_N4 VDD VSS BUF12CK
XSysClk__L3_I33 SysClk__L3_N33 SysClk__L2_N4 VDD VSS BUF12CK
XSysClk__L3_I32 SysClk__L3_N32 SysClk__L2_N4 VDD VSS BUF12CK
XSysClk__L3_I31 SysClk__L3_N31 SysClk__L2_N4 VDD VSS BUF12CK
XSysClk__L3_I30 SysClk__L3_N30 SysClk__L2_N3 VDD VSS BUF12CK
XSysClk__L3_I29 SysClk__L3_N29 SysClk__L2_N3 VDD VSS BUF12CK
XSysClk__L3_I28 SysClk__L3_N28 SysClk__L2_N3 VDD VSS BUF12CK
XSysClk__L3_I27 SysClk__L3_N27 SysClk__L2_N3 VDD VSS BUF12CK
XSysClk__L3_I26 SysClk__L3_N26 SysClk__L2_N3 VDD VSS BUF12CK
XSysClk__L3_I25 SysClk__L3_N25 SysClk__L2_N3 VDD VSS BUF12CK
XSysClk__L3_I24 SysClk__L3_N24 SysClk__L2_N3 VDD VSS BUF12CK
XSysClk__L3_I23 SysClk__L3_N23 SysClk__L2_N3 VDD VSS BUF12CK
XSysClk__L3_I22 SysClk__L3_N22 SysClk__L2_N3 VDD VSS BUF12CK
XSysClk__L3_I21 SysClk__L3_N21 SysClk__L2_N3 VDD VSS BUF12CK
XSysClk__L3_I20 SysClk__L3_N20 SysClk__L2_N2 VDD VSS BUF12CK
XSysClk__L3_I19 SysClk__L3_N19 SysClk__L2_N2 VDD VSS BUF12CK
XSysClk__L3_I18 SysClk__L3_N18 SysClk__L2_N2 VDD VSS BUF12CK
XSysClk__L3_I17 SysClk__L3_N17 SysClk__L2_N2 VDD VSS BUF12CK
XSysClk__L3_I16 SysClk__L3_N16 SysClk__L2_N2 VDD VSS BUF12CK
XSysClk__L3_I15 SysClk__L3_N15 SysClk__L2_N2 VDD VSS BUF12CK
XSysClk__L3_I14 SysClk__L3_N14 SysClk__L2_N2 VDD VSS BUF12CK
XSysClk__L3_I13 SysClk__L3_N13 SysClk__L2_N2 VDD VSS BUF12CK
XSysClk__L3_I12 SysClk__L3_N12 SysClk__L2_N2 VDD VSS BUF12CK
XSysClk__L3_I11 SysClk__L3_N11 SysClk__L2_N2 VDD VSS BUF12CK
XSysClk__L3_I10 SysClk__L3_N10 SysClk__L2_N2 VDD VSS BUF12CK
XSysClk__L3_I9 SysClk__L3_N9 SysClk__L2_N1 VDD VSS BUF12CK
XSysClk__L3_I8 SysClk__L3_N8 SysClk__L2_N0 VDD VSS BUF12CK
XSysClk__L3_I7 SysClk__L3_N7 SysClk__L2_N0 VDD VSS BUF12CK
XSysClk__L3_I6 SysClk__L3_N6 SysClk__L2_N0 VDD VSS BUF12CK
XSysClk__L3_I5 SysClk__L3_N5 SysClk__L2_N0 VDD VSS BUF12CK
XSysClk__L3_I4 SysClk__L3_N4 SysClk__L2_N0 VDD VSS BUF12CK
XSysClk__L3_I3 SysClk__L3_N3 SysClk__L2_N0 VDD VSS BUF12CK
XSysClk__L3_I2 SysClk__L3_N2 SysClk__L2_N0 VDD VSS BUF12CK
XSysClk__L3_I1 SysClk__L3_N1 SysClk__L2_N0 VDD VSS BUF12CK
XSysClk__L3_I0 SysClk__L3_N0 SysClk__L2_N0 VDD VSS BUF12CK
XSysClk__L2_I8 SysClk__L2_N8 SysClk__L1_N0 VDD VSS BUF12CK
XSysClk__L2_I7 SysClk__L2_N7 SysClk__L1_N0 VDD VSS BUF12CK
XSysClk__L2_I6 SysClk__L2_N6 SysClk__L1_N0 VDD VSS BUF12CK
XSysClk__L2_I5 SysClk__L2_N5 SysClk__L1_N0 VDD VSS BUF12CK
XSysClk__L2_I4 SysClk__L2_N4 SysClk__L1_N0 VDD VSS BUF12CK
XSysClk__L2_I3 SysClk__L2_N3 SysClk__L1_N0 VDD VSS BUF12CK
XSysClk__L2_I2 SysClk__L2_N2 SysClk__L1_N0 VDD VSS BUF12CK
XSysClk__L2_I1 SysClk__L2_N1 SysClk__L1_N0 VDD VSS BUF12CK
XSysClk__L2_I0 SysClk__L2_N0 SysClk__L1_N0 VDD VSS BUF12CK
XSysClk__L1_I0 SysClk__L1_N0 SysClk VDD VSS BUF12CK
.ENDS


*******************************************************************************
* Main Circuit Netlist:                                                       *
*                            24                                                 *
* Block: MIDC_7_VIRTUAL_C_VIRTUAL_C                                                        *
* Last Time Saved: Dec 19 09:16:36 2006                                       *
*******************************************************************************

.SUBCKT MIDC_7_VIRTUAL_C_VIRTUAL_C 177  178  179  180  181  182  183  184  185  186  187  188  189  190  191  192  193  194  195  196  197  198  199  200  201  202  203  204  205  206  207  208  669  671  672  673  675  677  679  680  681  685  687  688  689  692  693  695  696  697  700  701  703  704  705  707  708  709  711  712  713  717  719  720  721  724  725  726  727  728  729  730  731  732  733  734  735  736  737  738  739  740  741  742  743  744  745  766  767  768  769  770  771  772  773  774  775  776  1077  1078  1079  1080  1081  1082  1083  1084  1085  1086  1087  1088  1089  1090  1091  1092  1093  1094  1095  1096  1097  1098  1099  1100  1101  1102  1103  1104  1105  1106  1107  1108  1109  1110  1111  1112  1113  1114  1115  1116  1117  1118  1119  1120  1121  1122  1123  1124  1125  1126  1127  1128  1129  1130  1131  1132  1133  1134  1135  1136  1137  1138  1139  1140  1141  1142  1163  1164  1185  1186  1207  1208  1229  1230  1251  1252  1273  1274  1295  1296  1317  1318  1339  1340  1361  1362  1383  1384  1405  1406  1427  1428  1449  1450  1471  1472  1493  1494  1515  1516  1537  1538  1559  1560  1581  1582  1603  1604  1625  1626  1647  1648  1669  1670  1691  1692  1713  1714  1735  1736  1757  1758  1759  1760  1761  1762  1763  1764  1765  1766  1767  2388  2389  2390  2391  2392  2393  2394  2395  2396  2397  2398  2399  2400  2401  2402  2403  2404  2405  2406  2407  2408  2409  2410  
M0 177 1084 1082 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=3930
M1 177 1086 679 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=4800
M2 177 1094 1092 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=8930
M3 177 1096 687 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=9800
M4 177 1104 1102 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=13930
M5 177 1106 695 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=14800
M6 177 1114 1112 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=18930
M7 177 1116 703 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=19800
M8 177 1124 1122 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=23930
M9 177 1126 711 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=24800
M10 177 1134 1132 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=28930
M11 177 1136 719 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=29800
M12 177 1137 1077 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=33930
M13 177 1109 685 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=34800
M14 177 1123 1133 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=38930
M15 177 1113 709 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=39800
M16 177 1119 1083 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=43930
M17 177 1115 677 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=44800
M18 177 1135 1085 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=48930
M19 177 1099 708 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=230 $Y=49800
M20 178 1084 673 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=3930
M21 1088 1086 178 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=4790
M22 178 1094 681 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=8930
M23 1098 1096 178 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=9790
M24 178 1104 689 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=13930
M25 1108 1106 178 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=14790
M26 178 1114 697 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=18930
M27 1118 1116 178 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=19790
M28 178 1124 705 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=23930
M29 1128 1126 178 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=24790
M30 178 1134 713 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=28930
M31 1138 1136 178 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=29790
M32 178 1137 721 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=33930
M33 1129 1109 178 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=34790
M34 178 1123 717 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=38930
M35 1103 1113 178 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=39790
M36 178 1119 701 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=43930
M37 1125 1115 178 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=44790
M38 178 1135 669 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=48930
M39 1127 1099 178 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=760 $Y=49790
M40 180 1084 1176 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=3930
M41 180 1086 1165 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=4800
M42 180 1094 1177 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=8930
M43 180 1096 1166 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=9800
M44 180 1104 1178 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=13930
M45 180 1106 1167 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=14800
M46 180 1114 1179 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=18930
M47 180 1116 1168 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=19800
M48 180 1124 1180 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=23930
M49 180 1126 1169 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=24800
M50 180 1134 1181 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=28930
M51 180 1136 1170 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=29800
M52 180 1137 1182 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=33930
M53 180 1109 1171 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=34800
M54 180 1123 1183 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=38930
M55 180 1113 1172 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=39800
M56 180 1119 1184 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=43930
M57 180 1115 1173 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=44800
M58 180 1135 1175 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=48930
M59 180 1099 1174 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=2470 $Y=49800
M60 181 1084 1143 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=3930
M61 1144 1086 181 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=4790
M62 181 1094 1145 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=8930
M63 1146 1096 181 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=9790
M64 181 1104 1147 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=13930
M65 1148 1106 181 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=14790
M66 181 1114 1149 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=18930
M67 1150 1116 181 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=19790
M68 181 1124 1151 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=23930
M69 1152 1126 181 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=24790
M70 181 1134 1153 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=28930
M71 1154 1136 181 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=29790
M72 181 1137 1155 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=33930
M73 1156 1109 181 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=34790
M74 181 1123 1157 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=38930
M75 1158 1113 181 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=39790
M76 181 1119 1159 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=43930
M77 1160 1115 181 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=44790
M78 181 1135 1161 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=48930
M79 1162 1099 181 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=3000 $Y=49790
M80 182 1084 1220 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=3930
M81 182 1086 1209 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=4800
M82 182 1094 1221 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=8930
M83 182 1096 1210 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=9800
M84 182 1104 1222 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=13930
M85 182 1106 1211 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=14800
M86 182 1114 1223 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=18930
M87 182 1116 1212 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=19800
M88 182 1124 1224 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=23930
M89 182 1126 1213 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=24800
M90 182 1134 1225 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=28930
M91 182 1136 1214 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=29800
M92 182 1137 1226 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=33930
M93 182 1109 1215 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=34800
M94 182 1123 1227 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=38930
M95 182 1113 1216 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=39800
M96 182 1119 1228 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=43930
M97 182 1115 1217 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=44800
M98 182 1135 1219 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=48930
M99 182 1099 1218 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=4710 $Y=49800
M100 183 1084 1187 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=3930
M101 1188 1086 183 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=4790
M102 183 1094 1189 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=8930
M103 1190 1096 183 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=9790
M104 183 1104 1191 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=13930
M105 1192 1106 183 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=14790
M106 183 1114 1193 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=18930
M107 1194 1116 183 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=19790
M108 183 1124 1195 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=23930
M109 1196 1126 183 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=24790
M110 183 1134 1197 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=28930
M111 1198 1136 183 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=29790
M112 183 1137 1199 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=33930
M113 1200 1109 183 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=34790
M114 183 1123 1201 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=38930
M115 1202 1113 183 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=39790
M116 183 1119 1203 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=43930
M117 1204 1115 183 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=44790
M118 183 1135 1205 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=48930
M119 1206 1099 183 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=5240 $Y=49790
M120 184 1084 1264 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=3930
M121 184 1086 1253 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=4800
M122 184 1094 1265 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=8930
M123 184 1096 1254 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=9800
M124 184 1104 1266 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=13930
M125 184 1106 1255 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=14800
M126 184 1114 1267 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=18930
M127 184 1116 1256 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=19800
M128 184 1124 1268 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=23930
M129 184 1126 1257 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=24800
M130 184 1134 1269 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=28930
M131 184 1136 1258 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=29800
M132 184 1137 1270 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=33930
M133 184 1109 1259 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=34800
M134 184 1123 1271 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=38930
M135 184 1113 1260 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=39800
M136 184 1119 1272 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=43930
M137 184 1115 1261 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=44800
M138 184 1135 1263 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=48930
M139 184 1099 1262 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=6950 $Y=49800
M140 185 1084 1231 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=3930
M141 1232 1086 185 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=4790
M142 185 1094 1233 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=8930
M143 1234 1096 185 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=9790
M144 185 1104 1235 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=13930
M145 1236 1106 185 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=14790
M146 185 1114 1237 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=18930
M147 1238 1116 185 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=19790
M148 185 1124 1239 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=23930
M149 1240 1126 185 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=24790
M150 185 1134 1241 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=28930
M151 1242 1136 185 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=29790
M152 185 1137 1243 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=33930
M153 1244 1109 185 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=34790
M154 185 1123 1245 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=38930
M155 1246 1113 185 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=39790
M156 185 1119 1247 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=43930
M157 1248 1115 185 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=44790
M158 185 1135 1249 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=48930
M159 1250 1099 185 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=7480 $Y=49790
M160 186 1084 1308 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=3930
M161 186 1086 1297 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=4800
M162 186 1094 1309 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=8930
M163 186 1096 1298 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=9800
M164 186 1104 1310 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=13930
M165 186 1106 1299 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=14800
M166 186 1114 1311 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=18930
M167 186 1116 1300 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=19800
M168 186 1124 1312 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=23930
M169 186 1126 1301 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=24800
M170 186 1134 1313 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=28930
M171 186 1136 1302 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=29800
M172 186 1137 1314 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=33930
M173 186 1109 1303 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=34800
M174 186 1123 1315 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=38930
M175 186 1113 1304 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=39800
M176 186 1119 1316 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=43930
M177 186 1115 1305 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=44800
M178 186 1135 1307 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=48930
M179 186 1099 1306 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9190 $Y=49800
M180 187 1084 1275 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=3930
M181 1276 1086 187 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=4790
M182 187 1094 1277 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=8930
M183 1278 1096 187 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=9790
M184 187 1104 1279 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=13930
M185 1280 1106 187 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=14790
M186 187 1114 1281 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=18930
M187 1282 1116 187 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=19790
M188 187 1124 1283 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=23930
M189 1284 1126 187 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=24790
M190 187 1134 1285 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=28930
M191 1286 1136 187 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=29790
M192 187 1137 1287 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=33930
M193 1288 1109 187 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=34790
M194 187 1123 1289 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=38930
M195 1290 1113 187 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=39790
M196 187 1119 1291 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=43930
M197 1292 1115 187 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=44790
M198 187 1135 1293 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=48930
M199 1294 1099 187 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=9720 $Y=49790
M200 188 1084 1352 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=3930
M201 188 1086 1341 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=4800
M202 188 1094 1353 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=8930
M203 188 1096 1342 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=9800
M204 188 1104 1354 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=13930
M205 188 1106 1343 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=14800
M206 188 1114 1355 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=18930
M207 188 1116 1344 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=19800
M208 188 1124 1356 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=23930
M209 188 1126 1345 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=24800
M210 188 1134 1357 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=28930
M211 188 1136 1346 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=29800
M212 188 1137 1358 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=33930
M213 188 1109 1347 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=34800
M214 188 1123 1359 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=38930
M215 188 1113 1348 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=39800
M216 188 1119 1360 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=43930
M217 188 1115 1349 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=44800
M218 188 1135 1351 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=48930
M219 188 1099 1350 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11430 $Y=49800
M220 189 1084 1319 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=3930
M221 1320 1086 189 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=4790
M222 189 1094 1321 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=8930
M223 1322 1096 189 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=9790
M224 189 1104 1323 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=13930
M225 1324 1106 189 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=14790
M226 189 1114 1325 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=18930
M227 1326 1116 189 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=19790
M228 189 1124 1327 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=23930
M229 1328 1126 189 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=24790
M230 189 1134 1329 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=28930
M231 1330 1136 189 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=29790
M232 189 1137 1331 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=33930
M233 1332 1109 189 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=34790
M234 189 1123 1333 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=38930
M235 1334 1113 189 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=39790
M236 189 1119 1335 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=43930
M237 1336 1115 189 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=44790
M238 189 1135 1337 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=48930
M239 1338 1099 189 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=11960 $Y=49790
M240 190 1084 1396 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=3930
M241 190 1086 1385 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=4800
M242 190 1094 1397 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=8930
M243 190 1096 1386 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=9800
M244 190 1104 1398 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=13930
M245 190 1106 1387 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=14800
M246 190 1114 1399 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=18930
M247 190 1116 1388 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=19800
M248 190 1124 1400 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=23930
M249 190 1126 1389 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=24800
M250 190 1134 1401 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=28930
M251 190 1136 1390 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=29800
M252 190 1137 1402 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=33930
M253 190 1109 1391 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=34800
M254 190 1123 1403 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=38930
M255 190 1113 1392 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=39800
M256 190 1119 1404 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=43930
M257 190 1115 1393 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=44800
M258 190 1135 1395 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=48930
M259 190 1099 1394 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=13670 $Y=49800
M260 191 1084 1363 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=3930
M261 1364 1086 191 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=4790
M262 191 1094 1365 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=8930
M263 1366 1096 191 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=9790
M264 191 1104 1367 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=13930
M265 1368 1106 191 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=14790
M266 191 1114 1369 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=18930
M267 1370 1116 191 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=19790
M268 191 1124 1371 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=23930
M269 1372 1126 191 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=24790
M270 191 1134 1373 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=28930
M271 1374 1136 191 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=29790
M272 191 1137 1375 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=33930
M273 1376 1109 191 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=34790
M274 191 1123 1377 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=38930
M275 1378 1113 191 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=39790
M276 191 1119 1379 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=43930
M277 1380 1115 191 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=44790
M278 191 1135 1381 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=48930
M279 1382 1099 191 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=14200 $Y=49790
M280 192 1084 1440 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=3930
M281 192 1086 1429 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=4800
M282 192 1094 1441 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=8930
M283 192 1096 1430 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=9800
M284 192 1104 1442 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=13930
M285 192 1106 1431 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=14800
M286 192 1114 1443 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=18930
M287 192 1116 1432 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=19800
M288 192 1124 1444 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=23930
M289 192 1126 1433 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=24800
M290 192 1134 1445 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=28930
M291 192 1136 1434 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=29800
M292 192 1137 1446 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=33930
M293 192 1109 1435 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=34800
M294 192 1123 1447 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=38930
M295 192 1113 1436 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=39800
M296 192 1119 1448 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=43930
M297 192 1115 1437 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=44800
M298 192 1135 1439 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=48930
M299 192 1099 1438 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=15910 $Y=49800
M300 193 1084 1407 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=3930
M301 1408 1086 193 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=4790
M302 193 1094 1409 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=8930
M303 1410 1096 193 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=9790
M304 193 1104 1411 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=13930
M305 1412 1106 193 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=14790
M306 193 1114 1413 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=18930
M307 1414 1116 193 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=19790
M308 193 1124 1415 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=23930
M309 1416 1126 193 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=24790
M310 193 1134 1417 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=28930
M311 1418 1136 193 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=29790
M312 193 1137 1419 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=33930
M313 1420 1109 193 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=34790
M314 193 1123 1421 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=38930
M315 1422 1113 193 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=39790
M316 193 1119 1423 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=43930
M317 1424 1115 193 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=44790
M318 193 1135 1425 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=48930
M319 1426 1099 193 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=16440 $Y=49790
M320 194 1084 1484 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=3930
M321 194 1086 1473 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=4800
M322 194 1094 1485 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=8930
M323 194 1096 1474 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=9800
M324 194 1104 1486 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=13930
M325 194 1106 1475 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=14800
M326 194 1114 1487 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=18930
M327 194 1116 1476 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=19800
M328 194 1124 1488 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=23930
M329 194 1126 1477 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=24800
M330 194 1134 1489 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=28930
M331 194 1136 1478 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=29800
M332 194 1137 1490 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=33930
M333 194 1109 1479 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=34800
M334 194 1123 1491 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=38930
M335 194 1113 1480 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=39800
M336 194 1119 1492 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=43930
M337 194 1115 1481 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=44800
M338 194 1135 1483 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=48930
M339 194 1099 1482 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18150 $Y=49800
M340 195 1084 1451 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=3930
M341 1452 1086 195 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=4790
M342 195 1094 1453 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=8930
M343 1454 1096 195 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=9790
M344 195 1104 1455 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=13930
M345 1456 1106 195 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=14790
M346 195 1114 1457 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=18930
M347 1458 1116 195 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=19790
M348 195 1124 1459 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=23930
M349 1460 1126 195 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=24790
M350 195 1134 1461 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=28930
M351 1462 1136 195 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=29790
M352 195 1137 1463 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=33930
M353 1464 1109 195 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=34790
M354 195 1123 1465 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=38930
M355 1466 1113 195 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=39790
M356 195 1119 1467 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=43930
M357 1468 1115 195 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=44790
M358 195 1135 1469 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=48930
M359 1470 1099 195 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=18680 $Y=49790
M360 196 1084 1528 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=3930
M361 196 1086 1517 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=4800
M362 196 1094 1529 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=8930
M363 196 1096 1518 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=9800
M364 196 1104 1530 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=13930
M365 196 1106 1519 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=14800
M366 196 1114 1531 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=18930
M367 196 1116 1520 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=19800
M368 196 1124 1532 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=23930
M369 196 1126 1521 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=24800
M370 196 1134 1533 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=28930
M371 196 1136 1522 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=29800
M372 196 1137 1534 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=33930
M373 196 1109 1523 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=34800
M374 196 1123 1535 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=38930
M375 196 1113 1524 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=39800
M376 196 1119 1536 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=43930
M377 196 1115 1525 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=44800
M378 196 1135 1527 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=48930
M379 196 1099 1526 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20390 $Y=49800
M380 197 1084 1495 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=3930
M381 1496 1086 197 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=4790
M382 197 1094 1497 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=8930
M383 1498 1096 197 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=9790
M384 197 1104 1499 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=13930
M385 1500 1106 197 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=14790
M386 197 1114 1501 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=18930
M387 1502 1116 197 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=19790
M388 197 1124 1503 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=23930
M389 1504 1126 197 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=24790
M390 197 1134 1505 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=28930
M391 1506 1136 197 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=29790
M392 197 1137 1507 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=33930
M393 1508 1109 197 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=34790
M394 197 1123 1509 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=38930
M395 1510 1113 197 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=39790
M396 197 1119 1511 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=43930
M397 1512 1115 197 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=44790
M398 197 1135 1513 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=48930
M399 1514 1099 197 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=20920 $Y=49790
M400 198 1084 1572 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=3930
M401 198 1086 1561 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=4800
M402 198 1094 1573 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=8930
M403 198 1096 1562 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=9800
M404 198 1104 1574 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=13930
M405 198 1106 1563 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=14800
M406 198 1114 1575 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=18930
M407 198 1116 1564 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=19800
M408 198 1124 1576 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=23930
M409 198 1126 1565 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=24800
M410 198 1134 1577 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=28930
M411 198 1136 1566 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=29800
M412 198 1137 1578 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=33930
M413 198 1109 1567 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=34800
M414 198 1123 1579 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=38930
M415 198 1113 1568 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=39800
M416 198 1119 1580 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=43930
M417 198 1115 1569 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=44800
M418 198 1135 1571 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=48930
M419 198 1099 1570 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=22630 $Y=49800
M420 199 1084 1539 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=3930
M421 1540 1086 199 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=4790
M422 199 1094 1541 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=8930
M423 1542 1096 199 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=9790
M424 199 1104 1543 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=13930
M425 1544 1106 199 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=14790
M426 199 1114 1545 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=18930
M427 1546 1116 199 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=19790
M428 199 1124 1547 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=23930
M429 1548 1126 199 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=24790
M430 199 1134 1549 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=28930
M431 1550 1136 199 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=29790
M432 199 1137 1551 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=33930
M433 1552 1109 199 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=34790
M434 199 1123 1553 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=38930
M435 1554 1113 199 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=39790
M436 199 1119 1555 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=43930
M437 1556 1115 199 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=44790
M438 199 1135 1557 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=48930
M439 1558 1099 199 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=23160 $Y=49790
M440 200 1084 1616 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=3930
M441 200 1086 1605 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=4800
M442 200 1094 1617 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=8930
M443 200 1096 1606 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=9800
M444 200 1104 1618 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=13930
M445 200 1106 1607 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=14800
M446 200 1114 1619 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=18930
M447 200 1116 1608 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=19800
M448 200 1124 1620 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=23930
M449 200 1126 1609 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=24800
M450 200 1134 1621 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=28930
M451 200 1136 1610 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=29800
M452 200 1137 1622 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=33930
M453 200 1109 1611 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=34800
M454 200 1123 1623 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=38930
M455 200 1113 1612 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=39800
M456 200 1119 1624 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=43930
M457 200 1115 1613 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=44800
M458 200 1135 1615 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=48930
M459 200 1099 1614 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=24870 $Y=49800
M460 201 1084 1583 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=3930
M461 1584 1086 201 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=4790
M462 201 1094 1585 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=8930
M463 1586 1096 201 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=9790
M464 201 1104 1587 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=13930
M465 1588 1106 201 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=14790
M466 201 1114 1589 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=18930
M467 1590 1116 201 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=19790
M468 201 1124 1591 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=23930
M469 1592 1126 201 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=24790
M470 201 1134 1593 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=28930
M471 1594 1136 201 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=29790
M472 201 1137 1595 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=33930
M473 1596 1109 201 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=34790
M474 201 1123 1597 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=38930
M475 1598 1113 201 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=39790
M476 201 1119 1599 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=43930
M477 1600 1115 201 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=44790
M478 201 1135 1601 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=48930
M479 1602 1099 201 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=25400 $Y=49790
M480 202 1084 1660 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=3930
M481 202 1086 1649 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=4800
M482 202 1094 1661 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=8930
M483 202 1096 1650 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=9800
M484 202 1104 1662 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=13930
M485 202 1106 1651 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=14800
M486 202 1114 1663 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=18930
M487 202 1116 1652 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=19800
M488 202 1124 1664 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=23930
M489 202 1126 1653 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=24800
M490 202 1134 1665 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=28930
M491 202 1136 1654 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=29800
M492 202 1137 1666 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=33930
M493 202 1109 1655 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=34800
M494 202 1123 1667 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=38930
M495 202 1113 1656 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=39800
M496 202 1119 1668 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=43930
M497 202 1115 1657 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=44800
M498 202 1135 1659 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=48930
M499 202 1099 1658 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27110 $Y=49800
M500 203 1084 1627 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=3930
M501 1628 1086 203 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=4790
M502 203 1094 1629 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=8930
M503 1630 1096 203 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=9790
M504 203 1104 1631 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=13930
M505 1632 1106 203 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=14790
M506 203 1114 1633 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=18930
M507 1634 1116 203 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=19790
M508 203 1124 1635 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=23930
M509 1636 1126 203 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=24790
M510 203 1134 1637 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=28930
M511 1638 1136 203 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=29790
M512 203 1137 1639 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=33930
M513 1640 1109 203 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=34790
M514 203 1123 1641 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=38930
M515 1642 1113 203 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=39790
M516 203 1119 1643 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=43930
M517 1644 1115 203 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=44790
M518 203 1135 1645 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=48930
M519 1646 1099 203 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=27640 $Y=49790
M520 204 1084 1704 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=3930
M521 204 1086 1693 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=4800
M522 204 1094 1705 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=8930
M523 204 1096 1694 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=9800
M524 204 1104 1706 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=13930
M525 204 1106 1695 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=14800
M526 204 1114 1707 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=18930
M527 204 1116 1696 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=19800
M528 204 1124 1708 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=23930
M529 204 1126 1697 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=24800
M530 204 1134 1709 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=28930
M531 204 1136 1698 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=29800
M532 204 1137 1710 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=33930
M533 204 1109 1699 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=34800
M534 204 1123 1711 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=38930
M535 204 1113 1700 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=39800
M536 204 1119 1712 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=43930
M537 204 1115 1701 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=44800
M538 204 1135 1703 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=48930
M539 204 1099 1702 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29350 $Y=49800
M540 205 1084 1671 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=3930
M541 1672 1086 205 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=4790
M542 205 1094 1673 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=8930
M543 1674 1096 205 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=9790
M544 205 1104 1675 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=13930
M545 1676 1106 205 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=14790
M546 205 1114 1677 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=18930
M547 1678 1116 205 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=19790
M548 205 1124 1679 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=23930
M549 1680 1126 205 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=24790
M550 205 1134 1681 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=28930
M551 1682 1136 205 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=29790
M552 205 1137 1683 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=33930
M553 1684 1109 205 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=34790
M554 205 1123 1685 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=38930
M555 1686 1113 205 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=39790
M556 205 1119 1687 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=43930
M557 1688 1115 205 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=44790
M558 205 1135 1689 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=48930
M559 1690 1099 205 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=29880 $Y=49790
M560 206 1084 1748 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=3930
M561 206 1086 1737 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=4800
M562 206 1094 1749 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=8930
M563 206 1096 1738 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=9800
M564 206 1104 1750 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=13930
M565 206 1106 1739 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=14800
M566 206 1114 1751 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=18930
M567 206 1116 1740 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=19800
M568 206 1124 1752 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=23930
M569 206 1126 1741 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=24800
M570 206 1134 1753 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=28930
M571 206 1136 1742 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=29800
M572 206 1137 1754 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=33930
M573 206 1109 1743 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=34800
M574 206 1123 1755 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=38930
M575 206 1113 1744 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=39800
M576 206 1119 1756 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=43930
M577 206 1115 1745 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=44800
M578 206 1135 1747 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=48930
M579 206 1099 1746 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=31590 $Y=49800
M580 207 1084 1715 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=3930
M581 1716 1086 207 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=4790
M582 207 1094 1717 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=8930
M583 1718 1096 207 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=9790
M584 207 1104 1719 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=13930
M585 1720 1106 207 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=14790
M586 207 1114 1721 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=18930
M587 1722 1116 207 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=19790
M588 207 1124 1723 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=23930
M589 1724 1126 207 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=24790
M590 207 1134 1725 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=28930
M591 1726 1136 207 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=29790
M592 207 1137 1727 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=33930
M593 1728 1109 207 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=34790
M594 207 1123 1729 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=38930
M595 1730 1113 207 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=39790
M596 207 1119 1731 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=43930
M597 1732 1115 207 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=44790
M598 207 1135 1733 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=48930
M599 1734 1099 207 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=32120 $Y=49790
M600 208 1084 766 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=3930
M601 208 1086 736 2400 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=4800
M602 208 1094 767 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=8930
M603 208 1096 737 2401 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=9800
M604 208 1104 768 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=13930
M605 208 1106 738 2402 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=14800
M606 208 1114 769 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=18930
M607 208 1116 739 2403 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=19800
M608 208 1124 770 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=23930
M609 208 1126 740 2404 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=24800
M610 208 1134 771 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=28930
M611 208 1136 741 2405 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=29800
M612 208 1137 772 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=33930
M613 208 1109 742 2406 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=34800
M614 208 1123 773 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=38930
M615 208 1113 743 2407 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=39800
M616 208 1119 774 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=43930
M617 208 1115 744 2408 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=44800
M618 208 1135 775 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=48930
M619 208 1099 745 2409 N_18_G2 l=2.29302e-07 w=2.15e-07 $X=33830 $Y=49800
X620 179 692 700 708 734 745 1141 1174 1185 1218 1229 1262 1273 1306 1317 1350 1361 1394 1405 1438 1449 1482 1493 1526 1537 1570 1581 1614 1625 1658 1669 1702 1713 1746 776 1087 1127 1164 1162 1208 1206 1252 1250 1296 1294 1340 1338 1384 1382 1428 1426 1472 1470 1516 1514 1560 1558 1604 1602 1648 1646 1692 1690 1736 1734 1107 1097 1757 2398 2409 2410 MERGE_2_VIRTUAL_C_VIRTUAL_C $X=30 $Y=50000 $T=0 50000 0 0
X621 179 673 672 671 724 735 1143 1163 1187 1207 1231 1251 1275 1295 1319 1339 1363 1383 1407 1427 1451 1471 1495 1515 1539 1559 1583 1603 1627 1647 1671 1691 1715 1735 766 1082 1078 1176 1142 1220 1186 1264 1230 1308 1274 1352 1318 1396 1362 1440 1406 1484 1450 1528 1494 1572 1538 1616 1582 1660 1626 1704 1670 1748 1714 1080 1081 1758 2388 2399 2400 MERGE_2_VIRTUAL_C_VIRTUAL_C $X=30 $Y=0 $T=0 0 0 0
X622 179 681 680 679 725 736 1145 1165 1189 1209 1233 1253 1277 1297 1321 1341 1365 1385 1409 1429 1453 1473 1497 1517 1541 1561 1585 1605 1629 1649 1673 1693 1717 1737 767 1092 1088 1177 1144 1221 1188 1265 1232 1309 1276 1353 1320 1397 1364 1441 1408 1485 1452 1529 1496 1573 1540 1617 1584 1661 1628 1705 1672 1749 1716 1090 1091 1759 2389 2400 2401 MERGE_2_VIRTUAL_C_VIRTUAL_C $X=30 $Y=5000 $T=0 5000 0 0
X623 179 689 688 687 726 737 1147 1166 1191 1210 1235 1254 1279 1298 1323 1342 1367 1386 1411 1430 1455 1474 1499 1518 1543 1562 1587 1606 1631 1650 1675 1694 1719 1738 768 1102 1098 1178 1146 1222 1190 1266 1234 1310 1278 1354 1322 1398 1366 1442 1410 1486 1454 1530 1498 1574 1542 1618 1586 1662 1630 1706 1674 1750 1718 1100 1101 1760 2390 2401 2402 MERGE_2_VIRTUAL_C_VIRTUAL_C $X=30 $Y=10000 $T=0 10000 0 0
X624 179 697 696 695 727 738 1149 1167 1193 1211 1237 1255 1281 1299 1325 1343 1369 1387 1413 1431 1457 1475 1501 1519 1545 1563 1589 1607 1633 1651 1677 1695 1721 1739 769 1112 1108 1179 1148 1223 1192 1267 1236 1311 1280 1355 1324 1399 1368 1443 1412 1487 1456 1531 1500 1575 1544 1619 1588 1663 1632 1707 1676 1751 1720 1110 1111 1761 2391 2402 2403 MERGE_2_VIRTUAL_C_VIRTUAL_C $X=30 $Y=15000 $T=0 15000 0 0
X625 179 705 704 703 728 739 1151 1168 1195 1212 1239 1256 1283 1300 1327 1344 1371 1388 1415 1432 1459 1476 1503 1520 1547 1564 1591 1608 1635 1652 1679 1696 1723 1740 770 1122 1118 1180 1150 1224 1194 1268 1238 1312 1282 1356 1326 1400 1370 1444 1414 1488 1458 1532 1502 1576 1546 1620 1590 1664 1634 1708 1678 1752 1722 1120 1121 1762 2392 2403 2404 MERGE_2_VIRTUAL_C_VIRTUAL_C $X=30 $Y=20000 $T=0 20000 0 0
X626 179 713 712 711 729 740 1153 1169 1197 1213 1241 1257 1285 1301 1329 1345 1373 1389 1417 1433 1461 1477 1505 1521 1549 1565 1593 1609 1637 1653 1681 1697 1725 1741 771 1132 1128 1181 1152 1225 1196 1269 1240 1313 1284 1357 1328 1401 1372 1445 1416 1489 1460 1533 1504 1577 1548 1621 1592 1665 1636 1709 1680 1753 1724 1130 1131 1763 2393 2404 2405 MERGE_2_VIRTUAL_C_VIRTUAL_C $X=30 $Y=25000 $T=0 25000 0 0
X627 179 721 720 719 730 741 1155 1170 1199 1214 1243 1258 1287 1302 1331 1346 1375 1390 1419 1434 1463 1478 1507 1522 1551 1566 1595 1610 1639 1654 1683 1698 1727 1742 772 1077 1138 1182 1154 1226 1198 1270 1242 1314 1286 1358 1330 1402 1374 1446 1418 1490 1462 1534 1506 1578 1550 1622 1594 1666 1638 1710 1682 1754 1726 1140 1079 1764 2394 2405 2406 MERGE_2_VIRTUAL_C_VIRTUAL_C $X=30 $Y=30000 $T=0 30000 0 0
X628 179 717 693 685 731 742 1157 1171 1201 1215 1245 1259 1289 1303 1333 1347 1377 1391 1421 1435 1465 1479 1509 1523 1553 1567 1597 1611 1641 1655 1685 1699 1729 1743 773 1133 1129 1183 1156 1227 1200 1271 1244 1315 1288 1359 1332 1403 1376 1447 1420 1491 1464 1535 1508 1579 1552 1623 1596 1667 1640 1711 1684 1755 1728 1117 1139 1765 2395 2406 2407 MERGE_2_VIRTUAL_C_VIRTUAL_C $X=30 $Y=35000 $T=0 35000 0 0
X629 179 701 707 709 732 743 1159 1172 1203 1216 1247 1260 1291 1304 1335 1348 1379 1392 1423 1436 1467 1480 1511 1524 1555 1568 1599 1612 1643 1656 1687 1700 1731 1744 774 1083 1103 1184 1158 1228 1202 1272 1246 1316 1290 1360 1334 1404 1378 1448 1422 1492 1466 1536 1510 1580 1554 1624 1598 1668 1642 1712 1686 1756 1730 1093 1089 1766 2396 2407 2408 MERGE_2_VIRTUAL_C_VIRTUAL_C $X=30 $Y=40000 $T=0 40000 0 0
X630 179 669 675 677 733 744 1161 1173 1205 1217 1249 1261 1293 1305 1337 1349 1381 1393 1425 1437 1469 1481 1513 1525 1557 1569 1601 1613 1645 1657 1689 1701 1733 1745 775 1085 1125 1175 1160 1219 1204 1263 1248 1307 1292 1351 1336 1395 1380 1439 1424 1483 1468 1527 1512 1571 1556 1615 1600 1659 1644 1703 1688 1747 1732 1105 1095 1767 2397 2408 2409 MERGE_2_VIRTUAL_C_VIRTUAL_C $X=30 $Y=45000 $T=0 45000 0 0
.ENDS



*******************************************************************************
* Main Circuit Netlist:                                                       *
*                            25                                                 *
* Block: HN_ADFULHX2                                                        *
* Last Time Saved: Dec 19 09:16:36 2006                                       *
*******************************************************************************
.SUBCKT HN_ADFULHX2 A  B  CI  CO  VSS  VDD  S  
MM5 11 B 10 VSS N l=2.4e-07 w=2.32e-06
MM7 11 12 9 VSS N l=2.4e-07 w=2.32e-06
MM9 13 B 9 VSS N l=2.4e-07 w=2.32e-06
MM12 10 12 13 VSS N l=2.4e-07 w=2.31e-06
MM16 16 11 12 VSS N l=2.4e-07 w=1.14e-06
MM17 15 13 16 VSS N l=2.4e-07 w=1.14e-06
MM18 17 11 15 VSS N l=2.4e-07 w=1.14e-06
MM19 14 13 17 VSS N l=2.4e-07 w=1.14e-06
MM30 11 12 10 VDD P l=2.4e-07 w=3.2e-06
MM32 11 B 9 VDD P l=2.4e-07 w=3.21e-06
MM34 13 12 9 VDD P l=2.4e-07 w=3.21e-06
MM36 10 B 13 VDD P l=2.4e-07 w=3.21e-06
MM42 16 13 12 VDD P l=2.4e-07 w=1.68e-06
MM43 15 11 16 VDD P l=2.4e-07 w=1.68e-06
MM44 17 13 15 VDD P l=2.4e-07 w=1.68e-06
MM45 14 11 17 VDD P l=2.4e-07 w=1.68e-06
XG1 A 9 DECAP_INV_G1
XG2 A 8 DECAP_INV_G2
XG3 8 10 DECAP_INV_G1
XG4 B 12 DECAP_INV_G3
XG5 15 14 DECAP_INV_G4
XG6 CI 15 DECAP_INV_G5
XG7 16 CO DECAP_INV_G6
XG8 17 S DECAP_INV_G6
.ENDS

*******************************************************************************
* Main Circuit Netlist:                                                       *
*                            26                                                 *
* Block: HN_MUX2X4                                                          *
* Last Time Saved: Dec 19 09:16:36 2006                                       *
*******************************************************************************

.SUBCKT HN_MUX2X4 B  S0  A  Y  VSS  VDD  
MM2 10 S0 7 VSS N l=2.4e-07 w=1.1e-06
MM3 9 8 10 VSS N l=2.4e-07 w=1e-06
MM9 10 8 7 VDD P l=2.4e-07 w=1.26e-06
MM10 9 S0 10 VDD P l=2.4e-07 w=1.56e-06
XG229 S0 8 DECAP_INV_G166
XG230 B 7 DECAP_INV_G4
XG231 A 9 DECAP_INV_G6
XG232 10 Y DECAP_INV_G3
.ENDS

*******************************************************************************
* Main Circuit Netlist:                                                       *
*                            27                                                 *
* Block: SDC64X32H25_C4_MAINCTRL_C4                                                         *
* Last Time Saved: Dec 19 09:16:36 2006                                       *
*******************************************************************************

.SUBCKT SDC64X32H25_C4_MAINCTRL_C4 VDD  VSS  CLK  ZCLK  WLPULSEB  DLPRECH  SCLK  SCLK2  ZSCLK  ZSCLK2  CEB  ZWLODD  ZWLEVEN  WEB  WEPG  ZFPRECH  SAEN  X0[1]  X0[0]  20  
MM5 29 28 ZCLK VSS N l=2.4e-07 w=1.2e-05
MM14 CLK 28 30 VSS N l=2.4e-07 w=4e-06
MM17 VSS 21 30 VSS N l=4e-07 w=8e-07
MM39 28 ZCLK 43 VSS N l=2.4e-07 w=1.5e-06
MM54 21 CLK 22 VSS N l=2.4e-07 w=3e-06
MM66 WEPG 31 VSS VSS N l=4e-07 w=4e-06
MM69 CLK 35 50 VSS N l=2.4e-07 w=1.5e-06
MM76 25 CLK 32 VSS N l=2.4e-07 w=1.2e-06
MM82 53 ZCLK 52 VSS N l=2.4e-07 w=1.2e-06
MM122 VDD 28 29 VDD P l=2.4e-07 w=8e-07
MM130 29 21 ZCLK VDD P l=2.4e-07 w=4e-06
MM132 30 21 CLK VDD P l=2.4e-07 w=1.5e-05
MM157 28 CLK 43 VDD P l=2.4e-07 w=3e-06
MM172 21 ZCLK 22 VDD P l=2.4e-07 w=4e-06
MM183 50 35 VDD VDD P l=2.4e-07 w=8e-07
MM187 CLK 36 50 VDD P l=2.4e-07 w=3e-06
MM194 25 ZCLK 32 VDD P l=2.4e-07 w=2.5e-06
MM201 53 CLK 52 VDD P l=2.4e-07 w=2.4e-06
DX333D0 VSS CEB NP AREA=2.088e-12
DX649D0 VSS WEB NP AREA=2.088e-12
XG499 X0[1] 49 23 40 DECAP_NAND3_G305
XG500 21 22 24 DECAP_NAND2_G306
XG501 X0[0] 49 23 46 DECAP_NAND3_G305
XG502 DLPRECH 26 61 33 DECAP_NAND3_G305
XG503 20 24 50 35 DECAP_NAND3_G307
XG504 25 60 55 DECAP_NAND2_G299
XG505 27 35 37 59 DECAP_NAND3_G305
XG506 WLPULSEB 35 60 DECAP_NAND2_G308
XG507 35 37 61 DECAP_NAND2_G306
XG508 29 SCLK DECAP_INV_G309
XG509 CLK ZCLK DECAP_INV_G310
XG510 29 SCLK2 DECAP_INV_G311
XG511 30 ZSCLK DECAP_INV_G312
XG512 30 ZSCLK2 DECAP_INV_G313
XG513 44 ZWLODD DECAP_INV_G314
XG514 CEB 38 DECAP_INV_G304
XG515 38 42 DECAP_INV_G304
XG516 42 43 DECAP_INV_G315
XG517 40 44 DECAP_INV_G310
XG518 21 28 DECAP_INV_G298
XG519 46 45 DECAP_INV_G310
XG520 45 ZWLEVEN DECAP_INV_G314
XG521 28 21 DECAP_INV_G316
XG522 49 22 DECAP_INV_G298
XG523 22 49 DECAP_INV_G316
XG524 59 31 DECAP_INV_G315
XG525 51 27 DECAP_INV_G317
XG526 53 32 DECAP_INV_G318
XG527 33 WEPG DECAP_INV_G319
XG528 55 34 DECAP_INV_G315
XG529 31 DLPRECH DECAP_INV_G319
XG530 54 52 DECAP_INV_G302
XG531 37 51 DECAP_INV_G320
XG532 26 25 DECAP_INV_G298
XG533 32 53 DECAP_INV_G298
XG534 57 54 DECAP_INV_G304
XG535 25 26 DECAP_INV_G321
XG536 23 37 DECAP_INV_G322
XG537 WEB 57 DECAP_INV_G304
XG538 34 SAEN DECAP_INV_G319
XG539 WLPULSEB 23 DECAP_INV_G323
XG540 59 ZFPRECH DECAP_INV_G319
XG541 35 36 DECAP_INV_G302
XG542 36 WLPULSEB DECAP_INV_G316
.ENDS

*******************************************************************************
* Main Circuit Netlist:                                                       *
*                            28                                                 *
* Block: SDC64X32H25_C4_MAINCTRL_C4                                                         *
* Last Time Saved: Dec 19 09:16:36 2006                                       *
*******************************************************************************


