
.SUBCKT ram DOUT_7_  DOUT_6_  DOUT_5_  DOUT_4_  DOUT_3_  DOUT_2_  DOUT_1_  DOUT_0_  A_9_  A_8_  A_7_  A_6_  A_5_  A_4_  A_3_  A_2_  A_1_  A_0_  CLK  CS  DIN_7_  DIN_6_  DIN_5_  DIN_4_  DIN_3_  DIN_2_  DIN_1_  DIN_0_  RD  WR  gnd  vdd  
XI11_7/XI2/MN0_15 XI11_7/net21_0_ ysel_15_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll]
XI11_7/XI2/MN0_14 XI11_7/net21_1_ ysel_14_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_13 XI11_7/net21_2_ ysel_13_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_12 XI11_7/net21_3_ ysel_12_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_11 XI11_7/net21_4_ ysel_11_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_10 XI11_7/net21_5_ ysel_10_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_9 XI11_7/net21_6_ ysel_9_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_8 XI11_7/net21_7_ ysel_8_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_7 XI11_7/net21_8_ ysel_7_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_6 XI11_7/net21_9_ ysel_6_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_5 XI11_7/net21_10_ ysel_5_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_4 XI11_7/net21_11_ ysel_4_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_3 XI11_7/net21_12_ ysel_3_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_2 XI11_7/net21_13_ ysel_2_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_1 XI11_7/net21_14_ ysel_1_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_0 XI11_7/net21_15_ ysel_0_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_15 XI11_7/net20_0_ ysel_15_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_14 XI11_7/net20_1_ ysel_14_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_13 XI11_7/net20_2_ ysel_13_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_12 XI11_7/net20_3_ ysel_12_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_11 XI11_7/net20_4_ ysel_11_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_10 XI11_7/net20_5_ ysel_10_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_9 XI11_7/net20_6_ ysel_9_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_8 XI11_7/net20_7_ ysel_8_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_7 XI11_7/net20_8_ ysel_7_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_6 XI11_7/net20_9_ ysel_6_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_5 XI11_7/net20_10_ ysel_5_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_4 XI11_7/net20_11_ ysel_4_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_3 XI11_7/net20_12_ ysel_3_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_2 XI11_7/net20_13_ ysel_2_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_1 XI11_7/net20_14_ ysel_1_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_0 XI11_7/net20_15_ ysel_0_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI4/MN8 vdd XI11_7/XI4/net8 XI11_7/net12 vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_7/XI4/MP0 XI11_7/net9 XI11_7/XI4/net23 vdd vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_7/XI4/MP4 XI11_7/net12 XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI4/MP1 XI11_7/net9 XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI4/MP5 XI11_7/net12 XI11_7/preck XI11_7/net9 vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI4/MN7 vdd XI11_7/XI4/net090 DOUT_7_ vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_7/XI4/MP3 gnd XI11_7/XI4/net089 XI11_7/net12 gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_7/XI4/MN5 XI11_7/net9 XI11_7/XI4/net0103 gnd gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_7/XI4/MN4 XI11_7/XI4/data_out_ XI11_7/XI4/net32 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_7/XI4/MN0 XI11_7/XI4/data_out XI11_7/XI4/net52 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_7/XI4/MN9 gnd XI11_7/XI4/net0112 DOUT_7_ gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_7/XI1_15/MP2 XI11_7/net20_0_ XI11_7/preck XI11_7/net21_0_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_15/MP1 XI11_7/net20_0_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_15/MP0 XI11_7/net21_0_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_14/MP2 XI11_7/net20_1_ XI11_7/preck XI11_7/net21_1_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_14/MP1 XI11_7/net20_1_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_14/MP0 XI11_7/net21_1_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_13/MP2 XI11_7/net20_2_ XI11_7/preck XI11_7/net21_2_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_13/MP1 XI11_7/net20_2_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_13/MP0 XI11_7/net21_2_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_12/MP2 XI11_7/net20_3_ XI11_7/preck XI11_7/net21_3_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_12/MP1 XI11_7/net20_3_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_12/MP0 XI11_7/net21_3_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_11/MP2 XI11_7/net20_4_ XI11_7/preck XI11_7/net21_4_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_11/MP1 XI11_7/net20_4_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_11/MP0 XI11_7/net21_4_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_10/MP2 XI11_7/net20_5_ XI11_7/preck XI11_7/net21_5_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_10/MP1 XI11_7/net20_5_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_10/MP0 XI11_7/net21_5_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_9/MP2 XI11_7/net20_6_ XI11_7/preck XI11_7/net21_6_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_9/MP1 XI11_7/net20_6_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_9/MP0 XI11_7/net21_6_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_8/MP2 XI11_7/net20_7_ XI11_7/preck XI11_7/net21_7_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_8/MP1 XI11_7/net20_7_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_8/MP0 XI11_7/net21_7_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_7/MP2 XI11_7/net20_8_ XI11_7/preck XI11_7/net21_8_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_7/MP1 XI11_7/net20_8_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_7/MP0 XI11_7/net21_8_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_6/MP2 XI11_7/net20_9_ XI11_7/preck XI11_7/net21_9_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_6/MP1 XI11_7/net20_9_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_6/MP0 XI11_7/net21_9_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_5/MP2 XI11_7/net20_10_ XI11_7/preck XI11_7/net21_10_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_5/MP1 XI11_7/net20_10_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_5/MP0 XI11_7/net21_10_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_4/MP2 XI11_7/net20_11_ XI11_7/preck XI11_7/net21_11_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_4/MP1 XI11_7/net20_11_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_4/MP0 XI11_7/net21_11_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_3/MP2 XI11_7/net20_12_ XI11_7/preck XI11_7/net21_12_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_3/MP1 XI11_7/net20_12_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_3/MP0 XI11_7/net21_12_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_2/MP2 XI11_7/net20_13_ XI11_7/preck XI11_7/net21_13_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_2/MP1 XI11_7/net20_13_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_2/MP0 XI11_7/net21_13_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_1/MP2 XI11_7/net20_14_ XI11_7/preck XI11_7/net21_14_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_1/MP1 XI11_7/net20_14_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_1/MP0 XI11_7/net21_14_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_0/MP2 XI11_7/net20_15_ XI11_7/preck XI11_7/net21_15_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_0/MP1 XI11_7/net20_15_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_0/MP0 XI11_7/net21_15_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI0/MN0_15 gnd gnd XI11_7/net21_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_14 gnd gnd XI11_7/net21_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_13 gnd gnd XI11_7/net21_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_12 gnd gnd XI11_7/net21_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_11 gnd gnd XI11_7/net21_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_10 gnd gnd XI11_7/net21_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_9 gnd gnd XI11_7/net21_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_8 gnd gnd XI11_7/net21_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_7 gnd gnd XI11_7/net21_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_6 gnd gnd XI11_7/net21_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_5 gnd gnd XI11_7/net21_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_4 gnd gnd XI11_7/net21_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_3 gnd gnd XI11_7/net21_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_2 gnd gnd XI11_7/net21_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_1 gnd gnd XI11_7/net21_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_0 gnd gnd XI11_7/net21_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_15 gnd gnd XI11_7/net20_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_14 gnd gnd XI11_7/net20_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_13 gnd gnd XI11_7/net20_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_12 gnd gnd XI11_7/net20_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_11 gnd gnd XI11_7/net20_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_10 gnd gnd XI11_7/net20_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_9 gnd gnd XI11_7/net20_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_8 gnd gnd XI11_7/net20_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_7 gnd gnd XI11_7/net20_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_6 gnd gnd XI11_7/net20_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_5 gnd gnd XI11_7/net20_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_4 gnd gnd XI11_7/net20_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_3 gnd gnd XI11_7/net20_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_2 gnd gnd XI11_7/net20_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_1 gnd gnd XI11_7/net20_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_0 gnd gnd XI11_7/net20_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_15 XI11_7/net21_0_ xsel_63_ XI11_7/XI0/XI0_63/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_14 XI11_7/net21_1_ xsel_63_ XI11_7/XI0/XI0_63/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_13 XI11_7/net21_2_ xsel_63_ XI11_7/XI0/XI0_63/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_12 XI11_7/net21_3_ xsel_63_ XI11_7/XI0/XI0_63/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_11 XI11_7/net21_4_ xsel_63_ XI11_7/XI0/XI0_63/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_10 XI11_7/net21_5_ xsel_63_ XI11_7/XI0/XI0_63/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_9 XI11_7/net21_6_ xsel_63_ XI11_7/XI0/XI0_63/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_8 XI11_7/net21_7_ xsel_63_ XI11_7/XI0/XI0_63/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_7 XI11_7/net21_8_ xsel_63_ XI11_7/XI0/XI0_63/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_6 XI11_7/net21_9_ xsel_63_ XI11_7/XI0/XI0_63/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_5 XI11_7/net21_10_ xsel_63_ XI11_7/XI0/XI0_63/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_4 XI11_7/net21_11_ xsel_63_ XI11_7/XI0/XI0_63/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_3 XI11_7/net21_12_ xsel_63_ XI11_7/XI0/XI0_63/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_2 XI11_7/net21_13_ xsel_63_ XI11_7/XI0/XI0_63/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_1 XI11_7/net21_14_ xsel_63_ XI11_7/XI0/XI0_63/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_0 XI11_7/net21_15_ xsel_63_ XI11_7/XI0/XI0_63/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_15 XI11_7/XI0/XI0_63/d__15_ xsel_63_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_14 XI11_7/XI0/XI0_63/d__14_ xsel_63_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_13 XI11_7/XI0/XI0_63/d__13_ xsel_63_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_12 XI11_7/XI0/XI0_63/d__12_ xsel_63_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_11 XI11_7/XI0/XI0_63/d__11_ xsel_63_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_10 XI11_7/XI0/XI0_63/d__10_ xsel_63_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_9 XI11_7/XI0/XI0_63/d__9_ xsel_63_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_8 XI11_7/XI0/XI0_63/d__8_ xsel_63_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_7 XI11_7/XI0/XI0_63/d__7_ xsel_63_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_6 XI11_7/XI0/XI0_63/d__6_ xsel_63_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_5 XI11_7/XI0/XI0_63/d__5_ xsel_63_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_4 XI11_7/XI0/XI0_63/d__4_ xsel_63_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_3 XI11_7/XI0/XI0_63/d__3_ xsel_63_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_2 XI11_7/XI0/XI0_63/d__2_ xsel_63_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_1 XI11_7/XI0/XI0_63/d__1_ xsel_63_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_0 XI11_7/XI0/XI0_63/d__0_ xsel_63_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_15 XI11_7/net21_0_ xsel_62_ XI11_7/XI0/XI0_62/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_14 XI11_7/net21_1_ xsel_62_ XI11_7/XI0/XI0_62/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_13 XI11_7/net21_2_ xsel_62_ XI11_7/XI0/XI0_62/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_12 XI11_7/net21_3_ xsel_62_ XI11_7/XI0/XI0_62/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_11 XI11_7/net21_4_ xsel_62_ XI11_7/XI0/XI0_62/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_10 XI11_7/net21_5_ xsel_62_ XI11_7/XI0/XI0_62/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_9 XI11_7/net21_6_ xsel_62_ XI11_7/XI0/XI0_62/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_8 XI11_7/net21_7_ xsel_62_ XI11_7/XI0/XI0_62/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_7 XI11_7/net21_8_ xsel_62_ XI11_7/XI0/XI0_62/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_6 XI11_7/net21_9_ xsel_62_ XI11_7/XI0/XI0_62/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_5 XI11_7/net21_10_ xsel_62_ XI11_7/XI0/XI0_62/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_4 XI11_7/net21_11_ xsel_62_ XI11_7/XI0/XI0_62/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_3 XI11_7/net21_12_ xsel_62_ XI11_7/XI0/XI0_62/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_2 XI11_7/net21_13_ xsel_62_ XI11_7/XI0/XI0_62/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_1 XI11_7/net21_14_ xsel_62_ XI11_7/XI0/XI0_62/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_0 XI11_7/net21_15_ xsel_62_ XI11_7/XI0/XI0_62/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_15 XI11_7/XI0/XI0_62/d__15_ xsel_62_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_14 XI11_7/XI0/XI0_62/d__14_ xsel_62_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_13 XI11_7/XI0/XI0_62/d__13_ xsel_62_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_12 XI11_7/XI0/XI0_62/d__12_ xsel_62_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_11 XI11_7/XI0/XI0_62/d__11_ xsel_62_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_10 XI11_7/XI0/XI0_62/d__10_ xsel_62_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_9 XI11_7/XI0/XI0_62/d__9_ xsel_62_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_8 XI11_7/XI0/XI0_62/d__8_ xsel_62_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_7 XI11_7/XI0/XI0_62/d__7_ xsel_62_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_6 XI11_7/XI0/XI0_62/d__6_ xsel_62_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_5 XI11_7/XI0/XI0_62/d__5_ xsel_62_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_4 XI11_7/XI0/XI0_62/d__4_ xsel_62_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_3 XI11_7/XI0/XI0_62/d__3_ xsel_62_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_2 XI11_7/XI0/XI0_62/d__2_ xsel_62_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_1 XI11_7/XI0/XI0_62/d__1_ xsel_62_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_0 XI11_7/XI0/XI0_62/d__0_ xsel_62_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_15 XI11_7/net21_0_ xsel_61_ XI11_7/XI0/XI0_61/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_14 XI11_7/net21_1_ xsel_61_ XI11_7/XI0/XI0_61/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_13 XI11_7/net21_2_ xsel_61_ XI11_7/XI0/XI0_61/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_12 XI11_7/net21_3_ xsel_61_ XI11_7/XI0/XI0_61/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_11 XI11_7/net21_4_ xsel_61_ XI11_7/XI0/XI0_61/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_10 XI11_7/net21_5_ xsel_61_ XI11_7/XI0/XI0_61/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_9 XI11_7/net21_6_ xsel_61_ XI11_7/XI0/XI0_61/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_8 XI11_7/net21_7_ xsel_61_ XI11_7/XI0/XI0_61/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_7 XI11_7/net21_8_ xsel_61_ XI11_7/XI0/XI0_61/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_6 XI11_7/net21_9_ xsel_61_ XI11_7/XI0/XI0_61/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_5 XI11_7/net21_10_ xsel_61_ XI11_7/XI0/XI0_61/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_4 XI11_7/net21_11_ xsel_61_ XI11_7/XI0/XI0_61/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_3 XI11_7/net21_12_ xsel_61_ XI11_7/XI0/XI0_61/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_2 XI11_7/net21_13_ xsel_61_ XI11_7/XI0/XI0_61/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_1 XI11_7/net21_14_ xsel_61_ XI11_7/XI0/XI0_61/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_0 XI11_7/net21_15_ xsel_61_ XI11_7/XI0/XI0_61/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_15 XI11_7/XI0/XI0_61/d__15_ xsel_61_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_14 XI11_7/XI0/XI0_61/d__14_ xsel_61_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_13 XI11_7/XI0/XI0_61/d__13_ xsel_61_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_12 XI11_7/XI0/XI0_61/d__12_ xsel_61_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_11 XI11_7/XI0/XI0_61/d__11_ xsel_61_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_10 XI11_7/XI0/XI0_61/d__10_ xsel_61_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_9 XI11_7/XI0/XI0_61/d__9_ xsel_61_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_8 XI11_7/XI0/XI0_61/d__8_ xsel_61_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_7 XI11_7/XI0/XI0_61/d__7_ xsel_61_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_6 XI11_7/XI0/XI0_61/d__6_ xsel_61_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_5 XI11_7/XI0/XI0_61/d__5_ xsel_61_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_4 XI11_7/XI0/XI0_61/d__4_ xsel_61_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_3 XI11_7/XI0/XI0_61/d__3_ xsel_61_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_2 XI11_7/XI0/XI0_61/d__2_ xsel_61_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_1 XI11_7/XI0/XI0_61/d__1_ xsel_61_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_0 XI11_7/XI0/XI0_61/d__0_ xsel_61_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_15 XI11_7/net21_0_ xsel_60_ XI11_7/XI0/XI0_60/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_14 XI11_7/net21_1_ xsel_60_ XI11_7/XI0/XI0_60/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_13 XI11_7/net21_2_ xsel_60_ XI11_7/XI0/XI0_60/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_12 XI11_7/net21_3_ xsel_60_ XI11_7/XI0/XI0_60/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_11 XI11_7/net21_4_ xsel_60_ XI11_7/XI0/XI0_60/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_10 XI11_7/net21_5_ xsel_60_ XI11_7/XI0/XI0_60/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_9 XI11_7/net21_6_ xsel_60_ XI11_7/XI0/XI0_60/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_8 XI11_7/net21_7_ xsel_60_ XI11_7/XI0/XI0_60/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_7 XI11_7/net21_8_ xsel_60_ XI11_7/XI0/XI0_60/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_6 XI11_7/net21_9_ xsel_60_ XI11_7/XI0/XI0_60/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_5 XI11_7/net21_10_ xsel_60_ XI11_7/XI0/XI0_60/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_4 XI11_7/net21_11_ xsel_60_ XI11_7/XI0/XI0_60/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_3 XI11_7/net21_12_ xsel_60_ XI11_7/XI0/XI0_60/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_2 XI11_7/net21_13_ xsel_60_ XI11_7/XI0/XI0_60/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_1 XI11_7/net21_14_ xsel_60_ XI11_7/XI0/XI0_60/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_0 XI11_7/net21_15_ xsel_60_ XI11_7/XI0/XI0_60/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_15 XI11_7/XI0/XI0_60/d__15_ xsel_60_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_14 XI11_7/XI0/XI0_60/d__14_ xsel_60_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_13 XI11_7/XI0/XI0_60/d__13_ xsel_60_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_12 XI11_7/XI0/XI0_60/d__12_ xsel_60_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_11 XI11_7/XI0/XI0_60/d__11_ xsel_60_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_10 XI11_7/XI0/XI0_60/d__10_ xsel_60_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_9 XI11_7/XI0/XI0_60/d__9_ xsel_60_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_8 XI11_7/XI0/XI0_60/d__8_ xsel_60_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_7 XI11_7/XI0/XI0_60/d__7_ xsel_60_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_6 XI11_7/XI0/XI0_60/d__6_ xsel_60_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_5 XI11_7/XI0/XI0_60/d__5_ xsel_60_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_4 XI11_7/XI0/XI0_60/d__4_ xsel_60_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_3 XI11_7/XI0/XI0_60/d__3_ xsel_60_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_2 XI11_7/XI0/XI0_60/d__2_ xsel_60_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_1 XI11_7/XI0/XI0_60/d__1_ xsel_60_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_0 XI11_7/XI0/XI0_60/d__0_ xsel_60_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_15 XI11_7/net21_0_ xsel_59_ XI11_7/XI0/XI0_59/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_14 XI11_7/net21_1_ xsel_59_ XI11_7/XI0/XI0_59/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_13 XI11_7/net21_2_ xsel_59_ XI11_7/XI0/XI0_59/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_12 XI11_7/net21_3_ xsel_59_ XI11_7/XI0/XI0_59/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_11 XI11_7/net21_4_ xsel_59_ XI11_7/XI0/XI0_59/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_10 XI11_7/net21_5_ xsel_59_ XI11_7/XI0/XI0_59/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_9 XI11_7/net21_6_ xsel_59_ XI11_7/XI0/XI0_59/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_8 XI11_7/net21_7_ xsel_59_ XI11_7/XI0/XI0_59/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_7 XI11_7/net21_8_ xsel_59_ XI11_7/XI0/XI0_59/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_6 XI11_7/net21_9_ xsel_59_ XI11_7/XI0/XI0_59/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_5 XI11_7/net21_10_ xsel_59_ XI11_7/XI0/XI0_59/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_4 XI11_7/net21_11_ xsel_59_ XI11_7/XI0/XI0_59/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_3 XI11_7/net21_12_ xsel_59_ XI11_7/XI0/XI0_59/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_2 XI11_7/net21_13_ xsel_59_ XI11_7/XI0/XI0_59/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_1 XI11_7/net21_14_ xsel_59_ XI11_7/XI0/XI0_59/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_0 XI11_7/net21_15_ xsel_59_ XI11_7/XI0/XI0_59/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_15 XI11_7/XI0/XI0_59/d__15_ xsel_59_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_14 XI11_7/XI0/XI0_59/d__14_ xsel_59_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_13 XI11_7/XI0/XI0_59/d__13_ xsel_59_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_12 XI11_7/XI0/XI0_59/d__12_ xsel_59_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_11 XI11_7/XI0/XI0_59/d__11_ xsel_59_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_10 XI11_7/XI0/XI0_59/d__10_ xsel_59_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_9 XI11_7/XI0/XI0_59/d__9_ xsel_59_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_8 XI11_7/XI0/XI0_59/d__8_ xsel_59_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_7 XI11_7/XI0/XI0_59/d__7_ xsel_59_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_6 XI11_7/XI0/XI0_59/d__6_ xsel_59_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_5 XI11_7/XI0/XI0_59/d__5_ xsel_59_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_4 XI11_7/XI0/XI0_59/d__4_ xsel_59_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_3 XI11_7/XI0/XI0_59/d__3_ xsel_59_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_2 XI11_7/XI0/XI0_59/d__2_ xsel_59_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_1 XI11_7/XI0/XI0_59/d__1_ xsel_59_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_0 XI11_7/XI0/XI0_59/d__0_ xsel_59_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_15 XI11_7/net21_0_ xsel_58_ XI11_7/XI0/XI0_58/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_14 XI11_7/net21_1_ xsel_58_ XI11_7/XI0/XI0_58/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_13 XI11_7/net21_2_ xsel_58_ XI11_7/XI0/XI0_58/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_12 XI11_7/net21_3_ xsel_58_ XI11_7/XI0/XI0_58/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_11 XI11_7/net21_4_ xsel_58_ XI11_7/XI0/XI0_58/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_10 XI11_7/net21_5_ xsel_58_ XI11_7/XI0/XI0_58/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_9 XI11_7/net21_6_ xsel_58_ XI11_7/XI0/XI0_58/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_8 XI11_7/net21_7_ xsel_58_ XI11_7/XI0/XI0_58/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_7 XI11_7/net21_8_ xsel_58_ XI11_7/XI0/XI0_58/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_6 XI11_7/net21_9_ xsel_58_ XI11_7/XI0/XI0_58/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_5 XI11_7/net21_10_ xsel_58_ XI11_7/XI0/XI0_58/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_4 XI11_7/net21_11_ xsel_58_ XI11_7/XI0/XI0_58/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_3 XI11_7/net21_12_ xsel_58_ XI11_7/XI0/XI0_58/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_2 XI11_7/net21_13_ xsel_58_ XI11_7/XI0/XI0_58/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_1 XI11_7/net21_14_ xsel_58_ XI11_7/XI0/XI0_58/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_0 XI11_7/net21_15_ xsel_58_ XI11_7/XI0/XI0_58/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_15 XI11_7/XI0/XI0_58/d__15_ xsel_58_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_14 XI11_7/XI0/XI0_58/d__14_ xsel_58_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_13 XI11_7/XI0/XI0_58/d__13_ xsel_58_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_12 XI11_7/XI0/XI0_58/d__12_ xsel_58_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_11 XI11_7/XI0/XI0_58/d__11_ xsel_58_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_10 XI11_7/XI0/XI0_58/d__10_ xsel_58_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_9 XI11_7/XI0/XI0_58/d__9_ xsel_58_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_8 XI11_7/XI0/XI0_58/d__8_ xsel_58_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_7 XI11_7/XI0/XI0_58/d__7_ xsel_58_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_6 XI11_7/XI0/XI0_58/d__6_ xsel_58_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_5 XI11_7/XI0/XI0_58/d__5_ xsel_58_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_4 XI11_7/XI0/XI0_58/d__4_ xsel_58_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_3 XI11_7/XI0/XI0_58/d__3_ xsel_58_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_2 XI11_7/XI0/XI0_58/d__2_ xsel_58_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_1 XI11_7/XI0/XI0_58/d__1_ xsel_58_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_0 XI11_7/XI0/XI0_58/d__0_ xsel_58_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_15 XI11_7/net21_0_ xsel_57_ XI11_7/XI0/XI0_57/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_14 XI11_7/net21_1_ xsel_57_ XI11_7/XI0/XI0_57/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_13 XI11_7/net21_2_ xsel_57_ XI11_7/XI0/XI0_57/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_12 XI11_7/net21_3_ xsel_57_ XI11_7/XI0/XI0_57/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_11 XI11_7/net21_4_ xsel_57_ XI11_7/XI0/XI0_57/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_10 XI11_7/net21_5_ xsel_57_ XI11_7/XI0/XI0_57/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_9 XI11_7/net21_6_ xsel_57_ XI11_7/XI0/XI0_57/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_8 XI11_7/net21_7_ xsel_57_ XI11_7/XI0/XI0_57/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_7 XI11_7/net21_8_ xsel_57_ XI11_7/XI0/XI0_57/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_6 XI11_7/net21_9_ xsel_57_ XI11_7/XI0/XI0_57/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_5 XI11_7/net21_10_ xsel_57_ XI11_7/XI0/XI0_57/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_4 XI11_7/net21_11_ xsel_57_ XI11_7/XI0/XI0_57/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_3 XI11_7/net21_12_ xsel_57_ XI11_7/XI0/XI0_57/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_2 XI11_7/net21_13_ xsel_57_ XI11_7/XI0/XI0_57/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_1 XI11_7/net21_14_ xsel_57_ XI11_7/XI0/XI0_57/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_0 XI11_7/net21_15_ xsel_57_ XI11_7/XI0/XI0_57/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_15 XI11_7/XI0/XI0_57/d__15_ xsel_57_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_14 XI11_7/XI0/XI0_57/d__14_ xsel_57_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_13 XI11_7/XI0/XI0_57/d__13_ xsel_57_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_12 XI11_7/XI0/XI0_57/d__12_ xsel_57_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_11 XI11_7/XI0/XI0_57/d__11_ xsel_57_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_10 XI11_7/XI0/XI0_57/d__10_ xsel_57_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_9 XI11_7/XI0/XI0_57/d__9_ xsel_57_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_8 XI11_7/XI0/XI0_57/d__8_ xsel_57_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_7 XI11_7/XI0/XI0_57/d__7_ xsel_57_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_6 XI11_7/XI0/XI0_57/d__6_ xsel_57_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_5 XI11_7/XI0/XI0_57/d__5_ xsel_57_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_4 XI11_7/XI0/XI0_57/d__4_ xsel_57_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_3 XI11_7/XI0/XI0_57/d__3_ xsel_57_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_2 XI11_7/XI0/XI0_57/d__2_ xsel_57_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_1 XI11_7/XI0/XI0_57/d__1_ xsel_57_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_0 XI11_7/XI0/XI0_57/d__0_ xsel_57_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_15 XI11_7/net21_0_ xsel_56_ XI11_7/XI0/XI0_56/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_14 XI11_7/net21_1_ xsel_56_ XI11_7/XI0/XI0_56/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_13 XI11_7/net21_2_ xsel_56_ XI11_7/XI0/XI0_56/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_12 XI11_7/net21_3_ xsel_56_ XI11_7/XI0/XI0_56/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_11 XI11_7/net21_4_ xsel_56_ XI11_7/XI0/XI0_56/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_10 XI11_7/net21_5_ xsel_56_ XI11_7/XI0/XI0_56/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_9 XI11_7/net21_6_ xsel_56_ XI11_7/XI0/XI0_56/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_8 XI11_7/net21_7_ xsel_56_ XI11_7/XI0/XI0_56/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_7 XI11_7/net21_8_ xsel_56_ XI11_7/XI0/XI0_56/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_6 XI11_7/net21_9_ xsel_56_ XI11_7/XI0/XI0_56/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_5 XI11_7/net21_10_ xsel_56_ XI11_7/XI0/XI0_56/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_4 XI11_7/net21_11_ xsel_56_ XI11_7/XI0/XI0_56/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_3 XI11_7/net21_12_ xsel_56_ XI11_7/XI0/XI0_56/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_2 XI11_7/net21_13_ xsel_56_ XI11_7/XI0/XI0_56/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_1 XI11_7/net21_14_ xsel_56_ XI11_7/XI0/XI0_56/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_0 XI11_7/net21_15_ xsel_56_ XI11_7/XI0/XI0_56/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_15 XI11_7/XI0/XI0_56/d__15_ xsel_56_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_14 XI11_7/XI0/XI0_56/d__14_ xsel_56_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_13 XI11_7/XI0/XI0_56/d__13_ xsel_56_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_12 XI11_7/XI0/XI0_56/d__12_ xsel_56_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_11 XI11_7/XI0/XI0_56/d__11_ xsel_56_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_10 XI11_7/XI0/XI0_56/d__10_ xsel_56_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_9 XI11_7/XI0/XI0_56/d__9_ xsel_56_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_8 XI11_7/XI0/XI0_56/d__8_ xsel_56_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_7 XI11_7/XI0/XI0_56/d__7_ xsel_56_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_6 XI11_7/XI0/XI0_56/d__6_ xsel_56_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_5 XI11_7/XI0/XI0_56/d__5_ xsel_56_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_4 XI11_7/XI0/XI0_56/d__4_ xsel_56_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_3 XI11_7/XI0/XI0_56/d__3_ xsel_56_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_2 XI11_7/XI0/XI0_56/d__2_ xsel_56_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_1 XI11_7/XI0/XI0_56/d__1_ xsel_56_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_0 XI11_7/XI0/XI0_56/d__0_ xsel_56_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_15 XI11_7/net21_0_ xsel_55_ XI11_7/XI0/XI0_55/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_14 XI11_7/net21_1_ xsel_55_ XI11_7/XI0/XI0_55/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_13 XI11_7/net21_2_ xsel_55_ XI11_7/XI0/XI0_55/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_12 XI11_7/net21_3_ xsel_55_ XI11_7/XI0/XI0_55/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_11 XI11_7/net21_4_ xsel_55_ XI11_7/XI0/XI0_55/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_10 XI11_7/net21_5_ xsel_55_ XI11_7/XI0/XI0_55/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_9 XI11_7/net21_6_ xsel_55_ XI11_7/XI0/XI0_55/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_8 XI11_7/net21_7_ xsel_55_ XI11_7/XI0/XI0_55/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_7 XI11_7/net21_8_ xsel_55_ XI11_7/XI0/XI0_55/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_6 XI11_7/net21_9_ xsel_55_ XI11_7/XI0/XI0_55/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_5 XI11_7/net21_10_ xsel_55_ XI11_7/XI0/XI0_55/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_4 XI11_7/net21_11_ xsel_55_ XI11_7/XI0/XI0_55/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_3 XI11_7/net21_12_ xsel_55_ XI11_7/XI0/XI0_55/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_2 XI11_7/net21_13_ xsel_55_ XI11_7/XI0/XI0_55/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_1 XI11_7/net21_14_ xsel_55_ XI11_7/XI0/XI0_55/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_0 XI11_7/net21_15_ xsel_55_ XI11_7/XI0/XI0_55/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_15 XI11_7/XI0/XI0_55/d__15_ xsel_55_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_14 XI11_7/XI0/XI0_55/d__14_ xsel_55_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_13 XI11_7/XI0/XI0_55/d__13_ xsel_55_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_12 XI11_7/XI0/XI0_55/d__12_ xsel_55_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_11 XI11_7/XI0/XI0_55/d__11_ xsel_55_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_10 XI11_7/XI0/XI0_55/d__10_ xsel_55_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_9 XI11_7/XI0/XI0_55/d__9_ xsel_55_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_8 XI11_7/XI0/XI0_55/d__8_ xsel_55_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_7 XI11_7/XI0/XI0_55/d__7_ xsel_55_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_6 XI11_7/XI0/XI0_55/d__6_ xsel_55_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_5 XI11_7/XI0/XI0_55/d__5_ xsel_55_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_4 XI11_7/XI0/XI0_55/d__4_ xsel_55_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_3 XI11_7/XI0/XI0_55/d__3_ xsel_55_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_2 XI11_7/XI0/XI0_55/d__2_ xsel_55_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_1 XI11_7/XI0/XI0_55/d__1_ xsel_55_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_0 XI11_7/XI0/XI0_55/d__0_ xsel_55_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_15 XI11_7/net21_0_ xsel_54_ XI11_7/XI0/XI0_54/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_14 XI11_7/net21_1_ xsel_54_ XI11_7/XI0/XI0_54/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_13 XI11_7/net21_2_ xsel_54_ XI11_7/XI0/XI0_54/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_12 XI11_7/net21_3_ xsel_54_ XI11_7/XI0/XI0_54/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_11 XI11_7/net21_4_ xsel_54_ XI11_7/XI0/XI0_54/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_10 XI11_7/net21_5_ xsel_54_ XI11_7/XI0/XI0_54/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_9 XI11_7/net21_6_ xsel_54_ XI11_7/XI0/XI0_54/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_8 XI11_7/net21_7_ xsel_54_ XI11_7/XI0/XI0_54/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_7 XI11_7/net21_8_ xsel_54_ XI11_7/XI0/XI0_54/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_6 XI11_7/net21_9_ xsel_54_ XI11_7/XI0/XI0_54/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_5 XI11_7/net21_10_ xsel_54_ XI11_7/XI0/XI0_54/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_4 XI11_7/net21_11_ xsel_54_ XI11_7/XI0/XI0_54/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_3 XI11_7/net21_12_ xsel_54_ XI11_7/XI0/XI0_54/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_2 XI11_7/net21_13_ xsel_54_ XI11_7/XI0/XI0_54/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_1 XI11_7/net21_14_ xsel_54_ XI11_7/XI0/XI0_54/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_0 XI11_7/net21_15_ xsel_54_ XI11_7/XI0/XI0_54/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_15 XI11_7/XI0/XI0_54/d__15_ xsel_54_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_14 XI11_7/XI0/XI0_54/d__14_ xsel_54_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_13 XI11_7/XI0/XI0_54/d__13_ xsel_54_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_12 XI11_7/XI0/XI0_54/d__12_ xsel_54_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_11 XI11_7/XI0/XI0_54/d__11_ xsel_54_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_10 XI11_7/XI0/XI0_54/d__10_ xsel_54_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_9 XI11_7/XI0/XI0_54/d__9_ xsel_54_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_8 XI11_7/XI0/XI0_54/d__8_ xsel_54_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_7 XI11_7/XI0/XI0_54/d__7_ xsel_54_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_6 XI11_7/XI0/XI0_54/d__6_ xsel_54_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_5 XI11_7/XI0/XI0_54/d__5_ xsel_54_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_4 XI11_7/XI0/XI0_54/d__4_ xsel_54_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_3 XI11_7/XI0/XI0_54/d__3_ xsel_54_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_2 XI11_7/XI0/XI0_54/d__2_ xsel_54_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_1 XI11_7/XI0/XI0_54/d__1_ xsel_54_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_0 XI11_7/XI0/XI0_54/d__0_ xsel_54_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_15 XI11_7/net21_0_ xsel_53_ XI11_7/XI0/XI0_53/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_14 XI11_7/net21_1_ xsel_53_ XI11_7/XI0/XI0_53/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_13 XI11_7/net21_2_ xsel_53_ XI11_7/XI0/XI0_53/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_12 XI11_7/net21_3_ xsel_53_ XI11_7/XI0/XI0_53/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_11 XI11_7/net21_4_ xsel_53_ XI11_7/XI0/XI0_53/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_10 XI11_7/net21_5_ xsel_53_ XI11_7/XI0/XI0_53/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_9 XI11_7/net21_6_ xsel_53_ XI11_7/XI0/XI0_53/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_8 XI11_7/net21_7_ xsel_53_ XI11_7/XI0/XI0_53/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_7 XI11_7/net21_8_ xsel_53_ XI11_7/XI0/XI0_53/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_6 XI11_7/net21_9_ xsel_53_ XI11_7/XI0/XI0_53/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_5 XI11_7/net21_10_ xsel_53_ XI11_7/XI0/XI0_53/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_4 XI11_7/net21_11_ xsel_53_ XI11_7/XI0/XI0_53/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_3 XI11_7/net21_12_ xsel_53_ XI11_7/XI0/XI0_53/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_2 XI11_7/net21_13_ xsel_53_ XI11_7/XI0/XI0_53/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_1 XI11_7/net21_14_ xsel_53_ XI11_7/XI0/XI0_53/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_0 XI11_7/net21_15_ xsel_53_ XI11_7/XI0/XI0_53/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_15 XI11_7/XI0/XI0_53/d__15_ xsel_53_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_14 XI11_7/XI0/XI0_53/d__14_ xsel_53_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_13 XI11_7/XI0/XI0_53/d__13_ xsel_53_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_12 XI11_7/XI0/XI0_53/d__12_ xsel_53_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_11 XI11_7/XI0/XI0_53/d__11_ xsel_53_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_10 XI11_7/XI0/XI0_53/d__10_ xsel_53_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_9 XI11_7/XI0/XI0_53/d__9_ xsel_53_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_8 XI11_7/XI0/XI0_53/d__8_ xsel_53_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_7 XI11_7/XI0/XI0_53/d__7_ xsel_53_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_6 XI11_7/XI0/XI0_53/d__6_ xsel_53_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_5 XI11_7/XI0/XI0_53/d__5_ xsel_53_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_4 XI11_7/XI0/XI0_53/d__4_ xsel_53_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_3 XI11_7/XI0/XI0_53/d__3_ xsel_53_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_2 XI11_7/XI0/XI0_53/d__2_ xsel_53_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_1 XI11_7/XI0/XI0_53/d__1_ xsel_53_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_0 XI11_7/XI0/XI0_53/d__0_ xsel_53_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_15 XI11_7/net21_0_ xsel_52_ XI11_7/XI0/XI0_52/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_14 XI11_7/net21_1_ xsel_52_ XI11_7/XI0/XI0_52/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_13 XI11_7/net21_2_ xsel_52_ XI11_7/XI0/XI0_52/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_12 XI11_7/net21_3_ xsel_52_ XI11_7/XI0/XI0_52/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_11 XI11_7/net21_4_ xsel_52_ XI11_7/XI0/XI0_52/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_10 XI11_7/net21_5_ xsel_52_ XI11_7/XI0/XI0_52/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_9 XI11_7/net21_6_ xsel_52_ XI11_7/XI0/XI0_52/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_8 XI11_7/net21_7_ xsel_52_ XI11_7/XI0/XI0_52/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_7 XI11_7/net21_8_ xsel_52_ XI11_7/XI0/XI0_52/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_6 XI11_7/net21_9_ xsel_52_ XI11_7/XI0/XI0_52/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_5 XI11_7/net21_10_ xsel_52_ XI11_7/XI0/XI0_52/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_4 XI11_7/net21_11_ xsel_52_ XI11_7/XI0/XI0_52/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_3 XI11_7/net21_12_ xsel_52_ XI11_7/XI0/XI0_52/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_2 XI11_7/net21_13_ xsel_52_ XI11_7/XI0/XI0_52/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_1 XI11_7/net21_14_ xsel_52_ XI11_7/XI0/XI0_52/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_0 XI11_7/net21_15_ xsel_52_ XI11_7/XI0/XI0_52/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_15 XI11_7/XI0/XI0_52/d__15_ xsel_52_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_14 XI11_7/XI0/XI0_52/d__14_ xsel_52_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_13 XI11_7/XI0/XI0_52/d__13_ xsel_52_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_12 XI11_7/XI0/XI0_52/d__12_ xsel_52_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_11 XI11_7/XI0/XI0_52/d__11_ xsel_52_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_10 XI11_7/XI0/XI0_52/d__10_ xsel_52_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_9 XI11_7/XI0/XI0_52/d__9_ xsel_52_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_8 XI11_7/XI0/XI0_52/d__8_ xsel_52_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_7 XI11_7/XI0/XI0_52/d__7_ xsel_52_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_6 XI11_7/XI0/XI0_52/d__6_ xsel_52_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_5 XI11_7/XI0/XI0_52/d__5_ xsel_52_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_4 XI11_7/XI0/XI0_52/d__4_ xsel_52_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_3 XI11_7/XI0/XI0_52/d__3_ xsel_52_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_2 XI11_7/XI0/XI0_52/d__2_ xsel_52_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_1 XI11_7/XI0/XI0_52/d__1_ xsel_52_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_0 XI11_7/XI0/XI0_52/d__0_ xsel_52_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_15 XI11_7/net21_0_ xsel_51_ XI11_7/XI0/XI0_51/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_14 XI11_7/net21_1_ xsel_51_ XI11_7/XI0/XI0_51/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_13 XI11_7/net21_2_ xsel_51_ XI11_7/XI0/XI0_51/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_12 XI11_7/net21_3_ xsel_51_ XI11_7/XI0/XI0_51/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_11 XI11_7/net21_4_ xsel_51_ XI11_7/XI0/XI0_51/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_10 XI11_7/net21_5_ xsel_51_ XI11_7/XI0/XI0_51/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_9 XI11_7/net21_6_ xsel_51_ XI11_7/XI0/XI0_51/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_8 XI11_7/net21_7_ xsel_51_ XI11_7/XI0/XI0_51/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_7 XI11_7/net21_8_ xsel_51_ XI11_7/XI0/XI0_51/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_6 XI11_7/net21_9_ xsel_51_ XI11_7/XI0/XI0_51/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_5 XI11_7/net21_10_ xsel_51_ XI11_7/XI0/XI0_51/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_4 XI11_7/net21_11_ xsel_51_ XI11_7/XI0/XI0_51/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_3 XI11_7/net21_12_ xsel_51_ XI11_7/XI0/XI0_51/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_2 XI11_7/net21_13_ xsel_51_ XI11_7/XI0/XI0_51/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_1 XI11_7/net21_14_ xsel_51_ XI11_7/XI0/XI0_51/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_0 XI11_7/net21_15_ xsel_51_ XI11_7/XI0/XI0_51/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_15 XI11_7/XI0/XI0_51/d__15_ xsel_51_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_14 XI11_7/XI0/XI0_51/d__14_ xsel_51_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_13 XI11_7/XI0/XI0_51/d__13_ xsel_51_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_12 XI11_7/XI0/XI0_51/d__12_ xsel_51_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_11 XI11_7/XI0/XI0_51/d__11_ xsel_51_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_10 XI11_7/XI0/XI0_51/d__10_ xsel_51_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_9 XI11_7/XI0/XI0_51/d__9_ xsel_51_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_8 XI11_7/XI0/XI0_51/d__8_ xsel_51_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_7 XI11_7/XI0/XI0_51/d__7_ xsel_51_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_6 XI11_7/XI0/XI0_51/d__6_ xsel_51_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_5 XI11_7/XI0/XI0_51/d__5_ xsel_51_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_4 XI11_7/XI0/XI0_51/d__4_ xsel_51_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_3 XI11_7/XI0/XI0_51/d__3_ xsel_51_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_2 XI11_7/XI0/XI0_51/d__2_ xsel_51_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_1 XI11_7/XI0/XI0_51/d__1_ xsel_51_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_0 XI11_7/XI0/XI0_51/d__0_ xsel_51_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_15 XI11_7/net21_0_ xsel_50_ XI11_7/XI0/XI0_50/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_14 XI11_7/net21_1_ xsel_50_ XI11_7/XI0/XI0_50/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_13 XI11_7/net21_2_ xsel_50_ XI11_7/XI0/XI0_50/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_12 XI11_7/net21_3_ xsel_50_ XI11_7/XI0/XI0_50/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_11 XI11_7/net21_4_ xsel_50_ XI11_7/XI0/XI0_50/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_10 XI11_7/net21_5_ xsel_50_ XI11_7/XI0/XI0_50/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_9 XI11_7/net21_6_ xsel_50_ XI11_7/XI0/XI0_50/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_8 XI11_7/net21_7_ xsel_50_ XI11_7/XI0/XI0_50/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_7 XI11_7/net21_8_ xsel_50_ XI11_7/XI0/XI0_50/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_6 XI11_7/net21_9_ xsel_50_ XI11_7/XI0/XI0_50/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_5 XI11_7/net21_10_ xsel_50_ XI11_7/XI0/XI0_50/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_4 XI11_7/net21_11_ xsel_50_ XI11_7/XI0/XI0_50/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_3 XI11_7/net21_12_ xsel_50_ XI11_7/XI0/XI0_50/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_2 XI11_7/net21_13_ xsel_50_ XI11_7/XI0/XI0_50/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_1 XI11_7/net21_14_ xsel_50_ XI11_7/XI0/XI0_50/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_0 XI11_7/net21_15_ xsel_50_ XI11_7/XI0/XI0_50/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_15 XI11_7/XI0/XI0_50/d__15_ xsel_50_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_14 XI11_7/XI0/XI0_50/d__14_ xsel_50_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_13 XI11_7/XI0/XI0_50/d__13_ xsel_50_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_12 XI11_7/XI0/XI0_50/d__12_ xsel_50_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_11 XI11_7/XI0/XI0_50/d__11_ xsel_50_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_10 XI11_7/XI0/XI0_50/d__10_ xsel_50_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_9 XI11_7/XI0/XI0_50/d__9_ xsel_50_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_8 XI11_7/XI0/XI0_50/d__8_ xsel_50_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_7 XI11_7/XI0/XI0_50/d__7_ xsel_50_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_6 XI11_7/XI0/XI0_50/d__6_ xsel_50_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_5 XI11_7/XI0/XI0_50/d__5_ xsel_50_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_4 XI11_7/XI0/XI0_50/d__4_ xsel_50_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_3 XI11_7/XI0/XI0_50/d__3_ xsel_50_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_2 XI11_7/XI0/XI0_50/d__2_ xsel_50_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_1 XI11_7/XI0/XI0_50/d__1_ xsel_50_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_0 XI11_7/XI0/XI0_50/d__0_ xsel_50_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_15 XI11_7/net21_0_ xsel_49_ XI11_7/XI0/XI0_49/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_14 XI11_7/net21_1_ xsel_49_ XI11_7/XI0/XI0_49/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_13 XI11_7/net21_2_ xsel_49_ XI11_7/XI0/XI0_49/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_12 XI11_7/net21_3_ xsel_49_ XI11_7/XI0/XI0_49/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_11 XI11_7/net21_4_ xsel_49_ XI11_7/XI0/XI0_49/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_10 XI11_7/net21_5_ xsel_49_ XI11_7/XI0/XI0_49/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_9 XI11_7/net21_6_ xsel_49_ XI11_7/XI0/XI0_49/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_8 XI11_7/net21_7_ xsel_49_ XI11_7/XI0/XI0_49/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_7 XI11_7/net21_8_ xsel_49_ XI11_7/XI0/XI0_49/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_6 XI11_7/net21_9_ xsel_49_ XI11_7/XI0/XI0_49/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_5 XI11_7/net21_10_ xsel_49_ XI11_7/XI0/XI0_49/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_4 XI11_7/net21_11_ xsel_49_ XI11_7/XI0/XI0_49/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_3 XI11_7/net21_12_ xsel_49_ XI11_7/XI0/XI0_49/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_2 XI11_7/net21_13_ xsel_49_ XI11_7/XI0/XI0_49/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_1 XI11_7/net21_14_ xsel_49_ XI11_7/XI0/XI0_49/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_0 XI11_7/net21_15_ xsel_49_ XI11_7/XI0/XI0_49/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_15 XI11_7/XI0/XI0_49/d__15_ xsel_49_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_14 XI11_7/XI0/XI0_49/d__14_ xsel_49_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_13 XI11_7/XI0/XI0_49/d__13_ xsel_49_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_12 XI11_7/XI0/XI0_49/d__12_ xsel_49_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_11 XI11_7/XI0/XI0_49/d__11_ xsel_49_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_10 XI11_7/XI0/XI0_49/d__10_ xsel_49_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_9 XI11_7/XI0/XI0_49/d__9_ xsel_49_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_8 XI11_7/XI0/XI0_49/d__8_ xsel_49_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_7 XI11_7/XI0/XI0_49/d__7_ xsel_49_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_6 XI11_7/XI0/XI0_49/d__6_ xsel_49_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_5 XI11_7/XI0/XI0_49/d__5_ xsel_49_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_4 XI11_7/XI0/XI0_49/d__4_ xsel_49_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_3 XI11_7/XI0/XI0_49/d__3_ xsel_49_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_2 XI11_7/XI0/XI0_49/d__2_ xsel_49_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_1 XI11_7/XI0/XI0_49/d__1_ xsel_49_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_0 XI11_7/XI0/XI0_49/d__0_ xsel_49_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_15 XI11_7/net21_0_ xsel_48_ XI11_7/XI0/XI0_48/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_14 XI11_7/net21_1_ xsel_48_ XI11_7/XI0/XI0_48/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_13 XI11_7/net21_2_ xsel_48_ XI11_7/XI0/XI0_48/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_12 XI11_7/net21_3_ xsel_48_ XI11_7/XI0/XI0_48/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_11 XI11_7/net21_4_ xsel_48_ XI11_7/XI0/XI0_48/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_10 XI11_7/net21_5_ xsel_48_ XI11_7/XI0/XI0_48/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_9 XI11_7/net21_6_ xsel_48_ XI11_7/XI0/XI0_48/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_8 XI11_7/net21_7_ xsel_48_ XI11_7/XI0/XI0_48/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_7 XI11_7/net21_8_ xsel_48_ XI11_7/XI0/XI0_48/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_6 XI11_7/net21_9_ xsel_48_ XI11_7/XI0/XI0_48/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_5 XI11_7/net21_10_ xsel_48_ XI11_7/XI0/XI0_48/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_4 XI11_7/net21_11_ xsel_48_ XI11_7/XI0/XI0_48/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_3 XI11_7/net21_12_ xsel_48_ XI11_7/XI0/XI0_48/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_2 XI11_7/net21_13_ xsel_48_ XI11_7/XI0/XI0_48/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_1 XI11_7/net21_14_ xsel_48_ XI11_7/XI0/XI0_48/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_0 XI11_7/net21_15_ xsel_48_ XI11_7/XI0/XI0_48/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_15 XI11_7/XI0/XI0_48/d__15_ xsel_48_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_14 XI11_7/XI0/XI0_48/d__14_ xsel_48_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_13 XI11_7/XI0/XI0_48/d__13_ xsel_48_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_12 XI11_7/XI0/XI0_48/d__12_ xsel_48_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_11 XI11_7/XI0/XI0_48/d__11_ xsel_48_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_10 XI11_7/XI0/XI0_48/d__10_ xsel_48_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_9 XI11_7/XI0/XI0_48/d__9_ xsel_48_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_8 XI11_7/XI0/XI0_48/d__8_ xsel_48_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_7 XI11_7/XI0/XI0_48/d__7_ xsel_48_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_6 XI11_7/XI0/XI0_48/d__6_ xsel_48_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_5 XI11_7/XI0/XI0_48/d__5_ xsel_48_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_4 XI11_7/XI0/XI0_48/d__4_ xsel_48_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_3 XI11_7/XI0/XI0_48/d__3_ xsel_48_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_2 XI11_7/XI0/XI0_48/d__2_ xsel_48_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_1 XI11_7/XI0/XI0_48/d__1_ xsel_48_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_0 XI11_7/XI0/XI0_48/d__0_ xsel_48_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_15 XI11_7/net21_0_ xsel_47_ XI11_7/XI0/XI0_47/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_14 XI11_7/net21_1_ xsel_47_ XI11_7/XI0/XI0_47/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_13 XI11_7/net21_2_ xsel_47_ XI11_7/XI0/XI0_47/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_12 XI11_7/net21_3_ xsel_47_ XI11_7/XI0/XI0_47/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_11 XI11_7/net21_4_ xsel_47_ XI11_7/XI0/XI0_47/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_10 XI11_7/net21_5_ xsel_47_ XI11_7/XI0/XI0_47/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_9 XI11_7/net21_6_ xsel_47_ XI11_7/XI0/XI0_47/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_8 XI11_7/net21_7_ xsel_47_ XI11_7/XI0/XI0_47/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_7 XI11_7/net21_8_ xsel_47_ XI11_7/XI0/XI0_47/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_6 XI11_7/net21_9_ xsel_47_ XI11_7/XI0/XI0_47/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_5 XI11_7/net21_10_ xsel_47_ XI11_7/XI0/XI0_47/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_4 XI11_7/net21_11_ xsel_47_ XI11_7/XI0/XI0_47/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_3 XI11_7/net21_12_ xsel_47_ XI11_7/XI0/XI0_47/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_2 XI11_7/net21_13_ xsel_47_ XI11_7/XI0/XI0_47/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_1 XI11_7/net21_14_ xsel_47_ XI11_7/XI0/XI0_47/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_0 XI11_7/net21_15_ xsel_47_ XI11_7/XI0/XI0_47/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_15 XI11_7/XI0/XI0_47/d__15_ xsel_47_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_14 XI11_7/XI0/XI0_47/d__14_ xsel_47_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_13 XI11_7/XI0/XI0_47/d__13_ xsel_47_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_12 XI11_7/XI0/XI0_47/d__12_ xsel_47_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_11 XI11_7/XI0/XI0_47/d__11_ xsel_47_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_10 XI11_7/XI0/XI0_47/d__10_ xsel_47_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_9 XI11_7/XI0/XI0_47/d__9_ xsel_47_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_8 XI11_7/XI0/XI0_47/d__8_ xsel_47_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_7 XI11_7/XI0/XI0_47/d__7_ xsel_47_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_6 XI11_7/XI0/XI0_47/d__6_ xsel_47_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_5 XI11_7/XI0/XI0_47/d__5_ xsel_47_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_4 XI11_7/XI0/XI0_47/d__4_ xsel_47_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_3 XI11_7/XI0/XI0_47/d__3_ xsel_47_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_2 XI11_7/XI0/XI0_47/d__2_ xsel_47_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_1 XI11_7/XI0/XI0_47/d__1_ xsel_47_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_0 XI11_7/XI0/XI0_47/d__0_ xsel_47_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_15 XI11_7/net21_0_ xsel_46_ XI11_7/XI0/XI0_46/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_14 XI11_7/net21_1_ xsel_46_ XI11_7/XI0/XI0_46/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_13 XI11_7/net21_2_ xsel_46_ XI11_7/XI0/XI0_46/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_12 XI11_7/net21_3_ xsel_46_ XI11_7/XI0/XI0_46/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_11 XI11_7/net21_4_ xsel_46_ XI11_7/XI0/XI0_46/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_10 XI11_7/net21_5_ xsel_46_ XI11_7/XI0/XI0_46/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_9 XI11_7/net21_6_ xsel_46_ XI11_7/XI0/XI0_46/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_8 XI11_7/net21_7_ xsel_46_ XI11_7/XI0/XI0_46/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_7 XI11_7/net21_8_ xsel_46_ XI11_7/XI0/XI0_46/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_6 XI11_7/net21_9_ xsel_46_ XI11_7/XI0/XI0_46/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_5 XI11_7/net21_10_ xsel_46_ XI11_7/XI0/XI0_46/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_4 XI11_7/net21_11_ xsel_46_ XI11_7/XI0/XI0_46/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_3 XI11_7/net21_12_ xsel_46_ XI11_7/XI0/XI0_46/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_2 XI11_7/net21_13_ xsel_46_ XI11_7/XI0/XI0_46/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_1 XI11_7/net21_14_ xsel_46_ XI11_7/XI0/XI0_46/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_0 XI11_7/net21_15_ xsel_46_ XI11_7/XI0/XI0_46/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_15 XI11_7/XI0/XI0_46/d__15_ xsel_46_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_14 XI11_7/XI0/XI0_46/d__14_ xsel_46_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_13 XI11_7/XI0/XI0_46/d__13_ xsel_46_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_12 XI11_7/XI0/XI0_46/d__12_ xsel_46_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_11 XI11_7/XI0/XI0_46/d__11_ xsel_46_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_10 XI11_7/XI0/XI0_46/d__10_ xsel_46_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_9 XI11_7/XI0/XI0_46/d__9_ xsel_46_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_8 XI11_7/XI0/XI0_46/d__8_ xsel_46_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_7 XI11_7/XI0/XI0_46/d__7_ xsel_46_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_6 XI11_7/XI0/XI0_46/d__6_ xsel_46_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_5 XI11_7/XI0/XI0_46/d__5_ xsel_46_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_4 XI11_7/XI0/XI0_46/d__4_ xsel_46_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_3 XI11_7/XI0/XI0_46/d__3_ xsel_46_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_2 XI11_7/XI0/XI0_46/d__2_ xsel_46_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_1 XI11_7/XI0/XI0_46/d__1_ xsel_46_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_0 XI11_7/XI0/XI0_46/d__0_ xsel_46_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_15 XI11_7/net21_0_ xsel_45_ XI11_7/XI0/XI0_45/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_14 XI11_7/net21_1_ xsel_45_ XI11_7/XI0/XI0_45/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_13 XI11_7/net21_2_ xsel_45_ XI11_7/XI0/XI0_45/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_12 XI11_7/net21_3_ xsel_45_ XI11_7/XI0/XI0_45/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_11 XI11_7/net21_4_ xsel_45_ XI11_7/XI0/XI0_45/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_10 XI11_7/net21_5_ xsel_45_ XI11_7/XI0/XI0_45/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_9 XI11_7/net21_6_ xsel_45_ XI11_7/XI0/XI0_45/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_8 XI11_7/net21_7_ xsel_45_ XI11_7/XI0/XI0_45/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_7 XI11_7/net21_8_ xsel_45_ XI11_7/XI0/XI0_45/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_6 XI11_7/net21_9_ xsel_45_ XI11_7/XI0/XI0_45/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_5 XI11_7/net21_10_ xsel_45_ XI11_7/XI0/XI0_45/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_4 XI11_7/net21_11_ xsel_45_ XI11_7/XI0/XI0_45/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_3 XI11_7/net21_12_ xsel_45_ XI11_7/XI0/XI0_45/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_2 XI11_7/net21_13_ xsel_45_ XI11_7/XI0/XI0_45/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_1 XI11_7/net21_14_ xsel_45_ XI11_7/XI0/XI0_45/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_0 XI11_7/net21_15_ xsel_45_ XI11_7/XI0/XI0_45/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_15 XI11_7/XI0/XI0_45/d__15_ xsel_45_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_14 XI11_7/XI0/XI0_45/d__14_ xsel_45_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_13 XI11_7/XI0/XI0_45/d__13_ xsel_45_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_12 XI11_7/XI0/XI0_45/d__12_ xsel_45_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_11 XI11_7/XI0/XI0_45/d__11_ xsel_45_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_10 XI11_7/XI0/XI0_45/d__10_ xsel_45_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_9 XI11_7/XI0/XI0_45/d__9_ xsel_45_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_8 XI11_7/XI0/XI0_45/d__8_ xsel_45_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_7 XI11_7/XI0/XI0_45/d__7_ xsel_45_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_6 XI11_7/XI0/XI0_45/d__6_ xsel_45_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_5 XI11_7/XI0/XI0_45/d__5_ xsel_45_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_4 XI11_7/XI0/XI0_45/d__4_ xsel_45_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_3 XI11_7/XI0/XI0_45/d__3_ xsel_45_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_2 XI11_7/XI0/XI0_45/d__2_ xsel_45_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_1 XI11_7/XI0/XI0_45/d__1_ xsel_45_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_0 XI11_7/XI0/XI0_45/d__0_ xsel_45_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_15 XI11_7/net21_0_ xsel_44_ XI11_7/XI0/XI0_44/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_14 XI11_7/net21_1_ xsel_44_ XI11_7/XI0/XI0_44/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_13 XI11_7/net21_2_ xsel_44_ XI11_7/XI0/XI0_44/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_12 XI11_7/net21_3_ xsel_44_ XI11_7/XI0/XI0_44/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_11 XI11_7/net21_4_ xsel_44_ XI11_7/XI0/XI0_44/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_10 XI11_7/net21_5_ xsel_44_ XI11_7/XI0/XI0_44/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_9 XI11_7/net21_6_ xsel_44_ XI11_7/XI0/XI0_44/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_8 XI11_7/net21_7_ xsel_44_ XI11_7/XI0/XI0_44/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_7 XI11_7/net21_8_ xsel_44_ XI11_7/XI0/XI0_44/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_6 XI11_7/net21_9_ xsel_44_ XI11_7/XI0/XI0_44/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_5 XI11_7/net21_10_ xsel_44_ XI11_7/XI0/XI0_44/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_4 XI11_7/net21_11_ xsel_44_ XI11_7/XI0/XI0_44/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_3 XI11_7/net21_12_ xsel_44_ XI11_7/XI0/XI0_44/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_2 XI11_7/net21_13_ xsel_44_ XI11_7/XI0/XI0_44/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_1 XI11_7/net21_14_ xsel_44_ XI11_7/XI0/XI0_44/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_0 XI11_7/net21_15_ xsel_44_ XI11_7/XI0/XI0_44/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_15 XI11_7/XI0/XI0_44/d__15_ xsel_44_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_14 XI11_7/XI0/XI0_44/d__14_ xsel_44_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_13 XI11_7/XI0/XI0_44/d__13_ xsel_44_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_12 XI11_7/XI0/XI0_44/d__12_ xsel_44_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_11 XI11_7/XI0/XI0_44/d__11_ xsel_44_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_10 XI11_7/XI0/XI0_44/d__10_ xsel_44_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_9 XI11_7/XI0/XI0_44/d__9_ xsel_44_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_8 XI11_7/XI0/XI0_44/d__8_ xsel_44_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_7 XI11_7/XI0/XI0_44/d__7_ xsel_44_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_6 XI11_7/XI0/XI0_44/d__6_ xsel_44_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_5 XI11_7/XI0/XI0_44/d__5_ xsel_44_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_4 XI11_7/XI0/XI0_44/d__4_ xsel_44_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_3 XI11_7/XI0/XI0_44/d__3_ xsel_44_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_2 XI11_7/XI0/XI0_44/d__2_ xsel_44_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_1 XI11_7/XI0/XI0_44/d__1_ xsel_44_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_0 XI11_7/XI0/XI0_44/d__0_ xsel_44_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_15 XI11_7/net21_0_ xsel_43_ XI11_7/XI0/XI0_43/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_14 XI11_7/net21_1_ xsel_43_ XI11_7/XI0/XI0_43/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_13 XI11_7/net21_2_ xsel_43_ XI11_7/XI0/XI0_43/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_12 XI11_7/net21_3_ xsel_43_ XI11_7/XI0/XI0_43/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_11 XI11_7/net21_4_ xsel_43_ XI11_7/XI0/XI0_43/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_10 XI11_7/net21_5_ xsel_43_ XI11_7/XI0/XI0_43/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_9 XI11_7/net21_6_ xsel_43_ XI11_7/XI0/XI0_43/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_8 XI11_7/net21_7_ xsel_43_ XI11_7/XI0/XI0_43/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_7 XI11_7/net21_8_ xsel_43_ XI11_7/XI0/XI0_43/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_6 XI11_7/net21_9_ xsel_43_ XI11_7/XI0/XI0_43/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_5 XI11_7/net21_10_ xsel_43_ XI11_7/XI0/XI0_43/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_4 XI11_7/net21_11_ xsel_43_ XI11_7/XI0/XI0_43/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_3 XI11_7/net21_12_ xsel_43_ XI11_7/XI0/XI0_43/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_2 XI11_7/net21_13_ xsel_43_ XI11_7/XI0/XI0_43/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_1 XI11_7/net21_14_ xsel_43_ XI11_7/XI0/XI0_43/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_0 XI11_7/net21_15_ xsel_43_ XI11_7/XI0/XI0_43/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_15 XI11_7/XI0/XI0_43/d__15_ xsel_43_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_14 XI11_7/XI0/XI0_43/d__14_ xsel_43_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_13 XI11_7/XI0/XI0_43/d__13_ xsel_43_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_12 XI11_7/XI0/XI0_43/d__12_ xsel_43_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_11 XI11_7/XI0/XI0_43/d__11_ xsel_43_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_10 XI11_7/XI0/XI0_43/d__10_ xsel_43_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_9 XI11_7/XI0/XI0_43/d__9_ xsel_43_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_8 XI11_7/XI0/XI0_43/d__8_ xsel_43_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_7 XI11_7/XI0/XI0_43/d__7_ xsel_43_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_6 XI11_7/XI0/XI0_43/d__6_ xsel_43_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_5 XI11_7/XI0/XI0_43/d__5_ xsel_43_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_4 XI11_7/XI0/XI0_43/d__4_ xsel_43_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_3 XI11_7/XI0/XI0_43/d__3_ xsel_43_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_2 XI11_7/XI0/XI0_43/d__2_ xsel_43_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_1 XI11_7/XI0/XI0_43/d__1_ xsel_43_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_0 XI11_7/XI0/XI0_43/d__0_ xsel_43_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_15 XI11_7/net21_0_ xsel_42_ XI11_7/XI0/XI0_42/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_14 XI11_7/net21_1_ xsel_42_ XI11_7/XI0/XI0_42/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_13 XI11_7/net21_2_ xsel_42_ XI11_7/XI0/XI0_42/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_12 XI11_7/net21_3_ xsel_42_ XI11_7/XI0/XI0_42/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_11 XI11_7/net21_4_ xsel_42_ XI11_7/XI0/XI0_42/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_10 XI11_7/net21_5_ xsel_42_ XI11_7/XI0/XI0_42/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_9 XI11_7/net21_6_ xsel_42_ XI11_7/XI0/XI0_42/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_8 XI11_7/net21_7_ xsel_42_ XI11_7/XI0/XI0_42/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_7 XI11_7/net21_8_ xsel_42_ XI11_7/XI0/XI0_42/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_6 XI11_7/net21_9_ xsel_42_ XI11_7/XI0/XI0_42/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_5 XI11_7/net21_10_ xsel_42_ XI11_7/XI0/XI0_42/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_4 XI11_7/net21_11_ xsel_42_ XI11_7/XI0/XI0_42/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_3 XI11_7/net21_12_ xsel_42_ XI11_7/XI0/XI0_42/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_2 XI11_7/net21_13_ xsel_42_ XI11_7/XI0/XI0_42/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_1 XI11_7/net21_14_ xsel_42_ XI11_7/XI0/XI0_42/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_0 XI11_7/net21_15_ xsel_42_ XI11_7/XI0/XI0_42/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_15 XI11_7/XI0/XI0_42/d__15_ xsel_42_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_14 XI11_7/XI0/XI0_42/d__14_ xsel_42_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_13 XI11_7/XI0/XI0_42/d__13_ xsel_42_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_12 XI11_7/XI0/XI0_42/d__12_ xsel_42_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_11 XI11_7/XI0/XI0_42/d__11_ xsel_42_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_10 XI11_7/XI0/XI0_42/d__10_ xsel_42_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_9 XI11_7/XI0/XI0_42/d__9_ xsel_42_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_8 XI11_7/XI0/XI0_42/d__8_ xsel_42_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_7 XI11_7/XI0/XI0_42/d__7_ xsel_42_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_6 XI11_7/XI0/XI0_42/d__6_ xsel_42_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_5 XI11_7/XI0/XI0_42/d__5_ xsel_42_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_4 XI11_7/XI0/XI0_42/d__4_ xsel_42_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_3 XI11_7/XI0/XI0_42/d__3_ xsel_42_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_2 XI11_7/XI0/XI0_42/d__2_ xsel_42_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_1 XI11_7/XI0/XI0_42/d__1_ xsel_42_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_0 XI11_7/XI0/XI0_42/d__0_ xsel_42_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_15 XI11_7/net21_0_ xsel_41_ XI11_7/XI0/XI0_41/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_14 XI11_7/net21_1_ xsel_41_ XI11_7/XI0/XI0_41/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_13 XI11_7/net21_2_ xsel_41_ XI11_7/XI0/XI0_41/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_12 XI11_7/net21_3_ xsel_41_ XI11_7/XI0/XI0_41/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_11 XI11_7/net21_4_ xsel_41_ XI11_7/XI0/XI0_41/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_10 XI11_7/net21_5_ xsel_41_ XI11_7/XI0/XI0_41/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_9 XI11_7/net21_6_ xsel_41_ XI11_7/XI0/XI0_41/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_8 XI11_7/net21_7_ xsel_41_ XI11_7/XI0/XI0_41/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_7 XI11_7/net21_8_ xsel_41_ XI11_7/XI0/XI0_41/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_6 XI11_7/net21_9_ xsel_41_ XI11_7/XI0/XI0_41/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_5 XI11_7/net21_10_ xsel_41_ XI11_7/XI0/XI0_41/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_4 XI11_7/net21_11_ xsel_41_ XI11_7/XI0/XI0_41/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_3 XI11_7/net21_12_ xsel_41_ XI11_7/XI0/XI0_41/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_2 XI11_7/net21_13_ xsel_41_ XI11_7/XI0/XI0_41/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_1 XI11_7/net21_14_ xsel_41_ XI11_7/XI0/XI0_41/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_0 XI11_7/net21_15_ xsel_41_ XI11_7/XI0/XI0_41/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_15 XI11_7/XI0/XI0_41/d__15_ xsel_41_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_14 XI11_7/XI0/XI0_41/d__14_ xsel_41_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_13 XI11_7/XI0/XI0_41/d__13_ xsel_41_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_12 XI11_7/XI0/XI0_41/d__12_ xsel_41_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_11 XI11_7/XI0/XI0_41/d__11_ xsel_41_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_10 XI11_7/XI0/XI0_41/d__10_ xsel_41_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_9 XI11_7/XI0/XI0_41/d__9_ xsel_41_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_8 XI11_7/XI0/XI0_41/d__8_ xsel_41_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_7 XI11_7/XI0/XI0_41/d__7_ xsel_41_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_6 XI11_7/XI0/XI0_41/d__6_ xsel_41_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_5 XI11_7/XI0/XI0_41/d__5_ xsel_41_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_4 XI11_7/XI0/XI0_41/d__4_ xsel_41_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_3 XI11_7/XI0/XI0_41/d__3_ xsel_41_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_2 XI11_7/XI0/XI0_41/d__2_ xsel_41_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_1 XI11_7/XI0/XI0_41/d__1_ xsel_41_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_0 XI11_7/XI0/XI0_41/d__0_ xsel_41_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_15 XI11_7/net21_0_ xsel_40_ XI11_7/XI0/XI0_40/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_14 XI11_7/net21_1_ xsel_40_ XI11_7/XI0/XI0_40/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_13 XI11_7/net21_2_ xsel_40_ XI11_7/XI0/XI0_40/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_12 XI11_7/net21_3_ xsel_40_ XI11_7/XI0/XI0_40/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_11 XI11_7/net21_4_ xsel_40_ XI11_7/XI0/XI0_40/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_10 XI11_7/net21_5_ xsel_40_ XI11_7/XI0/XI0_40/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_9 XI11_7/net21_6_ xsel_40_ XI11_7/XI0/XI0_40/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_8 XI11_7/net21_7_ xsel_40_ XI11_7/XI0/XI0_40/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_7 XI11_7/net21_8_ xsel_40_ XI11_7/XI0/XI0_40/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_6 XI11_7/net21_9_ xsel_40_ XI11_7/XI0/XI0_40/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_5 XI11_7/net21_10_ xsel_40_ XI11_7/XI0/XI0_40/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_4 XI11_7/net21_11_ xsel_40_ XI11_7/XI0/XI0_40/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_3 XI11_7/net21_12_ xsel_40_ XI11_7/XI0/XI0_40/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_2 XI11_7/net21_13_ xsel_40_ XI11_7/XI0/XI0_40/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_1 XI11_7/net21_14_ xsel_40_ XI11_7/XI0/XI0_40/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_0 XI11_7/net21_15_ xsel_40_ XI11_7/XI0/XI0_40/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_15 XI11_7/XI0/XI0_40/d__15_ xsel_40_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_14 XI11_7/XI0/XI0_40/d__14_ xsel_40_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_13 XI11_7/XI0/XI0_40/d__13_ xsel_40_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_12 XI11_7/XI0/XI0_40/d__12_ xsel_40_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_11 XI11_7/XI0/XI0_40/d__11_ xsel_40_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_10 XI11_7/XI0/XI0_40/d__10_ xsel_40_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_9 XI11_7/XI0/XI0_40/d__9_ xsel_40_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_8 XI11_7/XI0/XI0_40/d__8_ xsel_40_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_7 XI11_7/XI0/XI0_40/d__7_ xsel_40_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_6 XI11_7/XI0/XI0_40/d__6_ xsel_40_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_5 XI11_7/XI0/XI0_40/d__5_ xsel_40_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_4 XI11_7/XI0/XI0_40/d__4_ xsel_40_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_3 XI11_7/XI0/XI0_40/d__3_ xsel_40_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_2 XI11_7/XI0/XI0_40/d__2_ xsel_40_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_1 XI11_7/XI0/XI0_40/d__1_ xsel_40_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_0 XI11_7/XI0/XI0_40/d__0_ xsel_40_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_15 XI11_7/net21_0_ xsel_39_ XI11_7/XI0/XI0_39/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_14 XI11_7/net21_1_ xsel_39_ XI11_7/XI0/XI0_39/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_13 XI11_7/net21_2_ xsel_39_ XI11_7/XI0/XI0_39/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_12 XI11_7/net21_3_ xsel_39_ XI11_7/XI0/XI0_39/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_11 XI11_7/net21_4_ xsel_39_ XI11_7/XI0/XI0_39/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_10 XI11_7/net21_5_ xsel_39_ XI11_7/XI0/XI0_39/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_9 XI11_7/net21_6_ xsel_39_ XI11_7/XI0/XI0_39/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_8 XI11_7/net21_7_ xsel_39_ XI11_7/XI0/XI0_39/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_7 XI11_7/net21_8_ xsel_39_ XI11_7/XI0/XI0_39/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_6 XI11_7/net21_9_ xsel_39_ XI11_7/XI0/XI0_39/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_5 XI11_7/net21_10_ xsel_39_ XI11_7/XI0/XI0_39/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_4 XI11_7/net21_11_ xsel_39_ XI11_7/XI0/XI0_39/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_3 XI11_7/net21_12_ xsel_39_ XI11_7/XI0/XI0_39/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_2 XI11_7/net21_13_ xsel_39_ XI11_7/XI0/XI0_39/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_1 XI11_7/net21_14_ xsel_39_ XI11_7/XI0/XI0_39/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_0 XI11_7/net21_15_ xsel_39_ XI11_7/XI0/XI0_39/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_15 XI11_7/XI0/XI0_39/d__15_ xsel_39_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_14 XI11_7/XI0/XI0_39/d__14_ xsel_39_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_13 XI11_7/XI0/XI0_39/d__13_ xsel_39_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_12 XI11_7/XI0/XI0_39/d__12_ xsel_39_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_11 XI11_7/XI0/XI0_39/d__11_ xsel_39_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_10 XI11_7/XI0/XI0_39/d__10_ xsel_39_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_9 XI11_7/XI0/XI0_39/d__9_ xsel_39_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_8 XI11_7/XI0/XI0_39/d__8_ xsel_39_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_7 XI11_7/XI0/XI0_39/d__7_ xsel_39_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_6 XI11_7/XI0/XI0_39/d__6_ xsel_39_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_5 XI11_7/XI0/XI0_39/d__5_ xsel_39_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_4 XI11_7/XI0/XI0_39/d__4_ xsel_39_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_3 XI11_7/XI0/XI0_39/d__3_ xsel_39_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_2 XI11_7/XI0/XI0_39/d__2_ xsel_39_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_1 XI11_7/XI0/XI0_39/d__1_ xsel_39_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_0 XI11_7/XI0/XI0_39/d__0_ xsel_39_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_15 XI11_7/net21_0_ xsel_38_ XI11_7/XI0/XI0_38/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_14 XI11_7/net21_1_ xsel_38_ XI11_7/XI0/XI0_38/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_13 XI11_7/net21_2_ xsel_38_ XI11_7/XI0/XI0_38/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_12 XI11_7/net21_3_ xsel_38_ XI11_7/XI0/XI0_38/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_11 XI11_7/net21_4_ xsel_38_ XI11_7/XI0/XI0_38/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_10 XI11_7/net21_5_ xsel_38_ XI11_7/XI0/XI0_38/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_9 XI11_7/net21_6_ xsel_38_ XI11_7/XI0/XI0_38/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_8 XI11_7/net21_7_ xsel_38_ XI11_7/XI0/XI0_38/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_7 XI11_7/net21_8_ xsel_38_ XI11_7/XI0/XI0_38/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_6 XI11_7/net21_9_ xsel_38_ XI11_7/XI0/XI0_38/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_5 XI11_7/net21_10_ xsel_38_ XI11_7/XI0/XI0_38/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_4 XI11_7/net21_11_ xsel_38_ XI11_7/XI0/XI0_38/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_3 XI11_7/net21_12_ xsel_38_ XI11_7/XI0/XI0_38/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_2 XI11_7/net21_13_ xsel_38_ XI11_7/XI0/XI0_38/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_1 XI11_7/net21_14_ xsel_38_ XI11_7/XI0/XI0_38/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_0 XI11_7/net21_15_ xsel_38_ XI11_7/XI0/XI0_38/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_15 XI11_7/XI0/XI0_38/d__15_ xsel_38_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_14 XI11_7/XI0/XI0_38/d__14_ xsel_38_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_13 XI11_7/XI0/XI0_38/d__13_ xsel_38_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_12 XI11_7/XI0/XI0_38/d__12_ xsel_38_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_11 XI11_7/XI0/XI0_38/d__11_ xsel_38_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_10 XI11_7/XI0/XI0_38/d__10_ xsel_38_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_9 XI11_7/XI0/XI0_38/d__9_ xsel_38_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_8 XI11_7/XI0/XI0_38/d__8_ xsel_38_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_7 XI11_7/XI0/XI0_38/d__7_ xsel_38_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_6 XI11_7/XI0/XI0_38/d__6_ xsel_38_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_5 XI11_7/XI0/XI0_38/d__5_ xsel_38_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_4 XI11_7/XI0/XI0_38/d__4_ xsel_38_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_3 XI11_7/XI0/XI0_38/d__3_ xsel_38_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_2 XI11_7/XI0/XI0_38/d__2_ xsel_38_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_1 XI11_7/XI0/XI0_38/d__1_ xsel_38_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_0 XI11_7/XI0/XI0_38/d__0_ xsel_38_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_15 XI11_7/net21_0_ xsel_37_ XI11_7/XI0/XI0_37/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_14 XI11_7/net21_1_ xsel_37_ XI11_7/XI0/XI0_37/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_13 XI11_7/net21_2_ xsel_37_ XI11_7/XI0/XI0_37/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_12 XI11_7/net21_3_ xsel_37_ XI11_7/XI0/XI0_37/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_11 XI11_7/net21_4_ xsel_37_ XI11_7/XI0/XI0_37/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_10 XI11_7/net21_5_ xsel_37_ XI11_7/XI0/XI0_37/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_9 XI11_7/net21_6_ xsel_37_ XI11_7/XI0/XI0_37/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_8 XI11_7/net21_7_ xsel_37_ XI11_7/XI0/XI0_37/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_7 XI11_7/net21_8_ xsel_37_ XI11_7/XI0/XI0_37/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_6 XI11_7/net21_9_ xsel_37_ XI11_7/XI0/XI0_37/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_5 XI11_7/net21_10_ xsel_37_ XI11_7/XI0/XI0_37/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_4 XI11_7/net21_11_ xsel_37_ XI11_7/XI0/XI0_37/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_3 XI11_7/net21_12_ xsel_37_ XI11_7/XI0/XI0_37/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_2 XI11_7/net21_13_ xsel_37_ XI11_7/XI0/XI0_37/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_1 XI11_7/net21_14_ xsel_37_ XI11_7/XI0/XI0_37/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_0 XI11_7/net21_15_ xsel_37_ XI11_7/XI0/XI0_37/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_15 XI11_7/XI0/XI0_37/d__15_ xsel_37_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_14 XI11_7/XI0/XI0_37/d__14_ xsel_37_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_13 XI11_7/XI0/XI0_37/d__13_ xsel_37_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_12 XI11_7/XI0/XI0_37/d__12_ xsel_37_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_11 XI11_7/XI0/XI0_37/d__11_ xsel_37_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_10 XI11_7/XI0/XI0_37/d__10_ xsel_37_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_9 XI11_7/XI0/XI0_37/d__9_ xsel_37_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_8 XI11_7/XI0/XI0_37/d__8_ xsel_37_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_7 XI11_7/XI0/XI0_37/d__7_ xsel_37_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_6 XI11_7/XI0/XI0_37/d__6_ xsel_37_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_5 XI11_7/XI0/XI0_37/d__5_ xsel_37_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_4 XI11_7/XI0/XI0_37/d__4_ xsel_37_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_3 XI11_7/XI0/XI0_37/d__3_ xsel_37_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_2 XI11_7/XI0/XI0_37/d__2_ xsel_37_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_1 XI11_7/XI0/XI0_37/d__1_ xsel_37_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_0 XI11_7/XI0/XI0_37/d__0_ xsel_37_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_15 XI11_7/net21_0_ xsel_36_ XI11_7/XI0/XI0_36/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_14 XI11_7/net21_1_ xsel_36_ XI11_7/XI0/XI0_36/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_13 XI11_7/net21_2_ xsel_36_ XI11_7/XI0/XI0_36/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_12 XI11_7/net21_3_ xsel_36_ XI11_7/XI0/XI0_36/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_11 XI11_7/net21_4_ xsel_36_ XI11_7/XI0/XI0_36/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_10 XI11_7/net21_5_ xsel_36_ XI11_7/XI0/XI0_36/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_9 XI11_7/net21_6_ xsel_36_ XI11_7/XI0/XI0_36/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_8 XI11_7/net21_7_ xsel_36_ XI11_7/XI0/XI0_36/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_7 XI11_7/net21_8_ xsel_36_ XI11_7/XI0/XI0_36/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_6 XI11_7/net21_9_ xsel_36_ XI11_7/XI0/XI0_36/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_5 XI11_7/net21_10_ xsel_36_ XI11_7/XI0/XI0_36/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_4 XI11_7/net21_11_ xsel_36_ XI11_7/XI0/XI0_36/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_3 XI11_7/net21_12_ xsel_36_ XI11_7/XI0/XI0_36/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_2 XI11_7/net21_13_ xsel_36_ XI11_7/XI0/XI0_36/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_1 XI11_7/net21_14_ xsel_36_ XI11_7/XI0/XI0_36/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_0 XI11_7/net21_15_ xsel_36_ XI11_7/XI0/XI0_36/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_15 XI11_7/XI0/XI0_36/d__15_ xsel_36_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_14 XI11_7/XI0/XI0_36/d__14_ xsel_36_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_13 XI11_7/XI0/XI0_36/d__13_ xsel_36_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_12 XI11_7/XI0/XI0_36/d__12_ xsel_36_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_11 XI11_7/XI0/XI0_36/d__11_ xsel_36_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_10 XI11_7/XI0/XI0_36/d__10_ xsel_36_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_9 XI11_7/XI0/XI0_36/d__9_ xsel_36_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_8 XI11_7/XI0/XI0_36/d__8_ xsel_36_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_7 XI11_7/XI0/XI0_36/d__7_ xsel_36_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_6 XI11_7/XI0/XI0_36/d__6_ xsel_36_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_5 XI11_7/XI0/XI0_36/d__5_ xsel_36_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_4 XI11_7/XI0/XI0_36/d__4_ xsel_36_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_3 XI11_7/XI0/XI0_36/d__3_ xsel_36_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_2 XI11_7/XI0/XI0_36/d__2_ xsel_36_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_1 XI11_7/XI0/XI0_36/d__1_ xsel_36_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_0 XI11_7/XI0/XI0_36/d__0_ xsel_36_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_15 XI11_7/net21_0_ xsel_35_ XI11_7/XI0/XI0_35/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_14 XI11_7/net21_1_ xsel_35_ XI11_7/XI0/XI0_35/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_13 XI11_7/net21_2_ xsel_35_ XI11_7/XI0/XI0_35/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_12 XI11_7/net21_3_ xsel_35_ XI11_7/XI0/XI0_35/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_11 XI11_7/net21_4_ xsel_35_ XI11_7/XI0/XI0_35/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_10 XI11_7/net21_5_ xsel_35_ XI11_7/XI0/XI0_35/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_9 XI11_7/net21_6_ xsel_35_ XI11_7/XI0/XI0_35/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_8 XI11_7/net21_7_ xsel_35_ XI11_7/XI0/XI0_35/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_7 XI11_7/net21_8_ xsel_35_ XI11_7/XI0/XI0_35/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_6 XI11_7/net21_9_ xsel_35_ XI11_7/XI0/XI0_35/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_5 XI11_7/net21_10_ xsel_35_ XI11_7/XI0/XI0_35/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_4 XI11_7/net21_11_ xsel_35_ XI11_7/XI0/XI0_35/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_3 XI11_7/net21_12_ xsel_35_ XI11_7/XI0/XI0_35/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_2 XI11_7/net21_13_ xsel_35_ XI11_7/XI0/XI0_35/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_1 XI11_7/net21_14_ xsel_35_ XI11_7/XI0/XI0_35/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_0 XI11_7/net21_15_ xsel_35_ XI11_7/XI0/XI0_35/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_15 XI11_7/XI0/XI0_35/d__15_ xsel_35_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_14 XI11_7/XI0/XI0_35/d__14_ xsel_35_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_13 XI11_7/XI0/XI0_35/d__13_ xsel_35_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_12 XI11_7/XI0/XI0_35/d__12_ xsel_35_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_11 XI11_7/XI0/XI0_35/d__11_ xsel_35_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_10 XI11_7/XI0/XI0_35/d__10_ xsel_35_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_9 XI11_7/XI0/XI0_35/d__9_ xsel_35_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_8 XI11_7/XI0/XI0_35/d__8_ xsel_35_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_7 XI11_7/XI0/XI0_35/d__7_ xsel_35_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_6 XI11_7/XI0/XI0_35/d__6_ xsel_35_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_5 XI11_7/XI0/XI0_35/d__5_ xsel_35_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_4 XI11_7/XI0/XI0_35/d__4_ xsel_35_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_3 XI11_7/XI0/XI0_35/d__3_ xsel_35_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_2 XI11_7/XI0/XI0_35/d__2_ xsel_35_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_1 XI11_7/XI0/XI0_35/d__1_ xsel_35_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_0 XI11_7/XI0/XI0_35/d__0_ xsel_35_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_15 XI11_7/net21_0_ xsel_34_ XI11_7/XI0/XI0_34/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_14 XI11_7/net21_1_ xsel_34_ XI11_7/XI0/XI0_34/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_13 XI11_7/net21_2_ xsel_34_ XI11_7/XI0/XI0_34/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_12 XI11_7/net21_3_ xsel_34_ XI11_7/XI0/XI0_34/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_11 XI11_7/net21_4_ xsel_34_ XI11_7/XI0/XI0_34/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_10 XI11_7/net21_5_ xsel_34_ XI11_7/XI0/XI0_34/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_9 XI11_7/net21_6_ xsel_34_ XI11_7/XI0/XI0_34/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_8 XI11_7/net21_7_ xsel_34_ XI11_7/XI0/XI0_34/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_7 XI11_7/net21_8_ xsel_34_ XI11_7/XI0/XI0_34/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_6 XI11_7/net21_9_ xsel_34_ XI11_7/XI0/XI0_34/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_5 XI11_7/net21_10_ xsel_34_ XI11_7/XI0/XI0_34/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_4 XI11_7/net21_11_ xsel_34_ XI11_7/XI0/XI0_34/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_3 XI11_7/net21_12_ xsel_34_ XI11_7/XI0/XI0_34/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_2 XI11_7/net21_13_ xsel_34_ XI11_7/XI0/XI0_34/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_1 XI11_7/net21_14_ xsel_34_ XI11_7/XI0/XI0_34/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_0 XI11_7/net21_15_ xsel_34_ XI11_7/XI0/XI0_34/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_15 XI11_7/XI0/XI0_34/d__15_ xsel_34_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_14 XI11_7/XI0/XI0_34/d__14_ xsel_34_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_13 XI11_7/XI0/XI0_34/d__13_ xsel_34_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_12 XI11_7/XI0/XI0_34/d__12_ xsel_34_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_11 XI11_7/XI0/XI0_34/d__11_ xsel_34_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_10 XI11_7/XI0/XI0_34/d__10_ xsel_34_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_9 XI11_7/XI0/XI0_34/d__9_ xsel_34_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_8 XI11_7/XI0/XI0_34/d__8_ xsel_34_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_7 XI11_7/XI0/XI0_34/d__7_ xsel_34_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_6 XI11_7/XI0/XI0_34/d__6_ xsel_34_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_5 XI11_7/XI0/XI0_34/d__5_ xsel_34_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_4 XI11_7/XI0/XI0_34/d__4_ xsel_34_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_3 XI11_7/XI0/XI0_34/d__3_ xsel_34_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_2 XI11_7/XI0/XI0_34/d__2_ xsel_34_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_1 XI11_7/XI0/XI0_34/d__1_ xsel_34_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_0 XI11_7/XI0/XI0_34/d__0_ xsel_34_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_15 XI11_7/net21_0_ xsel_33_ XI11_7/XI0/XI0_33/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_14 XI11_7/net21_1_ xsel_33_ XI11_7/XI0/XI0_33/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_13 XI11_7/net21_2_ xsel_33_ XI11_7/XI0/XI0_33/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_12 XI11_7/net21_3_ xsel_33_ XI11_7/XI0/XI0_33/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_11 XI11_7/net21_4_ xsel_33_ XI11_7/XI0/XI0_33/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_10 XI11_7/net21_5_ xsel_33_ XI11_7/XI0/XI0_33/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_9 XI11_7/net21_6_ xsel_33_ XI11_7/XI0/XI0_33/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_8 XI11_7/net21_7_ xsel_33_ XI11_7/XI0/XI0_33/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_7 XI11_7/net21_8_ xsel_33_ XI11_7/XI0/XI0_33/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_6 XI11_7/net21_9_ xsel_33_ XI11_7/XI0/XI0_33/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_5 XI11_7/net21_10_ xsel_33_ XI11_7/XI0/XI0_33/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_4 XI11_7/net21_11_ xsel_33_ XI11_7/XI0/XI0_33/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_3 XI11_7/net21_12_ xsel_33_ XI11_7/XI0/XI0_33/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_2 XI11_7/net21_13_ xsel_33_ XI11_7/XI0/XI0_33/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_1 XI11_7/net21_14_ xsel_33_ XI11_7/XI0/XI0_33/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_0 XI11_7/net21_15_ xsel_33_ XI11_7/XI0/XI0_33/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_15 XI11_7/XI0/XI0_33/d__15_ xsel_33_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_14 XI11_7/XI0/XI0_33/d__14_ xsel_33_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_13 XI11_7/XI0/XI0_33/d__13_ xsel_33_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_12 XI11_7/XI0/XI0_33/d__12_ xsel_33_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_11 XI11_7/XI0/XI0_33/d__11_ xsel_33_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_10 XI11_7/XI0/XI0_33/d__10_ xsel_33_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_9 XI11_7/XI0/XI0_33/d__9_ xsel_33_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_8 XI11_7/XI0/XI0_33/d__8_ xsel_33_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_7 XI11_7/XI0/XI0_33/d__7_ xsel_33_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_6 XI11_7/XI0/XI0_33/d__6_ xsel_33_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_5 XI11_7/XI0/XI0_33/d__5_ xsel_33_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_4 XI11_7/XI0/XI0_33/d__4_ xsel_33_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_3 XI11_7/XI0/XI0_33/d__3_ xsel_33_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_2 XI11_7/XI0/XI0_33/d__2_ xsel_33_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_1 XI11_7/XI0/XI0_33/d__1_ xsel_33_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_0 XI11_7/XI0/XI0_33/d__0_ xsel_33_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_15 XI11_7/net21_0_ xsel_32_ XI11_7/XI0/XI0_32/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_14 XI11_7/net21_1_ xsel_32_ XI11_7/XI0/XI0_32/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_13 XI11_7/net21_2_ xsel_32_ XI11_7/XI0/XI0_32/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_12 XI11_7/net21_3_ xsel_32_ XI11_7/XI0/XI0_32/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_11 XI11_7/net21_4_ xsel_32_ XI11_7/XI0/XI0_32/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_10 XI11_7/net21_5_ xsel_32_ XI11_7/XI0/XI0_32/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_9 XI11_7/net21_6_ xsel_32_ XI11_7/XI0/XI0_32/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_8 XI11_7/net21_7_ xsel_32_ XI11_7/XI0/XI0_32/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_7 XI11_7/net21_8_ xsel_32_ XI11_7/XI0/XI0_32/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_6 XI11_7/net21_9_ xsel_32_ XI11_7/XI0/XI0_32/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_5 XI11_7/net21_10_ xsel_32_ XI11_7/XI0/XI0_32/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_4 XI11_7/net21_11_ xsel_32_ XI11_7/XI0/XI0_32/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_3 XI11_7/net21_12_ xsel_32_ XI11_7/XI0/XI0_32/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_2 XI11_7/net21_13_ xsel_32_ XI11_7/XI0/XI0_32/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_1 XI11_7/net21_14_ xsel_32_ XI11_7/XI0/XI0_32/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_0 XI11_7/net21_15_ xsel_32_ XI11_7/XI0/XI0_32/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_15 XI11_7/XI0/XI0_32/d__15_ xsel_32_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_14 XI11_7/XI0/XI0_32/d__14_ xsel_32_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_13 XI11_7/XI0/XI0_32/d__13_ xsel_32_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_12 XI11_7/XI0/XI0_32/d__12_ xsel_32_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_11 XI11_7/XI0/XI0_32/d__11_ xsel_32_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_10 XI11_7/XI0/XI0_32/d__10_ xsel_32_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_9 XI11_7/XI0/XI0_32/d__9_ xsel_32_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_8 XI11_7/XI0/XI0_32/d__8_ xsel_32_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_7 XI11_7/XI0/XI0_32/d__7_ xsel_32_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_6 XI11_7/XI0/XI0_32/d__6_ xsel_32_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_5 XI11_7/XI0/XI0_32/d__5_ xsel_32_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_4 XI11_7/XI0/XI0_32/d__4_ xsel_32_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_3 XI11_7/XI0/XI0_32/d__3_ xsel_32_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_2 XI11_7/XI0/XI0_32/d__2_ xsel_32_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_1 XI11_7/XI0/XI0_32/d__1_ xsel_32_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_0 XI11_7/XI0/XI0_32/d__0_ xsel_32_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_15 XI11_7/net21_0_ xsel_31_ XI11_7/XI0/XI0_31/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_14 XI11_7/net21_1_ xsel_31_ XI11_7/XI0/XI0_31/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_13 XI11_7/net21_2_ xsel_31_ XI11_7/XI0/XI0_31/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_12 XI11_7/net21_3_ xsel_31_ XI11_7/XI0/XI0_31/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_11 XI11_7/net21_4_ xsel_31_ XI11_7/XI0/XI0_31/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_10 XI11_7/net21_5_ xsel_31_ XI11_7/XI0/XI0_31/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_9 XI11_7/net21_6_ xsel_31_ XI11_7/XI0/XI0_31/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_8 XI11_7/net21_7_ xsel_31_ XI11_7/XI0/XI0_31/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_7 XI11_7/net21_8_ xsel_31_ XI11_7/XI0/XI0_31/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_6 XI11_7/net21_9_ xsel_31_ XI11_7/XI0/XI0_31/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_5 XI11_7/net21_10_ xsel_31_ XI11_7/XI0/XI0_31/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_4 XI11_7/net21_11_ xsel_31_ XI11_7/XI0/XI0_31/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_3 XI11_7/net21_12_ xsel_31_ XI11_7/XI0/XI0_31/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_2 XI11_7/net21_13_ xsel_31_ XI11_7/XI0/XI0_31/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_1 XI11_7/net21_14_ xsel_31_ XI11_7/XI0/XI0_31/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_0 XI11_7/net21_15_ xsel_31_ XI11_7/XI0/XI0_31/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_15 XI11_7/XI0/XI0_31/d__15_ xsel_31_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_14 XI11_7/XI0/XI0_31/d__14_ xsel_31_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_13 XI11_7/XI0/XI0_31/d__13_ xsel_31_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_12 XI11_7/XI0/XI0_31/d__12_ xsel_31_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_11 XI11_7/XI0/XI0_31/d__11_ xsel_31_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_10 XI11_7/XI0/XI0_31/d__10_ xsel_31_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_9 XI11_7/XI0/XI0_31/d__9_ xsel_31_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_8 XI11_7/XI0/XI0_31/d__8_ xsel_31_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_7 XI11_7/XI0/XI0_31/d__7_ xsel_31_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_6 XI11_7/XI0/XI0_31/d__6_ xsel_31_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_5 XI11_7/XI0/XI0_31/d__5_ xsel_31_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_4 XI11_7/XI0/XI0_31/d__4_ xsel_31_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_3 XI11_7/XI0/XI0_31/d__3_ xsel_31_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_2 XI11_7/XI0/XI0_31/d__2_ xsel_31_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_1 XI11_7/XI0/XI0_31/d__1_ xsel_31_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_0 XI11_7/XI0/XI0_31/d__0_ xsel_31_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_15 XI11_7/net21_0_ xsel_30_ XI11_7/XI0/XI0_30/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_14 XI11_7/net21_1_ xsel_30_ XI11_7/XI0/XI0_30/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_13 XI11_7/net21_2_ xsel_30_ XI11_7/XI0/XI0_30/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_12 XI11_7/net21_3_ xsel_30_ XI11_7/XI0/XI0_30/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_11 XI11_7/net21_4_ xsel_30_ XI11_7/XI0/XI0_30/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_10 XI11_7/net21_5_ xsel_30_ XI11_7/XI0/XI0_30/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_9 XI11_7/net21_6_ xsel_30_ XI11_7/XI0/XI0_30/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_8 XI11_7/net21_7_ xsel_30_ XI11_7/XI0/XI0_30/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_7 XI11_7/net21_8_ xsel_30_ XI11_7/XI0/XI0_30/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_6 XI11_7/net21_9_ xsel_30_ XI11_7/XI0/XI0_30/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_5 XI11_7/net21_10_ xsel_30_ XI11_7/XI0/XI0_30/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_4 XI11_7/net21_11_ xsel_30_ XI11_7/XI0/XI0_30/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_3 XI11_7/net21_12_ xsel_30_ XI11_7/XI0/XI0_30/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_2 XI11_7/net21_13_ xsel_30_ XI11_7/XI0/XI0_30/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_1 XI11_7/net21_14_ xsel_30_ XI11_7/XI0/XI0_30/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_0 XI11_7/net21_15_ xsel_30_ XI11_7/XI0/XI0_30/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_15 XI11_7/XI0/XI0_30/d__15_ xsel_30_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_14 XI11_7/XI0/XI0_30/d__14_ xsel_30_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_13 XI11_7/XI0/XI0_30/d__13_ xsel_30_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_12 XI11_7/XI0/XI0_30/d__12_ xsel_30_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_11 XI11_7/XI0/XI0_30/d__11_ xsel_30_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_10 XI11_7/XI0/XI0_30/d__10_ xsel_30_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_9 XI11_7/XI0/XI0_30/d__9_ xsel_30_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_8 XI11_7/XI0/XI0_30/d__8_ xsel_30_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_7 XI11_7/XI0/XI0_30/d__7_ xsel_30_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_6 XI11_7/XI0/XI0_30/d__6_ xsel_30_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_5 XI11_7/XI0/XI0_30/d__5_ xsel_30_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_4 XI11_7/XI0/XI0_30/d__4_ xsel_30_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_3 XI11_7/XI0/XI0_30/d__3_ xsel_30_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_2 XI11_7/XI0/XI0_30/d__2_ xsel_30_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_1 XI11_7/XI0/XI0_30/d__1_ xsel_30_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_0 XI11_7/XI0/XI0_30/d__0_ xsel_30_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_15 XI11_7/net21_0_ xsel_29_ XI11_7/XI0/XI0_29/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_14 XI11_7/net21_1_ xsel_29_ XI11_7/XI0/XI0_29/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_13 XI11_7/net21_2_ xsel_29_ XI11_7/XI0/XI0_29/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_12 XI11_7/net21_3_ xsel_29_ XI11_7/XI0/XI0_29/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_11 XI11_7/net21_4_ xsel_29_ XI11_7/XI0/XI0_29/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_10 XI11_7/net21_5_ xsel_29_ XI11_7/XI0/XI0_29/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_9 XI11_7/net21_6_ xsel_29_ XI11_7/XI0/XI0_29/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_8 XI11_7/net21_7_ xsel_29_ XI11_7/XI0/XI0_29/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_7 XI11_7/net21_8_ xsel_29_ XI11_7/XI0/XI0_29/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_6 XI11_7/net21_9_ xsel_29_ XI11_7/XI0/XI0_29/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_5 XI11_7/net21_10_ xsel_29_ XI11_7/XI0/XI0_29/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_4 XI11_7/net21_11_ xsel_29_ XI11_7/XI0/XI0_29/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_3 XI11_7/net21_12_ xsel_29_ XI11_7/XI0/XI0_29/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_2 XI11_7/net21_13_ xsel_29_ XI11_7/XI0/XI0_29/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_1 XI11_7/net21_14_ xsel_29_ XI11_7/XI0/XI0_29/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_0 XI11_7/net21_15_ xsel_29_ XI11_7/XI0/XI0_29/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_15 XI11_7/XI0/XI0_29/d__15_ xsel_29_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_14 XI11_7/XI0/XI0_29/d__14_ xsel_29_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_13 XI11_7/XI0/XI0_29/d__13_ xsel_29_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_12 XI11_7/XI0/XI0_29/d__12_ xsel_29_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_11 XI11_7/XI0/XI0_29/d__11_ xsel_29_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_10 XI11_7/XI0/XI0_29/d__10_ xsel_29_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_9 XI11_7/XI0/XI0_29/d__9_ xsel_29_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_8 XI11_7/XI0/XI0_29/d__8_ xsel_29_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_7 XI11_7/XI0/XI0_29/d__7_ xsel_29_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_6 XI11_7/XI0/XI0_29/d__6_ xsel_29_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_5 XI11_7/XI0/XI0_29/d__5_ xsel_29_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_4 XI11_7/XI0/XI0_29/d__4_ xsel_29_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_3 XI11_7/XI0/XI0_29/d__3_ xsel_29_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_2 XI11_7/XI0/XI0_29/d__2_ xsel_29_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_1 XI11_7/XI0/XI0_29/d__1_ xsel_29_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_0 XI11_7/XI0/XI0_29/d__0_ xsel_29_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_15 XI11_7/net21_0_ xsel_28_ XI11_7/XI0/XI0_28/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_14 XI11_7/net21_1_ xsel_28_ XI11_7/XI0/XI0_28/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_13 XI11_7/net21_2_ xsel_28_ XI11_7/XI0/XI0_28/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_12 XI11_7/net21_3_ xsel_28_ XI11_7/XI0/XI0_28/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_11 XI11_7/net21_4_ xsel_28_ XI11_7/XI0/XI0_28/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_10 XI11_7/net21_5_ xsel_28_ XI11_7/XI0/XI0_28/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_9 XI11_7/net21_6_ xsel_28_ XI11_7/XI0/XI0_28/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_8 XI11_7/net21_7_ xsel_28_ XI11_7/XI0/XI0_28/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_7 XI11_7/net21_8_ xsel_28_ XI11_7/XI0/XI0_28/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_6 XI11_7/net21_9_ xsel_28_ XI11_7/XI0/XI0_28/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_5 XI11_7/net21_10_ xsel_28_ XI11_7/XI0/XI0_28/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_4 XI11_7/net21_11_ xsel_28_ XI11_7/XI0/XI0_28/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_3 XI11_7/net21_12_ xsel_28_ XI11_7/XI0/XI0_28/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_2 XI11_7/net21_13_ xsel_28_ XI11_7/XI0/XI0_28/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_1 XI11_7/net21_14_ xsel_28_ XI11_7/XI0/XI0_28/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_0 XI11_7/net21_15_ xsel_28_ XI11_7/XI0/XI0_28/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_15 XI11_7/XI0/XI0_28/d__15_ xsel_28_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_14 XI11_7/XI0/XI0_28/d__14_ xsel_28_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_13 XI11_7/XI0/XI0_28/d__13_ xsel_28_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_12 XI11_7/XI0/XI0_28/d__12_ xsel_28_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_11 XI11_7/XI0/XI0_28/d__11_ xsel_28_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_10 XI11_7/XI0/XI0_28/d__10_ xsel_28_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_9 XI11_7/XI0/XI0_28/d__9_ xsel_28_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_8 XI11_7/XI0/XI0_28/d__8_ xsel_28_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_7 XI11_7/XI0/XI0_28/d__7_ xsel_28_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_6 XI11_7/XI0/XI0_28/d__6_ xsel_28_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_5 XI11_7/XI0/XI0_28/d__5_ xsel_28_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_4 XI11_7/XI0/XI0_28/d__4_ xsel_28_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_3 XI11_7/XI0/XI0_28/d__3_ xsel_28_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_2 XI11_7/XI0/XI0_28/d__2_ xsel_28_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_1 XI11_7/XI0/XI0_28/d__1_ xsel_28_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_0 XI11_7/XI0/XI0_28/d__0_ xsel_28_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_15 XI11_7/net21_0_ xsel_27_ XI11_7/XI0/XI0_27/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_14 XI11_7/net21_1_ xsel_27_ XI11_7/XI0/XI0_27/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_13 XI11_7/net21_2_ xsel_27_ XI11_7/XI0/XI0_27/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_12 XI11_7/net21_3_ xsel_27_ XI11_7/XI0/XI0_27/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_11 XI11_7/net21_4_ xsel_27_ XI11_7/XI0/XI0_27/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_10 XI11_7/net21_5_ xsel_27_ XI11_7/XI0/XI0_27/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_9 XI11_7/net21_6_ xsel_27_ XI11_7/XI0/XI0_27/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_8 XI11_7/net21_7_ xsel_27_ XI11_7/XI0/XI0_27/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_7 XI11_7/net21_8_ xsel_27_ XI11_7/XI0/XI0_27/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_6 XI11_7/net21_9_ xsel_27_ XI11_7/XI0/XI0_27/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_5 XI11_7/net21_10_ xsel_27_ XI11_7/XI0/XI0_27/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_4 XI11_7/net21_11_ xsel_27_ XI11_7/XI0/XI0_27/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_3 XI11_7/net21_12_ xsel_27_ XI11_7/XI0/XI0_27/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_2 XI11_7/net21_13_ xsel_27_ XI11_7/XI0/XI0_27/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_1 XI11_7/net21_14_ xsel_27_ XI11_7/XI0/XI0_27/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_0 XI11_7/net21_15_ xsel_27_ XI11_7/XI0/XI0_27/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_15 XI11_7/XI0/XI0_27/d__15_ xsel_27_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_14 XI11_7/XI0/XI0_27/d__14_ xsel_27_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_13 XI11_7/XI0/XI0_27/d__13_ xsel_27_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_12 XI11_7/XI0/XI0_27/d__12_ xsel_27_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_11 XI11_7/XI0/XI0_27/d__11_ xsel_27_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_10 XI11_7/XI0/XI0_27/d__10_ xsel_27_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_9 XI11_7/XI0/XI0_27/d__9_ xsel_27_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_8 XI11_7/XI0/XI0_27/d__8_ xsel_27_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_7 XI11_7/XI0/XI0_27/d__7_ xsel_27_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_6 XI11_7/XI0/XI0_27/d__6_ xsel_27_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_5 XI11_7/XI0/XI0_27/d__5_ xsel_27_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_4 XI11_7/XI0/XI0_27/d__4_ xsel_27_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_3 XI11_7/XI0/XI0_27/d__3_ xsel_27_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_2 XI11_7/XI0/XI0_27/d__2_ xsel_27_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_1 XI11_7/XI0/XI0_27/d__1_ xsel_27_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_0 XI11_7/XI0/XI0_27/d__0_ xsel_27_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_15 XI11_7/net21_0_ xsel_26_ XI11_7/XI0/XI0_26/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_14 XI11_7/net21_1_ xsel_26_ XI11_7/XI0/XI0_26/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_13 XI11_7/net21_2_ xsel_26_ XI11_7/XI0/XI0_26/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_12 XI11_7/net21_3_ xsel_26_ XI11_7/XI0/XI0_26/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_11 XI11_7/net21_4_ xsel_26_ XI11_7/XI0/XI0_26/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_10 XI11_7/net21_5_ xsel_26_ XI11_7/XI0/XI0_26/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_9 XI11_7/net21_6_ xsel_26_ XI11_7/XI0/XI0_26/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_8 XI11_7/net21_7_ xsel_26_ XI11_7/XI0/XI0_26/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_7 XI11_7/net21_8_ xsel_26_ XI11_7/XI0/XI0_26/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_6 XI11_7/net21_9_ xsel_26_ XI11_7/XI0/XI0_26/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_5 XI11_7/net21_10_ xsel_26_ XI11_7/XI0/XI0_26/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_4 XI11_7/net21_11_ xsel_26_ XI11_7/XI0/XI0_26/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_3 XI11_7/net21_12_ xsel_26_ XI11_7/XI0/XI0_26/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_2 XI11_7/net21_13_ xsel_26_ XI11_7/XI0/XI0_26/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_1 XI11_7/net21_14_ xsel_26_ XI11_7/XI0/XI0_26/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_0 XI11_7/net21_15_ xsel_26_ XI11_7/XI0/XI0_26/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_15 XI11_7/XI0/XI0_26/d__15_ xsel_26_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_14 XI11_7/XI0/XI0_26/d__14_ xsel_26_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_13 XI11_7/XI0/XI0_26/d__13_ xsel_26_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_12 XI11_7/XI0/XI0_26/d__12_ xsel_26_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_11 XI11_7/XI0/XI0_26/d__11_ xsel_26_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_10 XI11_7/XI0/XI0_26/d__10_ xsel_26_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_9 XI11_7/XI0/XI0_26/d__9_ xsel_26_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_8 XI11_7/XI0/XI0_26/d__8_ xsel_26_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_7 XI11_7/XI0/XI0_26/d__7_ xsel_26_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_6 XI11_7/XI0/XI0_26/d__6_ xsel_26_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_5 XI11_7/XI0/XI0_26/d__5_ xsel_26_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_4 XI11_7/XI0/XI0_26/d__4_ xsel_26_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_3 XI11_7/XI0/XI0_26/d__3_ xsel_26_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_2 XI11_7/XI0/XI0_26/d__2_ xsel_26_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_1 XI11_7/XI0/XI0_26/d__1_ xsel_26_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_0 XI11_7/XI0/XI0_26/d__0_ xsel_26_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_15 XI11_7/net21_0_ xsel_25_ XI11_7/XI0/XI0_25/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_14 XI11_7/net21_1_ xsel_25_ XI11_7/XI0/XI0_25/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_13 XI11_7/net21_2_ xsel_25_ XI11_7/XI0/XI0_25/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_12 XI11_7/net21_3_ xsel_25_ XI11_7/XI0/XI0_25/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_11 XI11_7/net21_4_ xsel_25_ XI11_7/XI0/XI0_25/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_10 XI11_7/net21_5_ xsel_25_ XI11_7/XI0/XI0_25/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_9 XI11_7/net21_6_ xsel_25_ XI11_7/XI0/XI0_25/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_8 XI11_7/net21_7_ xsel_25_ XI11_7/XI0/XI0_25/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_7 XI11_7/net21_8_ xsel_25_ XI11_7/XI0/XI0_25/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_6 XI11_7/net21_9_ xsel_25_ XI11_7/XI0/XI0_25/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_5 XI11_7/net21_10_ xsel_25_ XI11_7/XI0/XI0_25/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_4 XI11_7/net21_11_ xsel_25_ XI11_7/XI0/XI0_25/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_3 XI11_7/net21_12_ xsel_25_ XI11_7/XI0/XI0_25/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_2 XI11_7/net21_13_ xsel_25_ XI11_7/XI0/XI0_25/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_1 XI11_7/net21_14_ xsel_25_ XI11_7/XI0/XI0_25/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_0 XI11_7/net21_15_ xsel_25_ XI11_7/XI0/XI0_25/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_15 XI11_7/XI0/XI0_25/d__15_ xsel_25_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_14 XI11_7/XI0/XI0_25/d__14_ xsel_25_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_13 XI11_7/XI0/XI0_25/d__13_ xsel_25_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_12 XI11_7/XI0/XI0_25/d__12_ xsel_25_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_11 XI11_7/XI0/XI0_25/d__11_ xsel_25_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_10 XI11_7/XI0/XI0_25/d__10_ xsel_25_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_9 XI11_7/XI0/XI0_25/d__9_ xsel_25_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_8 XI11_7/XI0/XI0_25/d__8_ xsel_25_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_7 XI11_7/XI0/XI0_25/d__7_ xsel_25_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_6 XI11_7/XI0/XI0_25/d__6_ xsel_25_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_5 XI11_7/XI0/XI0_25/d__5_ xsel_25_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_4 XI11_7/XI0/XI0_25/d__4_ xsel_25_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_3 XI11_7/XI0/XI0_25/d__3_ xsel_25_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_2 XI11_7/XI0/XI0_25/d__2_ xsel_25_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_1 XI11_7/XI0/XI0_25/d__1_ xsel_25_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_0 XI11_7/XI0/XI0_25/d__0_ xsel_25_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_15 XI11_7/net21_0_ xsel_24_ XI11_7/XI0/XI0_24/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_14 XI11_7/net21_1_ xsel_24_ XI11_7/XI0/XI0_24/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_13 XI11_7/net21_2_ xsel_24_ XI11_7/XI0/XI0_24/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_12 XI11_7/net21_3_ xsel_24_ XI11_7/XI0/XI0_24/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_11 XI11_7/net21_4_ xsel_24_ XI11_7/XI0/XI0_24/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_10 XI11_7/net21_5_ xsel_24_ XI11_7/XI0/XI0_24/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_9 XI11_7/net21_6_ xsel_24_ XI11_7/XI0/XI0_24/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_8 XI11_7/net21_7_ xsel_24_ XI11_7/XI0/XI0_24/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_7 XI11_7/net21_8_ xsel_24_ XI11_7/XI0/XI0_24/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_6 XI11_7/net21_9_ xsel_24_ XI11_7/XI0/XI0_24/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_5 XI11_7/net21_10_ xsel_24_ XI11_7/XI0/XI0_24/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_4 XI11_7/net21_11_ xsel_24_ XI11_7/XI0/XI0_24/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_3 XI11_7/net21_12_ xsel_24_ XI11_7/XI0/XI0_24/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_2 XI11_7/net21_13_ xsel_24_ XI11_7/XI0/XI0_24/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_1 XI11_7/net21_14_ xsel_24_ XI11_7/XI0/XI0_24/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_0 XI11_7/net21_15_ xsel_24_ XI11_7/XI0/XI0_24/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_15 XI11_7/XI0/XI0_24/d__15_ xsel_24_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_14 XI11_7/XI0/XI0_24/d__14_ xsel_24_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_13 XI11_7/XI0/XI0_24/d__13_ xsel_24_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_12 XI11_7/XI0/XI0_24/d__12_ xsel_24_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_11 XI11_7/XI0/XI0_24/d__11_ xsel_24_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_10 XI11_7/XI0/XI0_24/d__10_ xsel_24_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_9 XI11_7/XI0/XI0_24/d__9_ xsel_24_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_8 XI11_7/XI0/XI0_24/d__8_ xsel_24_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_7 XI11_7/XI0/XI0_24/d__7_ xsel_24_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_6 XI11_7/XI0/XI0_24/d__6_ xsel_24_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_5 XI11_7/XI0/XI0_24/d__5_ xsel_24_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_4 XI11_7/XI0/XI0_24/d__4_ xsel_24_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_3 XI11_7/XI0/XI0_24/d__3_ xsel_24_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_2 XI11_7/XI0/XI0_24/d__2_ xsel_24_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_1 XI11_7/XI0/XI0_24/d__1_ xsel_24_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_0 XI11_7/XI0/XI0_24/d__0_ xsel_24_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_15 XI11_7/net21_0_ xsel_23_ XI11_7/XI0/XI0_23/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_14 XI11_7/net21_1_ xsel_23_ XI11_7/XI0/XI0_23/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_13 XI11_7/net21_2_ xsel_23_ XI11_7/XI0/XI0_23/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_12 XI11_7/net21_3_ xsel_23_ XI11_7/XI0/XI0_23/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_11 XI11_7/net21_4_ xsel_23_ XI11_7/XI0/XI0_23/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_10 XI11_7/net21_5_ xsel_23_ XI11_7/XI0/XI0_23/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_9 XI11_7/net21_6_ xsel_23_ XI11_7/XI0/XI0_23/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_8 XI11_7/net21_7_ xsel_23_ XI11_7/XI0/XI0_23/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_7 XI11_7/net21_8_ xsel_23_ XI11_7/XI0/XI0_23/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_6 XI11_7/net21_9_ xsel_23_ XI11_7/XI0/XI0_23/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_5 XI11_7/net21_10_ xsel_23_ XI11_7/XI0/XI0_23/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_4 XI11_7/net21_11_ xsel_23_ XI11_7/XI0/XI0_23/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_3 XI11_7/net21_12_ xsel_23_ XI11_7/XI0/XI0_23/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_2 XI11_7/net21_13_ xsel_23_ XI11_7/XI0/XI0_23/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_1 XI11_7/net21_14_ xsel_23_ XI11_7/XI0/XI0_23/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_0 XI11_7/net21_15_ xsel_23_ XI11_7/XI0/XI0_23/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_15 XI11_7/XI0/XI0_23/d__15_ xsel_23_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_14 XI11_7/XI0/XI0_23/d__14_ xsel_23_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_13 XI11_7/XI0/XI0_23/d__13_ xsel_23_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_12 XI11_7/XI0/XI0_23/d__12_ xsel_23_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_11 XI11_7/XI0/XI0_23/d__11_ xsel_23_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_10 XI11_7/XI0/XI0_23/d__10_ xsel_23_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_9 XI11_7/XI0/XI0_23/d__9_ xsel_23_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_8 XI11_7/XI0/XI0_23/d__8_ xsel_23_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_7 XI11_7/XI0/XI0_23/d__7_ xsel_23_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_6 XI11_7/XI0/XI0_23/d__6_ xsel_23_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_5 XI11_7/XI0/XI0_23/d__5_ xsel_23_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_4 XI11_7/XI0/XI0_23/d__4_ xsel_23_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_3 XI11_7/XI0/XI0_23/d__3_ xsel_23_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_2 XI11_7/XI0/XI0_23/d__2_ xsel_23_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_1 XI11_7/XI0/XI0_23/d__1_ xsel_23_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_0 XI11_7/XI0/XI0_23/d__0_ xsel_23_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_15 XI11_7/net21_0_ xsel_22_ XI11_7/XI0/XI0_22/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_14 XI11_7/net21_1_ xsel_22_ XI11_7/XI0/XI0_22/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_13 XI11_7/net21_2_ xsel_22_ XI11_7/XI0/XI0_22/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_12 XI11_7/net21_3_ xsel_22_ XI11_7/XI0/XI0_22/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_11 XI11_7/net21_4_ xsel_22_ XI11_7/XI0/XI0_22/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_10 XI11_7/net21_5_ xsel_22_ XI11_7/XI0/XI0_22/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_9 XI11_7/net21_6_ xsel_22_ XI11_7/XI0/XI0_22/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_8 XI11_7/net21_7_ xsel_22_ XI11_7/XI0/XI0_22/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_7 XI11_7/net21_8_ xsel_22_ XI11_7/XI0/XI0_22/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_6 XI11_7/net21_9_ xsel_22_ XI11_7/XI0/XI0_22/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_5 XI11_7/net21_10_ xsel_22_ XI11_7/XI0/XI0_22/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_4 XI11_7/net21_11_ xsel_22_ XI11_7/XI0/XI0_22/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_3 XI11_7/net21_12_ xsel_22_ XI11_7/XI0/XI0_22/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_2 XI11_7/net21_13_ xsel_22_ XI11_7/XI0/XI0_22/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_1 XI11_7/net21_14_ xsel_22_ XI11_7/XI0/XI0_22/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_0 XI11_7/net21_15_ xsel_22_ XI11_7/XI0/XI0_22/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_15 XI11_7/XI0/XI0_22/d__15_ xsel_22_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_14 XI11_7/XI0/XI0_22/d__14_ xsel_22_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_13 XI11_7/XI0/XI0_22/d__13_ xsel_22_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_12 XI11_7/XI0/XI0_22/d__12_ xsel_22_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_11 XI11_7/XI0/XI0_22/d__11_ xsel_22_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_10 XI11_7/XI0/XI0_22/d__10_ xsel_22_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_9 XI11_7/XI0/XI0_22/d__9_ xsel_22_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_8 XI11_7/XI0/XI0_22/d__8_ xsel_22_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_7 XI11_7/XI0/XI0_22/d__7_ xsel_22_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_6 XI11_7/XI0/XI0_22/d__6_ xsel_22_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_5 XI11_7/XI0/XI0_22/d__5_ xsel_22_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_4 XI11_7/XI0/XI0_22/d__4_ xsel_22_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_3 XI11_7/XI0/XI0_22/d__3_ xsel_22_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_2 XI11_7/XI0/XI0_22/d__2_ xsel_22_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_1 XI11_7/XI0/XI0_22/d__1_ xsel_22_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_0 XI11_7/XI0/XI0_22/d__0_ xsel_22_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_15 XI11_7/net21_0_ xsel_21_ XI11_7/XI0/XI0_21/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_14 XI11_7/net21_1_ xsel_21_ XI11_7/XI0/XI0_21/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_13 XI11_7/net21_2_ xsel_21_ XI11_7/XI0/XI0_21/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_12 XI11_7/net21_3_ xsel_21_ XI11_7/XI0/XI0_21/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_11 XI11_7/net21_4_ xsel_21_ XI11_7/XI0/XI0_21/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_10 XI11_7/net21_5_ xsel_21_ XI11_7/XI0/XI0_21/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_9 XI11_7/net21_6_ xsel_21_ XI11_7/XI0/XI0_21/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_8 XI11_7/net21_7_ xsel_21_ XI11_7/XI0/XI0_21/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_7 XI11_7/net21_8_ xsel_21_ XI11_7/XI0/XI0_21/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_6 XI11_7/net21_9_ xsel_21_ XI11_7/XI0/XI0_21/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_5 XI11_7/net21_10_ xsel_21_ XI11_7/XI0/XI0_21/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_4 XI11_7/net21_11_ xsel_21_ XI11_7/XI0/XI0_21/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_3 XI11_7/net21_12_ xsel_21_ XI11_7/XI0/XI0_21/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_2 XI11_7/net21_13_ xsel_21_ XI11_7/XI0/XI0_21/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_1 XI11_7/net21_14_ xsel_21_ XI11_7/XI0/XI0_21/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_0 XI11_7/net21_15_ xsel_21_ XI11_7/XI0/XI0_21/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_15 XI11_7/XI0/XI0_21/d__15_ xsel_21_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_14 XI11_7/XI0/XI0_21/d__14_ xsel_21_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_13 XI11_7/XI0/XI0_21/d__13_ xsel_21_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_12 XI11_7/XI0/XI0_21/d__12_ xsel_21_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_11 XI11_7/XI0/XI0_21/d__11_ xsel_21_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_10 XI11_7/XI0/XI0_21/d__10_ xsel_21_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_9 XI11_7/XI0/XI0_21/d__9_ xsel_21_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_8 XI11_7/XI0/XI0_21/d__8_ xsel_21_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_7 XI11_7/XI0/XI0_21/d__7_ xsel_21_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_6 XI11_7/XI0/XI0_21/d__6_ xsel_21_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_5 XI11_7/XI0/XI0_21/d__5_ xsel_21_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_4 XI11_7/XI0/XI0_21/d__4_ xsel_21_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_3 XI11_7/XI0/XI0_21/d__3_ xsel_21_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_2 XI11_7/XI0/XI0_21/d__2_ xsel_21_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_1 XI11_7/XI0/XI0_21/d__1_ xsel_21_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_0 XI11_7/XI0/XI0_21/d__0_ xsel_21_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_15 XI11_7/net21_0_ xsel_20_ XI11_7/XI0/XI0_20/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_14 XI11_7/net21_1_ xsel_20_ XI11_7/XI0/XI0_20/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_13 XI11_7/net21_2_ xsel_20_ XI11_7/XI0/XI0_20/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_12 XI11_7/net21_3_ xsel_20_ XI11_7/XI0/XI0_20/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_11 XI11_7/net21_4_ xsel_20_ XI11_7/XI0/XI0_20/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_10 XI11_7/net21_5_ xsel_20_ XI11_7/XI0/XI0_20/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_9 XI11_7/net21_6_ xsel_20_ XI11_7/XI0/XI0_20/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_8 XI11_7/net21_7_ xsel_20_ XI11_7/XI0/XI0_20/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_7 XI11_7/net21_8_ xsel_20_ XI11_7/XI0/XI0_20/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_6 XI11_7/net21_9_ xsel_20_ XI11_7/XI0/XI0_20/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_5 XI11_7/net21_10_ xsel_20_ XI11_7/XI0/XI0_20/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_4 XI11_7/net21_11_ xsel_20_ XI11_7/XI0/XI0_20/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_3 XI11_7/net21_12_ xsel_20_ XI11_7/XI0/XI0_20/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_2 XI11_7/net21_13_ xsel_20_ XI11_7/XI0/XI0_20/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_1 XI11_7/net21_14_ xsel_20_ XI11_7/XI0/XI0_20/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_0 XI11_7/net21_15_ xsel_20_ XI11_7/XI0/XI0_20/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_15 XI11_7/XI0/XI0_20/d__15_ xsel_20_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_14 XI11_7/XI0/XI0_20/d__14_ xsel_20_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_13 XI11_7/XI0/XI0_20/d__13_ xsel_20_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_12 XI11_7/XI0/XI0_20/d__12_ xsel_20_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_11 XI11_7/XI0/XI0_20/d__11_ xsel_20_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_10 XI11_7/XI0/XI0_20/d__10_ xsel_20_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_9 XI11_7/XI0/XI0_20/d__9_ xsel_20_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_8 XI11_7/XI0/XI0_20/d__8_ xsel_20_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_7 XI11_7/XI0/XI0_20/d__7_ xsel_20_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_6 XI11_7/XI0/XI0_20/d__6_ xsel_20_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_5 XI11_7/XI0/XI0_20/d__5_ xsel_20_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_4 XI11_7/XI0/XI0_20/d__4_ xsel_20_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_3 XI11_7/XI0/XI0_20/d__3_ xsel_20_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_2 XI11_7/XI0/XI0_20/d__2_ xsel_20_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_1 XI11_7/XI0/XI0_20/d__1_ xsel_20_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_0 XI11_7/XI0/XI0_20/d__0_ xsel_20_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_15 XI11_7/net21_0_ xsel_19_ XI11_7/XI0/XI0_19/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_14 XI11_7/net21_1_ xsel_19_ XI11_7/XI0/XI0_19/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_13 XI11_7/net21_2_ xsel_19_ XI11_7/XI0/XI0_19/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_12 XI11_7/net21_3_ xsel_19_ XI11_7/XI0/XI0_19/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_11 XI11_7/net21_4_ xsel_19_ XI11_7/XI0/XI0_19/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_10 XI11_7/net21_5_ xsel_19_ XI11_7/XI0/XI0_19/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_9 XI11_7/net21_6_ xsel_19_ XI11_7/XI0/XI0_19/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_8 XI11_7/net21_7_ xsel_19_ XI11_7/XI0/XI0_19/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_7 XI11_7/net21_8_ xsel_19_ XI11_7/XI0/XI0_19/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_6 XI11_7/net21_9_ xsel_19_ XI11_7/XI0/XI0_19/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_5 XI11_7/net21_10_ xsel_19_ XI11_7/XI0/XI0_19/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_4 XI11_7/net21_11_ xsel_19_ XI11_7/XI0/XI0_19/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_3 XI11_7/net21_12_ xsel_19_ XI11_7/XI0/XI0_19/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_2 XI11_7/net21_13_ xsel_19_ XI11_7/XI0/XI0_19/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_1 XI11_7/net21_14_ xsel_19_ XI11_7/XI0/XI0_19/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_0 XI11_7/net21_15_ xsel_19_ XI11_7/XI0/XI0_19/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_15 XI11_7/XI0/XI0_19/d__15_ xsel_19_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_14 XI11_7/XI0/XI0_19/d__14_ xsel_19_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_13 XI11_7/XI0/XI0_19/d__13_ xsel_19_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_12 XI11_7/XI0/XI0_19/d__12_ xsel_19_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_11 XI11_7/XI0/XI0_19/d__11_ xsel_19_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_10 XI11_7/XI0/XI0_19/d__10_ xsel_19_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_9 XI11_7/XI0/XI0_19/d__9_ xsel_19_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_8 XI11_7/XI0/XI0_19/d__8_ xsel_19_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_7 XI11_7/XI0/XI0_19/d__7_ xsel_19_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_6 XI11_7/XI0/XI0_19/d__6_ xsel_19_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_5 XI11_7/XI0/XI0_19/d__5_ xsel_19_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_4 XI11_7/XI0/XI0_19/d__4_ xsel_19_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_3 XI11_7/XI0/XI0_19/d__3_ xsel_19_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_2 XI11_7/XI0/XI0_19/d__2_ xsel_19_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_1 XI11_7/XI0/XI0_19/d__1_ xsel_19_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_0 XI11_7/XI0/XI0_19/d__0_ xsel_19_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_15 XI11_7/net21_0_ xsel_18_ XI11_7/XI0/XI0_18/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_14 XI11_7/net21_1_ xsel_18_ XI11_7/XI0/XI0_18/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_13 XI11_7/net21_2_ xsel_18_ XI11_7/XI0/XI0_18/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_12 XI11_7/net21_3_ xsel_18_ XI11_7/XI0/XI0_18/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_11 XI11_7/net21_4_ xsel_18_ XI11_7/XI0/XI0_18/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_10 XI11_7/net21_5_ xsel_18_ XI11_7/XI0/XI0_18/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_9 XI11_7/net21_6_ xsel_18_ XI11_7/XI0/XI0_18/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_8 XI11_7/net21_7_ xsel_18_ XI11_7/XI0/XI0_18/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_7 XI11_7/net21_8_ xsel_18_ XI11_7/XI0/XI0_18/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_6 XI11_7/net21_9_ xsel_18_ XI11_7/XI0/XI0_18/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_5 XI11_7/net21_10_ xsel_18_ XI11_7/XI0/XI0_18/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_4 XI11_7/net21_11_ xsel_18_ XI11_7/XI0/XI0_18/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_3 XI11_7/net21_12_ xsel_18_ XI11_7/XI0/XI0_18/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_2 XI11_7/net21_13_ xsel_18_ XI11_7/XI0/XI0_18/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_1 XI11_7/net21_14_ xsel_18_ XI11_7/XI0/XI0_18/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_0 XI11_7/net21_15_ xsel_18_ XI11_7/XI0/XI0_18/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_15 XI11_7/XI0/XI0_18/d__15_ xsel_18_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_14 XI11_7/XI0/XI0_18/d__14_ xsel_18_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_13 XI11_7/XI0/XI0_18/d__13_ xsel_18_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_12 XI11_7/XI0/XI0_18/d__12_ xsel_18_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_11 XI11_7/XI0/XI0_18/d__11_ xsel_18_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_10 XI11_7/XI0/XI0_18/d__10_ xsel_18_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_9 XI11_7/XI0/XI0_18/d__9_ xsel_18_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_8 XI11_7/XI0/XI0_18/d__8_ xsel_18_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_7 XI11_7/XI0/XI0_18/d__7_ xsel_18_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_6 XI11_7/XI0/XI0_18/d__6_ xsel_18_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_5 XI11_7/XI0/XI0_18/d__5_ xsel_18_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_4 XI11_7/XI0/XI0_18/d__4_ xsel_18_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_3 XI11_7/XI0/XI0_18/d__3_ xsel_18_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_2 XI11_7/XI0/XI0_18/d__2_ xsel_18_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_1 XI11_7/XI0/XI0_18/d__1_ xsel_18_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_0 XI11_7/XI0/XI0_18/d__0_ xsel_18_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_15 XI11_7/net21_0_ xsel_17_ XI11_7/XI0/XI0_17/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_14 XI11_7/net21_1_ xsel_17_ XI11_7/XI0/XI0_17/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_13 XI11_7/net21_2_ xsel_17_ XI11_7/XI0/XI0_17/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_12 XI11_7/net21_3_ xsel_17_ XI11_7/XI0/XI0_17/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_11 XI11_7/net21_4_ xsel_17_ XI11_7/XI0/XI0_17/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_10 XI11_7/net21_5_ xsel_17_ XI11_7/XI0/XI0_17/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_9 XI11_7/net21_6_ xsel_17_ XI11_7/XI0/XI0_17/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_8 XI11_7/net21_7_ xsel_17_ XI11_7/XI0/XI0_17/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_7 XI11_7/net21_8_ xsel_17_ XI11_7/XI0/XI0_17/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_6 XI11_7/net21_9_ xsel_17_ XI11_7/XI0/XI0_17/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_5 XI11_7/net21_10_ xsel_17_ XI11_7/XI0/XI0_17/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_4 XI11_7/net21_11_ xsel_17_ XI11_7/XI0/XI0_17/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_3 XI11_7/net21_12_ xsel_17_ XI11_7/XI0/XI0_17/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_2 XI11_7/net21_13_ xsel_17_ XI11_7/XI0/XI0_17/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_1 XI11_7/net21_14_ xsel_17_ XI11_7/XI0/XI0_17/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_0 XI11_7/net21_15_ xsel_17_ XI11_7/XI0/XI0_17/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_15 XI11_7/XI0/XI0_17/d__15_ xsel_17_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_14 XI11_7/XI0/XI0_17/d__14_ xsel_17_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_13 XI11_7/XI0/XI0_17/d__13_ xsel_17_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_12 XI11_7/XI0/XI0_17/d__12_ xsel_17_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_11 XI11_7/XI0/XI0_17/d__11_ xsel_17_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_10 XI11_7/XI0/XI0_17/d__10_ xsel_17_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_9 XI11_7/XI0/XI0_17/d__9_ xsel_17_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_8 XI11_7/XI0/XI0_17/d__8_ xsel_17_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_7 XI11_7/XI0/XI0_17/d__7_ xsel_17_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_6 XI11_7/XI0/XI0_17/d__6_ xsel_17_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_5 XI11_7/XI0/XI0_17/d__5_ xsel_17_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_4 XI11_7/XI0/XI0_17/d__4_ xsel_17_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_3 XI11_7/XI0/XI0_17/d__3_ xsel_17_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_2 XI11_7/XI0/XI0_17/d__2_ xsel_17_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_1 XI11_7/XI0/XI0_17/d__1_ xsel_17_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_0 XI11_7/XI0/XI0_17/d__0_ xsel_17_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_15 XI11_7/net21_0_ xsel_16_ XI11_7/XI0/XI0_16/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_14 XI11_7/net21_1_ xsel_16_ XI11_7/XI0/XI0_16/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_13 XI11_7/net21_2_ xsel_16_ XI11_7/XI0/XI0_16/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_12 XI11_7/net21_3_ xsel_16_ XI11_7/XI0/XI0_16/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_11 XI11_7/net21_4_ xsel_16_ XI11_7/XI0/XI0_16/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_10 XI11_7/net21_5_ xsel_16_ XI11_7/XI0/XI0_16/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_9 XI11_7/net21_6_ xsel_16_ XI11_7/XI0/XI0_16/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_8 XI11_7/net21_7_ xsel_16_ XI11_7/XI0/XI0_16/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_7 XI11_7/net21_8_ xsel_16_ XI11_7/XI0/XI0_16/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_6 XI11_7/net21_9_ xsel_16_ XI11_7/XI0/XI0_16/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_5 XI11_7/net21_10_ xsel_16_ XI11_7/XI0/XI0_16/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_4 XI11_7/net21_11_ xsel_16_ XI11_7/XI0/XI0_16/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_3 XI11_7/net21_12_ xsel_16_ XI11_7/XI0/XI0_16/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_2 XI11_7/net21_13_ xsel_16_ XI11_7/XI0/XI0_16/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_1 XI11_7/net21_14_ xsel_16_ XI11_7/XI0/XI0_16/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_0 XI11_7/net21_15_ xsel_16_ XI11_7/XI0/XI0_16/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_15 XI11_7/XI0/XI0_16/d__15_ xsel_16_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_14 XI11_7/XI0/XI0_16/d__14_ xsel_16_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_13 XI11_7/XI0/XI0_16/d__13_ xsel_16_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_12 XI11_7/XI0/XI0_16/d__12_ xsel_16_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_11 XI11_7/XI0/XI0_16/d__11_ xsel_16_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_10 XI11_7/XI0/XI0_16/d__10_ xsel_16_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_9 XI11_7/XI0/XI0_16/d__9_ xsel_16_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_8 XI11_7/XI0/XI0_16/d__8_ xsel_16_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_7 XI11_7/XI0/XI0_16/d__7_ xsel_16_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_6 XI11_7/XI0/XI0_16/d__6_ xsel_16_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_5 XI11_7/XI0/XI0_16/d__5_ xsel_16_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_4 XI11_7/XI0/XI0_16/d__4_ xsel_16_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_3 XI11_7/XI0/XI0_16/d__3_ xsel_16_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_2 XI11_7/XI0/XI0_16/d__2_ xsel_16_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_1 XI11_7/XI0/XI0_16/d__1_ xsel_16_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_0 XI11_7/XI0/XI0_16/d__0_ xsel_16_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_15 XI11_7/net21_0_ xsel_15_ XI11_7/XI0/XI0_15/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_14 XI11_7/net21_1_ xsel_15_ XI11_7/XI0/XI0_15/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_13 XI11_7/net21_2_ xsel_15_ XI11_7/XI0/XI0_15/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_12 XI11_7/net21_3_ xsel_15_ XI11_7/XI0/XI0_15/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_11 XI11_7/net21_4_ xsel_15_ XI11_7/XI0/XI0_15/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_10 XI11_7/net21_5_ xsel_15_ XI11_7/XI0/XI0_15/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_9 XI11_7/net21_6_ xsel_15_ XI11_7/XI0/XI0_15/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_8 XI11_7/net21_7_ xsel_15_ XI11_7/XI0/XI0_15/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_7 XI11_7/net21_8_ xsel_15_ XI11_7/XI0/XI0_15/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_6 XI11_7/net21_9_ xsel_15_ XI11_7/XI0/XI0_15/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_5 XI11_7/net21_10_ xsel_15_ XI11_7/XI0/XI0_15/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_4 XI11_7/net21_11_ xsel_15_ XI11_7/XI0/XI0_15/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_3 XI11_7/net21_12_ xsel_15_ XI11_7/XI0/XI0_15/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_2 XI11_7/net21_13_ xsel_15_ XI11_7/XI0/XI0_15/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_1 XI11_7/net21_14_ xsel_15_ XI11_7/XI0/XI0_15/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_0 XI11_7/net21_15_ xsel_15_ XI11_7/XI0/XI0_15/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_15 XI11_7/XI0/XI0_15/d__15_ xsel_15_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_14 XI11_7/XI0/XI0_15/d__14_ xsel_15_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_13 XI11_7/XI0/XI0_15/d__13_ xsel_15_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_12 XI11_7/XI0/XI0_15/d__12_ xsel_15_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_11 XI11_7/XI0/XI0_15/d__11_ xsel_15_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_10 XI11_7/XI0/XI0_15/d__10_ xsel_15_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_9 XI11_7/XI0/XI0_15/d__9_ xsel_15_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_8 XI11_7/XI0/XI0_15/d__8_ xsel_15_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_7 XI11_7/XI0/XI0_15/d__7_ xsel_15_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_6 XI11_7/XI0/XI0_15/d__6_ xsel_15_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_5 XI11_7/XI0/XI0_15/d__5_ xsel_15_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_4 XI11_7/XI0/XI0_15/d__4_ xsel_15_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_3 XI11_7/XI0/XI0_15/d__3_ xsel_15_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_2 XI11_7/XI0/XI0_15/d__2_ xsel_15_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_1 XI11_7/XI0/XI0_15/d__1_ xsel_15_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_0 XI11_7/XI0/XI0_15/d__0_ xsel_15_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_15 XI11_7/net21_0_ xsel_14_ XI11_7/XI0/XI0_14/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_14 XI11_7/net21_1_ xsel_14_ XI11_7/XI0/XI0_14/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_13 XI11_7/net21_2_ xsel_14_ XI11_7/XI0/XI0_14/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_12 XI11_7/net21_3_ xsel_14_ XI11_7/XI0/XI0_14/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_11 XI11_7/net21_4_ xsel_14_ XI11_7/XI0/XI0_14/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_10 XI11_7/net21_5_ xsel_14_ XI11_7/XI0/XI0_14/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_9 XI11_7/net21_6_ xsel_14_ XI11_7/XI0/XI0_14/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_8 XI11_7/net21_7_ xsel_14_ XI11_7/XI0/XI0_14/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_7 XI11_7/net21_8_ xsel_14_ XI11_7/XI0/XI0_14/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_6 XI11_7/net21_9_ xsel_14_ XI11_7/XI0/XI0_14/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_5 XI11_7/net21_10_ xsel_14_ XI11_7/XI0/XI0_14/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_4 XI11_7/net21_11_ xsel_14_ XI11_7/XI0/XI0_14/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_3 XI11_7/net21_12_ xsel_14_ XI11_7/XI0/XI0_14/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_2 XI11_7/net21_13_ xsel_14_ XI11_7/XI0/XI0_14/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_1 XI11_7/net21_14_ xsel_14_ XI11_7/XI0/XI0_14/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_0 XI11_7/net21_15_ xsel_14_ XI11_7/XI0/XI0_14/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_15 XI11_7/XI0/XI0_14/d__15_ xsel_14_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_14 XI11_7/XI0/XI0_14/d__14_ xsel_14_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_13 XI11_7/XI0/XI0_14/d__13_ xsel_14_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_12 XI11_7/XI0/XI0_14/d__12_ xsel_14_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_11 XI11_7/XI0/XI0_14/d__11_ xsel_14_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_10 XI11_7/XI0/XI0_14/d__10_ xsel_14_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_9 XI11_7/XI0/XI0_14/d__9_ xsel_14_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_8 XI11_7/XI0/XI0_14/d__8_ xsel_14_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_7 XI11_7/XI0/XI0_14/d__7_ xsel_14_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_6 XI11_7/XI0/XI0_14/d__6_ xsel_14_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_5 XI11_7/XI0/XI0_14/d__5_ xsel_14_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_4 XI11_7/XI0/XI0_14/d__4_ xsel_14_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_3 XI11_7/XI0/XI0_14/d__3_ xsel_14_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_2 XI11_7/XI0/XI0_14/d__2_ xsel_14_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_1 XI11_7/XI0/XI0_14/d__1_ xsel_14_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_0 XI11_7/XI0/XI0_14/d__0_ xsel_14_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_15 XI11_7/net21_0_ xsel_13_ XI11_7/XI0/XI0_13/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_14 XI11_7/net21_1_ xsel_13_ XI11_7/XI0/XI0_13/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_13 XI11_7/net21_2_ xsel_13_ XI11_7/XI0/XI0_13/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_12 XI11_7/net21_3_ xsel_13_ XI11_7/XI0/XI0_13/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_11 XI11_7/net21_4_ xsel_13_ XI11_7/XI0/XI0_13/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_10 XI11_7/net21_5_ xsel_13_ XI11_7/XI0/XI0_13/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_9 XI11_7/net21_6_ xsel_13_ XI11_7/XI0/XI0_13/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_8 XI11_7/net21_7_ xsel_13_ XI11_7/XI0/XI0_13/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_7 XI11_7/net21_8_ xsel_13_ XI11_7/XI0/XI0_13/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_6 XI11_7/net21_9_ xsel_13_ XI11_7/XI0/XI0_13/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_5 XI11_7/net21_10_ xsel_13_ XI11_7/XI0/XI0_13/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_4 XI11_7/net21_11_ xsel_13_ XI11_7/XI0/XI0_13/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_3 XI11_7/net21_12_ xsel_13_ XI11_7/XI0/XI0_13/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_2 XI11_7/net21_13_ xsel_13_ XI11_7/XI0/XI0_13/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_1 XI11_7/net21_14_ xsel_13_ XI11_7/XI0/XI0_13/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_0 XI11_7/net21_15_ xsel_13_ XI11_7/XI0/XI0_13/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_15 XI11_7/XI0/XI0_13/d__15_ xsel_13_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_14 XI11_7/XI0/XI0_13/d__14_ xsel_13_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_13 XI11_7/XI0/XI0_13/d__13_ xsel_13_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_12 XI11_7/XI0/XI0_13/d__12_ xsel_13_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_11 XI11_7/XI0/XI0_13/d__11_ xsel_13_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_10 XI11_7/XI0/XI0_13/d__10_ xsel_13_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_9 XI11_7/XI0/XI0_13/d__9_ xsel_13_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_8 XI11_7/XI0/XI0_13/d__8_ xsel_13_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_7 XI11_7/XI0/XI0_13/d__7_ xsel_13_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_6 XI11_7/XI0/XI0_13/d__6_ xsel_13_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_5 XI11_7/XI0/XI0_13/d__5_ xsel_13_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_4 XI11_7/XI0/XI0_13/d__4_ xsel_13_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_3 XI11_7/XI0/XI0_13/d__3_ xsel_13_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_2 XI11_7/XI0/XI0_13/d__2_ xsel_13_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_1 XI11_7/XI0/XI0_13/d__1_ xsel_13_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_0 XI11_7/XI0/XI0_13/d__0_ xsel_13_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_15 XI11_7/net21_0_ xsel_12_ XI11_7/XI0/XI0_12/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_14 XI11_7/net21_1_ xsel_12_ XI11_7/XI0/XI0_12/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_13 XI11_7/net21_2_ xsel_12_ XI11_7/XI0/XI0_12/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_12 XI11_7/net21_3_ xsel_12_ XI11_7/XI0/XI0_12/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_11 XI11_7/net21_4_ xsel_12_ XI11_7/XI0/XI0_12/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_10 XI11_7/net21_5_ xsel_12_ XI11_7/XI0/XI0_12/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_9 XI11_7/net21_6_ xsel_12_ XI11_7/XI0/XI0_12/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_8 XI11_7/net21_7_ xsel_12_ XI11_7/XI0/XI0_12/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_7 XI11_7/net21_8_ xsel_12_ XI11_7/XI0/XI0_12/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_6 XI11_7/net21_9_ xsel_12_ XI11_7/XI0/XI0_12/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_5 XI11_7/net21_10_ xsel_12_ XI11_7/XI0/XI0_12/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_4 XI11_7/net21_11_ xsel_12_ XI11_7/XI0/XI0_12/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_3 XI11_7/net21_12_ xsel_12_ XI11_7/XI0/XI0_12/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_2 XI11_7/net21_13_ xsel_12_ XI11_7/XI0/XI0_12/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_1 XI11_7/net21_14_ xsel_12_ XI11_7/XI0/XI0_12/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_0 XI11_7/net21_15_ xsel_12_ XI11_7/XI0/XI0_12/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_15 XI11_7/XI0/XI0_12/d__15_ xsel_12_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_14 XI11_7/XI0/XI0_12/d__14_ xsel_12_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_13 XI11_7/XI0/XI0_12/d__13_ xsel_12_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_12 XI11_7/XI0/XI0_12/d__12_ xsel_12_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_11 XI11_7/XI0/XI0_12/d__11_ xsel_12_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_10 XI11_7/XI0/XI0_12/d__10_ xsel_12_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_9 XI11_7/XI0/XI0_12/d__9_ xsel_12_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_8 XI11_7/XI0/XI0_12/d__8_ xsel_12_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_7 XI11_7/XI0/XI0_12/d__7_ xsel_12_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_6 XI11_7/XI0/XI0_12/d__6_ xsel_12_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_5 XI11_7/XI0/XI0_12/d__5_ xsel_12_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_4 XI11_7/XI0/XI0_12/d__4_ xsel_12_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_3 XI11_7/XI0/XI0_12/d__3_ xsel_12_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_2 XI11_7/XI0/XI0_12/d__2_ xsel_12_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_1 XI11_7/XI0/XI0_12/d__1_ xsel_12_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_0 XI11_7/XI0/XI0_12/d__0_ xsel_12_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_15 XI11_7/net21_0_ xsel_11_ XI11_7/XI0/XI0_11/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_14 XI11_7/net21_1_ xsel_11_ XI11_7/XI0/XI0_11/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_13 XI11_7/net21_2_ xsel_11_ XI11_7/XI0/XI0_11/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_12 XI11_7/net21_3_ xsel_11_ XI11_7/XI0/XI0_11/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_11 XI11_7/net21_4_ xsel_11_ XI11_7/XI0/XI0_11/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_10 XI11_7/net21_5_ xsel_11_ XI11_7/XI0/XI0_11/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_9 XI11_7/net21_6_ xsel_11_ XI11_7/XI0/XI0_11/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_8 XI11_7/net21_7_ xsel_11_ XI11_7/XI0/XI0_11/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_7 XI11_7/net21_8_ xsel_11_ XI11_7/XI0/XI0_11/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_6 XI11_7/net21_9_ xsel_11_ XI11_7/XI0/XI0_11/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_5 XI11_7/net21_10_ xsel_11_ XI11_7/XI0/XI0_11/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_4 XI11_7/net21_11_ xsel_11_ XI11_7/XI0/XI0_11/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_3 XI11_7/net21_12_ xsel_11_ XI11_7/XI0/XI0_11/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_2 XI11_7/net21_13_ xsel_11_ XI11_7/XI0/XI0_11/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_1 XI11_7/net21_14_ xsel_11_ XI11_7/XI0/XI0_11/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_0 XI11_7/net21_15_ xsel_11_ XI11_7/XI0/XI0_11/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_15 XI11_7/XI0/XI0_11/d__15_ xsel_11_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_14 XI11_7/XI0/XI0_11/d__14_ xsel_11_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_13 XI11_7/XI0/XI0_11/d__13_ xsel_11_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_12 XI11_7/XI0/XI0_11/d__12_ xsel_11_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_11 XI11_7/XI0/XI0_11/d__11_ xsel_11_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_10 XI11_7/XI0/XI0_11/d__10_ xsel_11_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_9 XI11_7/XI0/XI0_11/d__9_ xsel_11_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_8 XI11_7/XI0/XI0_11/d__8_ xsel_11_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_7 XI11_7/XI0/XI0_11/d__7_ xsel_11_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_6 XI11_7/XI0/XI0_11/d__6_ xsel_11_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_5 XI11_7/XI0/XI0_11/d__5_ xsel_11_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_4 XI11_7/XI0/XI0_11/d__4_ xsel_11_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_3 XI11_7/XI0/XI0_11/d__3_ xsel_11_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_2 XI11_7/XI0/XI0_11/d__2_ xsel_11_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_1 XI11_7/XI0/XI0_11/d__1_ xsel_11_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_0 XI11_7/XI0/XI0_11/d__0_ xsel_11_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_15 XI11_7/net21_0_ xsel_10_ XI11_7/XI0/XI0_10/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_14 XI11_7/net21_1_ xsel_10_ XI11_7/XI0/XI0_10/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_13 XI11_7/net21_2_ xsel_10_ XI11_7/XI0/XI0_10/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_12 XI11_7/net21_3_ xsel_10_ XI11_7/XI0/XI0_10/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_11 XI11_7/net21_4_ xsel_10_ XI11_7/XI0/XI0_10/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_10 XI11_7/net21_5_ xsel_10_ XI11_7/XI0/XI0_10/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_9 XI11_7/net21_6_ xsel_10_ XI11_7/XI0/XI0_10/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_8 XI11_7/net21_7_ xsel_10_ XI11_7/XI0/XI0_10/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_7 XI11_7/net21_8_ xsel_10_ XI11_7/XI0/XI0_10/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_6 XI11_7/net21_9_ xsel_10_ XI11_7/XI0/XI0_10/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_5 XI11_7/net21_10_ xsel_10_ XI11_7/XI0/XI0_10/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_4 XI11_7/net21_11_ xsel_10_ XI11_7/XI0/XI0_10/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_3 XI11_7/net21_12_ xsel_10_ XI11_7/XI0/XI0_10/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_2 XI11_7/net21_13_ xsel_10_ XI11_7/XI0/XI0_10/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_1 XI11_7/net21_14_ xsel_10_ XI11_7/XI0/XI0_10/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_0 XI11_7/net21_15_ xsel_10_ XI11_7/XI0/XI0_10/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_15 XI11_7/XI0/XI0_10/d__15_ xsel_10_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_14 XI11_7/XI0/XI0_10/d__14_ xsel_10_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_13 XI11_7/XI0/XI0_10/d__13_ xsel_10_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_12 XI11_7/XI0/XI0_10/d__12_ xsel_10_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_11 XI11_7/XI0/XI0_10/d__11_ xsel_10_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_10 XI11_7/XI0/XI0_10/d__10_ xsel_10_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_9 XI11_7/XI0/XI0_10/d__9_ xsel_10_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_8 XI11_7/XI0/XI0_10/d__8_ xsel_10_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_7 XI11_7/XI0/XI0_10/d__7_ xsel_10_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_6 XI11_7/XI0/XI0_10/d__6_ xsel_10_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_5 XI11_7/XI0/XI0_10/d__5_ xsel_10_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_4 XI11_7/XI0/XI0_10/d__4_ xsel_10_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_3 XI11_7/XI0/XI0_10/d__3_ xsel_10_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_2 XI11_7/XI0/XI0_10/d__2_ xsel_10_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_1 XI11_7/XI0/XI0_10/d__1_ xsel_10_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_0 XI11_7/XI0/XI0_10/d__0_ xsel_10_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_15 XI11_7/net21_0_ xsel_9_ XI11_7/XI0/XI0_9/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_14 XI11_7/net21_1_ xsel_9_ XI11_7/XI0/XI0_9/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_13 XI11_7/net21_2_ xsel_9_ XI11_7/XI0/XI0_9/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_12 XI11_7/net21_3_ xsel_9_ XI11_7/XI0/XI0_9/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_11 XI11_7/net21_4_ xsel_9_ XI11_7/XI0/XI0_9/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_10 XI11_7/net21_5_ xsel_9_ XI11_7/XI0/XI0_9/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_9 XI11_7/net21_6_ xsel_9_ XI11_7/XI0/XI0_9/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_8 XI11_7/net21_7_ xsel_9_ XI11_7/XI0/XI0_9/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_7 XI11_7/net21_8_ xsel_9_ XI11_7/XI0/XI0_9/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_6 XI11_7/net21_9_ xsel_9_ XI11_7/XI0/XI0_9/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_5 XI11_7/net21_10_ xsel_9_ XI11_7/XI0/XI0_9/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_4 XI11_7/net21_11_ xsel_9_ XI11_7/XI0/XI0_9/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_3 XI11_7/net21_12_ xsel_9_ XI11_7/XI0/XI0_9/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_2 XI11_7/net21_13_ xsel_9_ XI11_7/XI0/XI0_9/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_1 XI11_7/net21_14_ xsel_9_ XI11_7/XI0/XI0_9/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_0 XI11_7/net21_15_ xsel_9_ XI11_7/XI0/XI0_9/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_15 XI11_7/XI0/XI0_9/d__15_ xsel_9_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_14 XI11_7/XI0/XI0_9/d__14_ xsel_9_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_13 XI11_7/XI0/XI0_9/d__13_ xsel_9_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_12 XI11_7/XI0/XI0_9/d__12_ xsel_9_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_11 XI11_7/XI0/XI0_9/d__11_ xsel_9_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_10 XI11_7/XI0/XI0_9/d__10_ xsel_9_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_9 XI11_7/XI0/XI0_9/d__9_ xsel_9_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_8 XI11_7/XI0/XI0_9/d__8_ xsel_9_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_7 XI11_7/XI0/XI0_9/d__7_ xsel_9_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_6 XI11_7/XI0/XI0_9/d__6_ xsel_9_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_5 XI11_7/XI0/XI0_9/d__5_ xsel_9_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_4 XI11_7/XI0/XI0_9/d__4_ xsel_9_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_3 XI11_7/XI0/XI0_9/d__3_ xsel_9_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_2 XI11_7/XI0/XI0_9/d__2_ xsel_9_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_1 XI11_7/XI0/XI0_9/d__1_ xsel_9_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_0 XI11_7/XI0/XI0_9/d__0_ xsel_9_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_15 XI11_7/net21_0_ xsel_8_ XI11_7/XI0/XI0_8/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_14 XI11_7/net21_1_ xsel_8_ XI11_7/XI0/XI0_8/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_13 XI11_7/net21_2_ xsel_8_ XI11_7/XI0/XI0_8/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_12 XI11_7/net21_3_ xsel_8_ XI11_7/XI0/XI0_8/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_11 XI11_7/net21_4_ xsel_8_ XI11_7/XI0/XI0_8/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_10 XI11_7/net21_5_ xsel_8_ XI11_7/XI0/XI0_8/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_9 XI11_7/net21_6_ xsel_8_ XI11_7/XI0/XI0_8/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_8 XI11_7/net21_7_ xsel_8_ XI11_7/XI0/XI0_8/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_7 XI11_7/net21_8_ xsel_8_ XI11_7/XI0/XI0_8/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_6 XI11_7/net21_9_ xsel_8_ XI11_7/XI0/XI0_8/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_5 XI11_7/net21_10_ xsel_8_ XI11_7/XI0/XI0_8/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_4 XI11_7/net21_11_ xsel_8_ XI11_7/XI0/XI0_8/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_3 XI11_7/net21_12_ xsel_8_ XI11_7/XI0/XI0_8/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_2 XI11_7/net21_13_ xsel_8_ XI11_7/XI0/XI0_8/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_1 XI11_7/net21_14_ xsel_8_ XI11_7/XI0/XI0_8/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_0 XI11_7/net21_15_ xsel_8_ XI11_7/XI0/XI0_8/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_15 XI11_7/XI0/XI0_8/d__15_ xsel_8_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_14 XI11_7/XI0/XI0_8/d__14_ xsel_8_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_13 XI11_7/XI0/XI0_8/d__13_ xsel_8_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_12 XI11_7/XI0/XI0_8/d__12_ xsel_8_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_11 XI11_7/XI0/XI0_8/d__11_ xsel_8_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_10 XI11_7/XI0/XI0_8/d__10_ xsel_8_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_9 XI11_7/XI0/XI0_8/d__9_ xsel_8_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_8 XI11_7/XI0/XI0_8/d__8_ xsel_8_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_7 XI11_7/XI0/XI0_8/d__7_ xsel_8_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_6 XI11_7/XI0/XI0_8/d__6_ xsel_8_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_5 XI11_7/XI0/XI0_8/d__5_ xsel_8_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_4 XI11_7/XI0/XI0_8/d__4_ xsel_8_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_3 XI11_7/XI0/XI0_8/d__3_ xsel_8_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_2 XI11_7/XI0/XI0_8/d__2_ xsel_8_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_1 XI11_7/XI0/XI0_8/d__1_ xsel_8_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_0 XI11_7/XI0/XI0_8/d__0_ xsel_8_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_15 XI11_7/net21_0_ xsel_7_ XI11_7/XI0/XI0_7/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_14 XI11_7/net21_1_ xsel_7_ XI11_7/XI0/XI0_7/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_13 XI11_7/net21_2_ xsel_7_ XI11_7/XI0/XI0_7/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_12 XI11_7/net21_3_ xsel_7_ XI11_7/XI0/XI0_7/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_11 XI11_7/net21_4_ xsel_7_ XI11_7/XI0/XI0_7/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_10 XI11_7/net21_5_ xsel_7_ XI11_7/XI0/XI0_7/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_9 XI11_7/net21_6_ xsel_7_ XI11_7/XI0/XI0_7/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_8 XI11_7/net21_7_ xsel_7_ XI11_7/XI0/XI0_7/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_7 XI11_7/net21_8_ xsel_7_ XI11_7/XI0/XI0_7/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_6 XI11_7/net21_9_ xsel_7_ XI11_7/XI0/XI0_7/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_5 XI11_7/net21_10_ xsel_7_ XI11_7/XI0/XI0_7/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_4 XI11_7/net21_11_ xsel_7_ XI11_7/XI0/XI0_7/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_3 XI11_7/net21_12_ xsel_7_ XI11_7/XI0/XI0_7/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_2 XI11_7/net21_13_ xsel_7_ XI11_7/XI0/XI0_7/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_1 XI11_7/net21_14_ xsel_7_ XI11_7/XI0/XI0_7/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_0 XI11_7/net21_15_ xsel_7_ XI11_7/XI0/XI0_7/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_15 XI11_7/XI0/XI0_7/d__15_ xsel_7_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_14 XI11_7/XI0/XI0_7/d__14_ xsel_7_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_13 XI11_7/XI0/XI0_7/d__13_ xsel_7_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_12 XI11_7/XI0/XI0_7/d__12_ xsel_7_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_11 XI11_7/XI0/XI0_7/d__11_ xsel_7_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_10 XI11_7/XI0/XI0_7/d__10_ xsel_7_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_9 XI11_7/XI0/XI0_7/d__9_ xsel_7_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_8 XI11_7/XI0/XI0_7/d__8_ xsel_7_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_7 XI11_7/XI0/XI0_7/d__7_ xsel_7_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_6 XI11_7/XI0/XI0_7/d__6_ xsel_7_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_5 XI11_7/XI0/XI0_7/d__5_ xsel_7_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_4 XI11_7/XI0/XI0_7/d__4_ xsel_7_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_3 XI11_7/XI0/XI0_7/d__3_ xsel_7_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_2 XI11_7/XI0/XI0_7/d__2_ xsel_7_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_1 XI11_7/XI0/XI0_7/d__1_ xsel_7_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_0 XI11_7/XI0/XI0_7/d__0_ xsel_7_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_15 XI11_7/net21_0_ xsel_6_ XI11_7/XI0/XI0_6/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_14 XI11_7/net21_1_ xsel_6_ XI11_7/XI0/XI0_6/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_13 XI11_7/net21_2_ xsel_6_ XI11_7/XI0/XI0_6/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_12 XI11_7/net21_3_ xsel_6_ XI11_7/XI0/XI0_6/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_11 XI11_7/net21_4_ xsel_6_ XI11_7/XI0/XI0_6/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_10 XI11_7/net21_5_ xsel_6_ XI11_7/XI0/XI0_6/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_9 XI11_7/net21_6_ xsel_6_ XI11_7/XI0/XI0_6/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_8 XI11_7/net21_7_ xsel_6_ XI11_7/XI0/XI0_6/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_7 XI11_7/net21_8_ xsel_6_ XI11_7/XI0/XI0_6/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_6 XI11_7/net21_9_ xsel_6_ XI11_7/XI0/XI0_6/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_5 XI11_7/net21_10_ xsel_6_ XI11_7/XI0/XI0_6/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_4 XI11_7/net21_11_ xsel_6_ XI11_7/XI0/XI0_6/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_3 XI11_7/net21_12_ xsel_6_ XI11_7/XI0/XI0_6/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_2 XI11_7/net21_13_ xsel_6_ XI11_7/XI0/XI0_6/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_1 XI11_7/net21_14_ xsel_6_ XI11_7/XI0/XI0_6/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_0 XI11_7/net21_15_ xsel_6_ XI11_7/XI0/XI0_6/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_15 XI11_7/XI0/XI0_6/d__15_ xsel_6_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_14 XI11_7/XI0/XI0_6/d__14_ xsel_6_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_13 XI11_7/XI0/XI0_6/d__13_ xsel_6_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_12 XI11_7/XI0/XI0_6/d__12_ xsel_6_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_11 XI11_7/XI0/XI0_6/d__11_ xsel_6_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_10 XI11_7/XI0/XI0_6/d__10_ xsel_6_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_9 XI11_7/XI0/XI0_6/d__9_ xsel_6_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_8 XI11_7/XI0/XI0_6/d__8_ xsel_6_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_7 XI11_7/XI0/XI0_6/d__7_ xsel_6_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_6 XI11_7/XI0/XI0_6/d__6_ xsel_6_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_5 XI11_7/XI0/XI0_6/d__5_ xsel_6_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_4 XI11_7/XI0/XI0_6/d__4_ xsel_6_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_3 XI11_7/XI0/XI0_6/d__3_ xsel_6_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_2 XI11_7/XI0/XI0_6/d__2_ xsel_6_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_1 XI11_7/XI0/XI0_6/d__1_ xsel_6_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_0 XI11_7/XI0/XI0_6/d__0_ xsel_6_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_15 XI11_7/net21_0_ xsel_5_ XI11_7/XI0/XI0_5/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_14 XI11_7/net21_1_ xsel_5_ XI11_7/XI0/XI0_5/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_13 XI11_7/net21_2_ xsel_5_ XI11_7/XI0/XI0_5/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_12 XI11_7/net21_3_ xsel_5_ XI11_7/XI0/XI0_5/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_11 XI11_7/net21_4_ xsel_5_ XI11_7/XI0/XI0_5/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_10 XI11_7/net21_5_ xsel_5_ XI11_7/XI0/XI0_5/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_9 XI11_7/net21_6_ xsel_5_ XI11_7/XI0/XI0_5/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_8 XI11_7/net21_7_ xsel_5_ XI11_7/XI0/XI0_5/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_7 XI11_7/net21_8_ xsel_5_ XI11_7/XI0/XI0_5/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_6 XI11_7/net21_9_ xsel_5_ XI11_7/XI0/XI0_5/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_5 XI11_7/net21_10_ xsel_5_ XI11_7/XI0/XI0_5/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_4 XI11_7/net21_11_ xsel_5_ XI11_7/XI0/XI0_5/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_3 XI11_7/net21_12_ xsel_5_ XI11_7/XI0/XI0_5/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_2 XI11_7/net21_13_ xsel_5_ XI11_7/XI0/XI0_5/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_1 XI11_7/net21_14_ xsel_5_ XI11_7/XI0/XI0_5/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_0 XI11_7/net21_15_ xsel_5_ XI11_7/XI0/XI0_5/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_15 XI11_7/XI0/XI0_5/d__15_ xsel_5_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_14 XI11_7/XI0/XI0_5/d__14_ xsel_5_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_13 XI11_7/XI0/XI0_5/d__13_ xsel_5_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_12 XI11_7/XI0/XI0_5/d__12_ xsel_5_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_11 XI11_7/XI0/XI0_5/d__11_ xsel_5_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_10 XI11_7/XI0/XI0_5/d__10_ xsel_5_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_9 XI11_7/XI0/XI0_5/d__9_ xsel_5_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_8 XI11_7/XI0/XI0_5/d__8_ xsel_5_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_7 XI11_7/XI0/XI0_5/d__7_ xsel_5_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_6 XI11_7/XI0/XI0_5/d__6_ xsel_5_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_5 XI11_7/XI0/XI0_5/d__5_ xsel_5_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_4 XI11_7/XI0/XI0_5/d__4_ xsel_5_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_3 XI11_7/XI0/XI0_5/d__3_ xsel_5_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_2 XI11_7/XI0/XI0_5/d__2_ xsel_5_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_1 XI11_7/XI0/XI0_5/d__1_ xsel_5_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_0 XI11_7/XI0/XI0_5/d__0_ xsel_5_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_15 XI11_7/net21_0_ xsel_4_ XI11_7/XI0/XI0_4/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_14 XI11_7/net21_1_ xsel_4_ XI11_7/XI0/XI0_4/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_13 XI11_7/net21_2_ xsel_4_ XI11_7/XI0/XI0_4/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_12 XI11_7/net21_3_ xsel_4_ XI11_7/XI0/XI0_4/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_11 XI11_7/net21_4_ xsel_4_ XI11_7/XI0/XI0_4/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_10 XI11_7/net21_5_ xsel_4_ XI11_7/XI0/XI0_4/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_9 XI11_7/net21_6_ xsel_4_ XI11_7/XI0/XI0_4/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_8 XI11_7/net21_7_ xsel_4_ XI11_7/XI0/XI0_4/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_7 XI11_7/net21_8_ xsel_4_ XI11_7/XI0/XI0_4/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_6 XI11_7/net21_9_ xsel_4_ XI11_7/XI0/XI0_4/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_5 XI11_7/net21_10_ xsel_4_ XI11_7/XI0/XI0_4/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_4 XI11_7/net21_11_ xsel_4_ XI11_7/XI0/XI0_4/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_3 XI11_7/net21_12_ xsel_4_ XI11_7/XI0/XI0_4/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_2 XI11_7/net21_13_ xsel_4_ XI11_7/XI0/XI0_4/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_1 XI11_7/net21_14_ xsel_4_ XI11_7/XI0/XI0_4/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_0 XI11_7/net21_15_ xsel_4_ XI11_7/XI0/XI0_4/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_15 XI11_7/XI0/XI0_4/d__15_ xsel_4_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_14 XI11_7/XI0/XI0_4/d__14_ xsel_4_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_13 XI11_7/XI0/XI0_4/d__13_ xsel_4_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_12 XI11_7/XI0/XI0_4/d__12_ xsel_4_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_11 XI11_7/XI0/XI0_4/d__11_ xsel_4_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_10 XI11_7/XI0/XI0_4/d__10_ xsel_4_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_9 XI11_7/XI0/XI0_4/d__9_ xsel_4_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_8 XI11_7/XI0/XI0_4/d__8_ xsel_4_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_7 XI11_7/XI0/XI0_4/d__7_ xsel_4_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_6 XI11_7/XI0/XI0_4/d__6_ xsel_4_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_5 XI11_7/XI0/XI0_4/d__5_ xsel_4_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_4 XI11_7/XI0/XI0_4/d__4_ xsel_4_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_3 XI11_7/XI0/XI0_4/d__3_ xsel_4_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_2 XI11_7/XI0/XI0_4/d__2_ xsel_4_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_1 XI11_7/XI0/XI0_4/d__1_ xsel_4_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_0 XI11_7/XI0/XI0_4/d__0_ xsel_4_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_15 XI11_7/net21_0_ xsel_3_ XI11_7/XI0/XI0_3/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_14 XI11_7/net21_1_ xsel_3_ XI11_7/XI0/XI0_3/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_13 XI11_7/net21_2_ xsel_3_ XI11_7/XI0/XI0_3/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_12 XI11_7/net21_3_ xsel_3_ XI11_7/XI0/XI0_3/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_11 XI11_7/net21_4_ xsel_3_ XI11_7/XI0/XI0_3/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_10 XI11_7/net21_5_ xsel_3_ XI11_7/XI0/XI0_3/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_9 XI11_7/net21_6_ xsel_3_ XI11_7/XI0/XI0_3/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_8 XI11_7/net21_7_ xsel_3_ XI11_7/XI0/XI0_3/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_7 XI11_7/net21_8_ xsel_3_ XI11_7/XI0/XI0_3/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_6 XI11_7/net21_9_ xsel_3_ XI11_7/XI0/XI0_3/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_5 XI11_7/net21_10_ xsel_3_ XI11_7/XI0/XI0_3/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_4 XI11_7/net21_11_ xsel_3_ XI11_7/XI0/XI0_3/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_3 XI11_7/net21_12_ xsel_3_ XI11_7/XI0/XI0_3/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_2 XI11_7/net21_13_ xsel_3_ XI11_7/XI0/XI0_3/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_1 XI11_7/net21_14_ xsel_3_ XI11_7/XI0/XI0_3/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_0 XI11_7/net21_15_ xsel_3_ XI11_7/XI0/XI0_3/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_15 XI11_7/XI0/XI0_3/d__15_ xsel_3_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_14 XI11_7/XI0/XI0_3/d__14_ xsel_3_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_13 XI11_7/XI0/XI0_3/d__13_ xsel_3_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_12 XI11_7/XI0/XI0_3/d__12_ xsel_3_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_11 XI11_7/XI0/XI0_3/d__11_ xsel_3_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_10 XI11_7/XI0/XI0_3/d__10_ xsel_3_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_9 XI11_7/XI0/XI0_3/d__9_ xsel_3_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_8 XI11_7/XI0/XI0_3/d__8_ xsel_3_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_7 XI11_7/XI0/XI0_3/d__7_ xsel_3_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_6 XI11_7/XI0/XI0_3/d__6_ xsel_3_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_5 XI11_7/XI0/XI0_3/d__5_ xsel_3_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_4 XI11_7/XI0/XI0_3/d__4_ xsel_3_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_3 XI11_7/XI0/XI0_3/d__3_ xsel_3_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_2 XI11_7/XI0/XI0_3/d__2_ xsel_3_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_1 XI11_7/XI0/XI0_3/d__1_ xsel_3_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_0 XI11_7/XI0/XI0_3/d__0_ xsel_3_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_15 XI11_7/net21_0_ xsel_2_ XI11_7/XI0/XI0_2/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_14 XI11_7/net21_1_ xsel_2_ XI11_7/XI0/XI0_2/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_13 XI11_7/net21_2_ xsel_2_ XI11_7/XI0/XI0_2/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_12 XI11_7/net21_3_ xsel_2_ XI11_7/XI0/XI0_2/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_11 XI11_7/net21_4_ xsel_2_ XI11_7/XI0/XI0_2/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_10 XI11_7/net21_5_ xsel_2_ XI11_7/XI0/XI0_2/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_9 XI11_7/net21_6_ xsel_2_ XI11_7/XI0/XI0_2/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_8 XI11_7/net21_7_ xsel_2_ XI11_7/XI0/XI0_2/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_7 XI11_7/net21_8_ xsel_2_ XI11_7/XI0/XI0_2/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_6 XI11_7/net21_9_ xsel_2_ XI11_7/XI0/XI0_2/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_5 XI11_7/net21_10_ xsel_2_ XI11_7/XI0/XI0_2/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_4 XI11_7/net21_11_ xsel_2_ XI11_7/XI0/XI0_2/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_3 XI11_7/net21_12_ xsel_2_ XI11_7/XI0/XI0_2/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_2 XI11_7/net21_13_ xsel_2_ XI11_7/XI0/XI0_2/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_1 XI11_7/net21_14_ xsel_2_ XI11_7/XI0/XI0_2/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_0 XI11_7/net21_15_ xsel_2_ XI11_7/XI0/XI0_2/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_15 XI11_7/XI0/XI0_2/d__15_ xsel_2_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_14 XI11_7/XI0/XI0_2/d__14_ xsel_2_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_13 XI11_7/XI0/XI0_2/d__13_ xsel_2_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_12 XI11_7/XI0/XI0_2/d__12_ xsel_2_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_11 XI11_7/XI0/XI0_2/d__11_ xsel_2_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_10 XI11_7/XI0/XI0_2/d__10_ xsel_2_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_9 XI11_7/XI0/XI0_2/d__9_ xsel_2_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_8 XI11_7/XI0/XI0_2/d__8_ xsel_2_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_7 XI11_7/XI0/XI0_2/d__7_ xsel_2_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_6 XI11_7/XI0/XI0_2/d__6_ xsel_2_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_5 XI11_7/XI0/XI0_2/d__5_ xsel_2_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_4 XI11_7/XI0/XI0_2/d__4_ xsel_2_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_3 XI11_7/XI0/XI0_2/d__3_ xsel_2_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_2 XI11_7/XI0/XI0_2/d__2_ xsel_2_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_1 XI11_7/XI0/XI0_2/d__1_ xsel_2_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_0 XI11_7/XI0/XI0_2/d__0_ xsel_2_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_15 XI11_7/net21_0_ xsel_1_ XI11_7/XI0/XI0_1/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_14 XI11_7/net21_1_ xsel_1_ XI11_7/XI0/XI0_1/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_13 XI11_7/net21_2_ xsel_1_ XI11_7/XI0/XI0_1/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_12 XI11_7/net21_3_ xsel_1_ XI11_7/XI0/XI0_1/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_11 XI11_7/net21_4_ xsel_1_ XI11_7/XI0/XI0_1/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_10 XI11_7/net21_5_ xsel_1_ XI11_7/XI0/XI0_1/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_9 XI11_7/net21_6_ xsel_1_ XI11_7/XI0/XI0_1/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_8 XI11_7/net21_7_ xsel_1_ XI11_7/XI0/XI0_1/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_7 XI11_7/net21_8_ xsel_1_ XI11_7/XI0/XI0_1/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_6 XI11_7/net21_9_ xsel_1_ XI11_7/XI0/XI0_1/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_5 XI11_7/net21_10_ xsel_1_ XI11_7/XI0/XI0_1/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_4 XI11_7/net21_11_ xsel_1_ XI11_7/XI0/XI0_1/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_3 XI11_7/net21_12_ xsel_1_ XI11_7/XI0/XI0_1/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_2 XI11_7/net21_13_ xsel_1_ XI11_7/XI0/XI0_1/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_1 XI11_7/net21_14_ xsel_1_ XI11_7/XI0/XI0_1/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_0 XI11_7/net21_15_ xsel_1_ XI11_7/XI0/XI0_1/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_15 XI11_7/XI0/XI0_1/d__15_ xsel_1_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_14 XI11_7/XI0/XI0_1/d__14_ xsel_1_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_13 XI11_7/XI0/XI0_1/d__13_ xsel_1_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_12 XI11_7/XI0/XI0_1/d__12_ xsel_1_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_11 XI11_7/XI0/XI0_1/d__11_ xsel_1_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_10 XI11_7/XI0/XI0_1/d__10_ xsel_1_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_9 XI11_7/XI0/XI0_1/d__9_ xsel_1_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_8 XI11_7/XI0/XI0_1/d__8_ xsel_1_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_7 XI11_7/XI0/XI0_1/d__7_ xsel_1_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_6 XI11_7/XI0/XI0_1/d__6_ xsel_1_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_5 XI11_7/XI0/XI0_1/d__5_ xsel_1_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_4 XI11_7/XI0/XI0_1/d__4_ xsel_1_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_3 XI11_7/XI0/XI0_1/d__3_ xsel_1_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_2 XI11_7/XI0/XI0_1/d__2_ xsel_1_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_1 XI11_7/XI0/XI0_1/d__1_ xsel_1_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_0 XI11_7/XI0/XI0_1/d__0_ xsel_1_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_15 XI11_7/net21_0_ xsel_0_ XI11_7/XI0/XI0_0/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_14 XI11_7/net21_1_ xsel_0_ XI11_7/XI0/XI0_0/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_13 XI11_7/net21_2_ xsel_0_ XI11_7/XI0/XI0_0/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_12 XI11_7/net21_3_ xsel_0_ XI11_7/XI0/XI0_0/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_11 XI11_7/net21_4_ xsel_0_ XI11_7/XI0/XI0_0/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_10 XI11_7/net21_5_ xsel_0_ XI11_7/XI0/XI0_0/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_9 XI11_7/net21_6_ xsel_0_ XI11_7/XI0/XI0_0/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_8 XI11_7/net21_7_ xsel_0_ XI11_7/XI0/XI0_0/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_7 XI11_7/net21_8_ xsel_0_ XI11_7/XI0/XI0_0/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_6 XI11_7/net21_9_ xsel_0_ XI11_7/XI0/XI0_0/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_5 XI11_7/net21_10_ xsel_0_ XI11_7/XI0/XI0_0/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_4 XI11_7/net21_11_ xsel_0_ XI11_7/XI0/XI0_0/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_3 XI11_7/net21_12_ xsel_0_ XI11_7/XI0/XI0_0/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_2 XI11_7/net21_13_ xsel_0_ XI11_7/XI0/XI0_0/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_1 XI11_7/net21_14_ xsel_0_ XI11_7/XI0/XI0_0/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_0 XI11_7/net21_15_ xsel_0_ XI11_7/XI0/XI0_0/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_15 XI11_7/XI0/XI0_0/d__15_ xsel_0_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_14 XI11_7/XI0/XI0_0/d__14_ xsel_0_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_13 XI11_7/XI0/XI0_0/d__13_ xsel_0_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_12 XI11_7/XI0/XI0_0/d__12_ xsel_0_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_11 XI11_7/XI0/XI0_0/d__11_ xsel_0_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_10 XI11_7/XI0/XI0_0/d__10_ xsel_0_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_9 XI11_7/XI0/XI0_0/d__9_ xsel_0_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_8 XI11_7/XI0/XI0_0/d__8_ xsel_0_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_7 XI11_7/XI0/XI0_0/d__7_ xsel_0_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_6 XI11_7/XI0/XI0_0/d__6_ xsel_0_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_5 XI11_7/XI0/XI0_0/d__5_ xsel_0_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_4 XI11_7/XI0/XI0_0/d__4_ xsel_0_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_3 XI11_7/XI0/XI0_0/d__3_ xsel_0_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_2 XI11_7/XI0/XI0_0/d__2_ xsel_0_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_1 XI11_7/XI0/XI0_0/d__1_ xsel_0_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_0 XI11_7/XI0/XI0_0/d__0_ xsel_0_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI2/MN0_15 XI11_6/net21_0_ ysel_15_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_14 XI11_6/net21_1_ ysel_14_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_13 XI11_6/net21_2_ ysel_13_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_12 XI11_6/net21_3_ ysel_12_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_11 XI11_6/net21_4_ ysel_11_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_10 XI11_6/net21_5_ ysel_10_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_9 XI11_6/net21_6_ ysel_9_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_8 XI11_6/net21_7_ ysel_8_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_7 XI11_6/net21_8_ ysel_7_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_6 XI11_6/net21_9_ ysel_6_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_5 XI11_6/net21_10_ ysel_5_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_4 XI11_6/net21_11_ ysel_4_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_3 XI11_6/net21_12_ ysel_3_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_2 XI11_6/net21_13_ ysel_2_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_1 XI11_6/net21_14_ ysel_1_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_0 XI11_6/net21_15_ ysel_0_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_15 XI11_6/net20_0_ ysel_15_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_14 XI11_6/net20_1_ ysel_14_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_13 XI11_6/net20_2_ ysel_13_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_12 XI11_6/net20_3_ ysel_12_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_11 XI11_6/net20_4_ ysel_11_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_10 XI11_6/net20_5_ ysel_10_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_9 XI11_6/net20_6_ ysel_9_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_8 XI11_6/net20_7_ ysel_8_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_7 XI11_6/net20_8_ ysel_7_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_6 XI11_6/net20_9_ ysel_6_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_5 XI11_6/net20_10_ ysel_5_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_4 XI11_6/net20_11_ ysel_4_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_3 XI11_6/net20_12_ ysel_3_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_2 XI11_6/net20_13_ ysel_2_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_1 XI11_6/net20_14_ ysel_1_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_0 XI11_6/net20_15_ ysel_0_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI4/MN8 vdd XI11_6/XI4/net8 XI11_6/net12 vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_6/XI4/MP0 XI11_6/net9 XI11_6/XI4/net23 vdd vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_6/XI4/MP4 XI11_6/net12 XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI4/MP1 XI11_6/net9 XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI4/MP5 XI11_6/net12 XI11_6/preck XI11_6/net9 vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI4/MN7 vdd XI11_6/XI4/net090 DOUT_6_ vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_6/XI4/MP3 gnd XI11_6/XI4/net089 XI11_6/net12 gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_6/XI4/MN5 XI11_6/net9 XI11_6/XI4/net0103 gnd gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_6/XI4/MN4 XI11_6/XI4/data_out_ XI11_6/XI4/net32 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_6/XI4/MN0 XI11_6/XI4/data_out XI11_6/XI4/net52 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_6/XI4/MN9 gnd XI11_6/XI4/net0112 DOUT_6_ gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_6/XI1_15/MP2 XI11_6/net20_0_ XI11_6/preck XI11_6/net21_0_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_15/MP1 XI11_6/net20_0_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_15/MP0 XI11_6/net21_0_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_14/MP2 XI11_6/net20_1_ XI11_6/preck XI11_6/net21_1_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_14/MP1 XI11_6/net20_1_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_14/MP0 XI11_6/net21_1_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_13/MP2 XI11_6/net20_2_ XI11_6/preck XI11_6/net21_2_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_13/MP1 XI11_6/net20_2_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_13/MP0 XI11_6/net21_2_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_12/MP2 XI11_6/net20_3_ XI11_6/preck XI11_6/net21_3_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_12/MP1 XI11_6/net20_3_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_12/MP0 XI11_6/net21_3_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_11/MP2 XI11_6/net20_4_ XI11_6/preck XI11_6/net21_4_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_11/MP1 XI11_6/net20_4_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_11/MP0 XI11_6/net21_4_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_10/MP2 XI11_6/net20_5_ XI11_6/preck XI11_6/net21_5_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_10/MP1 XI11_6/net20_5_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_10/MP0 XI11_6/net21_5_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_9/MP2 XI11_6/net20_6_ XI11_6/preck XI11_6/net21_6_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_9/MP1 XI11_6/net20_6_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_9/MP0 XI11_6/net21_6_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_8/MP2 XI11_6/net20_7_ XI11_6/preck XI11_6/net21_7_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_8/MP1 XI11_6/net20_7_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_8/MP0 XI11_6/net21_7_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_7/MP2 XI11_6/net20_8_ XI11_6/preck XI11_6/net21_8_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_7/MP1 XI11_6/net20_8_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_7/MP0 XI11_6/net21_8_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_6/MP2 XI11_6/net20_9_ XI11_6/preck XI11_6/net21_9_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_6/MP1 XI11_6/net20_9_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_6/MP0 XI11_6/net21_9_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_5/MP2 XI11_6/net20_10_ XI11_6/preck XI11_6/net21_10_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_5/MP1 XI11_6/net20_10_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_5/MP0 XI11_6/net21_10_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_4/MP2 XI11_6/net20_11_ XI11_6/preck XI11_6/net21_11_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_4/MP1 XI11_6/net20_11_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_4/MP0 XI11_6/net21_11_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_3/MP2 XI11_6/net20_12_ XI11_6/preck XI11_6/net21_12_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_3/MP1 XI11_6/net20_12_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_3/MP0 XI11_6/net21_12_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_2/MP2 XI11_6/net20_13_ XI11_6/preck XI11_6/net21_13_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_2/MP1 XI11_6/net20_13_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_2/MP0 XI11_6/net21_13_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_1/MP2 XI11_6/net20_14_ XI11_6/preck XI11_6/net21_14_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_1/MP1 XI11_6/net20_14_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_1/MP0 XI11_6/net21_14_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_0/MP2 XI11_6/net20_15_ XI11_6/preck XI11_6/net21_15_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_0/MP1 XI11_6/net20_15_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_0/MP0 XI11_6/net21_15_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI0/MN0_15 gnd gnd XI11_6/net21_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_14 gnd gnd XI11_6/net21_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_13 gnd gnd XI11_6/net21_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_12 gnd gnd XI11_6/net21_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_11 gnd gnd XI11_6/net21_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_10 gnd gnd XI11_6/net21_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_9 gnd gnd XI11_6/net21_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_8 gnd gnd XI11_6/net21_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_7 gnd gnd XI11_6/net21_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_6 gnd gnd XI11_6/net21_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_5 gnd gnd XI11_6/net21_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_4 gnd gnd XI11_6/net21_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_3 gnd gnd XI11_6/net21_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_2 gnd gnd XI11_6/net21_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_1 gnd gnd XI11_6/net21_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_0 gnd gnd XI11_6/net21_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_15 gnd gnd XI11_6/net20_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_14 gnd gnd XI11_6/net20_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_13 gnd gnd XI11_6/net20_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_12 gnd gnd XI11_6/net20_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_11 gnd gnd XI11_6/net20_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_10 gnd gnd XI11_6/net20_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_9 gnd gnd XI11_6/net20_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_8 gnd gnd XI11_6/net20_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_7 gnd gnd XI11_6/net20_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_6 gnd gnd XI11_6/net20_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_5 gnd gnd XI11_6/net20_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_4 gnd gnd XI11_6/net20_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_3 gnd gnd XI11_6/net20_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_2 gnd gnd XI11_6/net20_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_1 gnd gnd XI11_6/net20_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_0 gnd gnd XI11_6/net20_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_15 XI11_6/net21_0_ xsel_63_ XI11_6/XI0/XI0_63/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_14 XI11_6/net21_1_ xsel_63_ XI11_6/XI0/XI0_63/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_13 XI11_6/net21_2_ xsel_63_ XI11_6/XI0/XI0_63/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_12 XI11_6/net21_3_ xsel_63_ XI11_6/XI0/XI0_63/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_11 XI11_6/net21_4_ xsel_63_ XI11_6/XI0/XI0_63/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_10 XI11_6/net21_5_ xsel_63_ XI11_6/XI0/XI0_63/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_9 XI11_6/net21_6_ xsel_63_ XI11_6/XI0/XI0_63/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_8 XI11_6/net21_7_ xsel_63_ XI11_6/XI0/XI0_63/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_7 XI11_6/net21_8_ xsel_63_ XI11_6/XI0/XI0_63/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_6 XI11_6/net21_9_ xsel_63_ XI11_6/XI0/XI0_63/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_5 XI11_6/net21_10_ xsel_63_ XI11_6/XI0/XI0_63/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_4 XI11_6/net21_11_ xsel_63_ XI11_6/XI0/XI0_63/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_3 XI11_6/net21_12_ xsel_63_ XI11_6/XI0/XI0_63/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_2 XI11_6/net21_13_ xsel_63_ XI11_6/XI0/XI0_63/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_1 XI11_6/net21_14_ xsel_63_ XI11_6/XI0/XI0_63/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_0 XI11_6/net21_15_ xsel_63_ XI11_6/XI0/XI0_63/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_15 XI11_6/XI0/XI0_63/d__15_ xsel_63_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_14 XI11_6/XI0/XI0_63/d__14_ xsel_63_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_13 XI11_6/XI0/XI0_63/d__13_ xsel_63_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_12 XI11_6/XI0/XI0_63/d__12_ xsel_63_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_11 XI11_6/XI0/XI0_63/d__11_ xsel_63_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_10 XI11_6/XI0/XI0_63/d__10_ xsel_63_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_9 XI11_6/XI0/XI0_63/d__9_ xsel_63_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_8 XI11_6/XI0/XI0_63/d__8_ xsel_63_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_7 XI11_6/XI0/XI0_63/d__7_ xsel_63_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_6 XI11_6/XI0/XI0_63/d__6_ xsel_63_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_5 XI11_6/XI0/XI0_63/d__5_ xsel_63_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_4 XI11_6/XI0/XI0_63/d__4_ xsel_63_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_3 XI11_6/XI0/XI0_63/d__3_ xsel_63_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_2 XI11_6/XI0/XI0_63/d__2_ xsel_63_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_1 XI11_6/XI0/XI0_63/d__1_ xsel_63_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_0 XI11_6/XI0/XI0_63/d__0_ xsel_63_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_15 XI11_6/net21_0_ xsel_62_ XI11_6/XI0/XI0_62/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_14 XI11_6/net21_1_ xsel_62_ XI11_6/XI0/XI0_62/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_13 XI11_6/net21_2_ xsel_62_ XI11_6/XI0/XI0_62/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_12 XI11_6/net21_3_ xsel_62_ XI11_6/XI0/XI0_62/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_11 XI11_6/net21_4_ xsel_62_ XI11_6/XI0/XI0_62/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_10 XI11_6/net21_5_ xsel_62_ XI11_6/XI0/XI0_62/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_9 XI11_6/net21_6_ xsel_62_ XI11_6/XI0/XI0_62/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_8 XI11_6/net21_7_ xsel_62_ XI11_6/XI0/XI0_62/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_7 XI11_6/net21_8_ xsel_62_ XI11_6/XI0/XI0_62/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_6 XI11_6/net21_9_ xsel_62_ XI11_6/XI0/XI0_62/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_5 XI11_6/net21_10_ xsel_62_ XI11_6/XI0/XI0_62/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_4 XI11_6/net21_11_ xsel_62_ XI11_6/XI0/XI0_62/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_3 XI11_6/net21_12_ xsel_62_ XI11_6/XI0/XI0_62/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_2 XI11_6/net21_13_ xsel_62_ XI11_6/XI0/XI0_62/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_1 XI11_6/net21_14_ xsel_62_ XI11_6/XI0/XI0_62/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_0 XI11_6/net21_15_ xsel_62_ XI11_6/XI0/XI0_62/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_15 XI11_6/XI0/XI0_62/d__15_ xsel_62_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_14 XI11_6/XI0/XI0_62/d__14_ xsel_62_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_13 XI11_6/XI0/XI0_62/d__13_ xsel_62_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_12 XI11_6/XI0/XI0_62/d__12_ xsel_62_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_11 XI11_6/XI0/XI0_62/d__11_ xsel_62_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_10 XI11_6/XI0/XI0_62/d__10_ xsel_62_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_9 XI11_6/XI0/XI0_62/d__9_ xsel_62_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_8 XI11_6/XI0/XI0_62/d__8_ xsel_62_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_7 XI11_6/XI0/XI0_62/d__7_ xsel_62_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_6 XI11_6/XI0/XI0_62/d__6_ xsel_62_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_5 XI11_6/XI0/XI0_62/d__5_ xsel_62_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_4 XI11_6/XI0/XI0_62/d__4_ xsel_62_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_3 XI11_6/XI0/XI0_62/d__3_ xsel_62_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_2 XI11_6/XI0/XI0_62/d__2_ xsel_62_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_1 XI11_6/XI0/XI0_62/d__1_ xsel_62_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_0 XI11_6/XI0/XI0_62/d__0_ xsel_62_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_15 XI11_6/net21_0_ xsel_61_ XI11_6/XI0/XI0_61/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_14 XI11_6/net21_1_ xsel_61_ XI11_6/XI0/XI0_61/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_13 XI11_6/net21_2_ xsel_61_ XI11_6/XI0/XI0_61/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_12 XI11_6/net21_3_ xsel_61_ XI11_6/XI0/XI0_61/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_11 XI11_6/net21_4_ xsel_61_ XI11_6/XI0/XI0_61/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_10 XI11_6/net21_5_ xsel_61_ XI11_6/XI0/XI0_61/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_9 XI11_6/net21_6_ xsel_61_ XI11_6/XI0/XI0_61/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_8 XI11_6/net21_7_ xsel_61_ XI11_6/XI0/XI0_61/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_7 XI11_6/net21_8_ xsel_61_ XI11_6/XI0/XI0_61/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_6 XI11_6/net21_9_ xsel_61_ XI11_6/XI0/XI0_61/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_5 XI11_6/net21_10_ xsel_61_ XI11_6/XI0/XI0_61/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_4 XI11_6/net21_11_ xsel_61_ XI11_6/XI0/XI0_61/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_3 XI11_6/net21_12_ xsel_61_ XI11_6/XI0/XI0_61/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_2 XI11_6/net21_13_ xsel_61_ XI11_6/XI0/XI0_61/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_1 XI11_6/net21_14_ xsel_61_ XI11_6/XI0/XI0_61/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_0 XI11_6/net21_15_ xsel_61_ XI11_6/XI0/XI0_61/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_15 XI11_6/XI0/XI0_61/d__15_ xsel_61_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_14 XI11_6/XI0/XI0_61/d__14_ xsel_61_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_13 XI11_6/XI0/XI0_61/d__13_ xsel_61_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_12 XI11_6/XI0/XI0_61/d__12_ xsel_61_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_11 XI11_6/XI0/XI0_61/d__11_ xsel_61_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_10 XI11_6/XI0/XI0_61/d__10_ xsel_61_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_9 XI11_6/XI0/XI0_61/d__9_ xsel_61_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_8 XI11_6/XI0/XI0_61/d__8_ xsel_61_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_7 XI11_6/XI0/XI0_61/d__7_ xsel_61_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_6 XI11_6/XI0/XI0_61/d__6_ xsel_61_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_5 XI11_6/XI0/XI0_61/d__5_ xsel_61_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_4 XI11_6/XI0/XI0_61/d__4_ xsel_61_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_3 XI11_6/XI0/XI0_61/d__3_ xsel_61_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_2 XI11_6/XI0/XI0_61/d__2_ xsel_61_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_1 XI11_6/XI0/XI0_61/d__1_ xsel_61_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_0 XI11_6/XI0/XI0_61/d__0_ xsel_61_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_15 XI11_6/net21_0_ xsel_60_ XI11_6/XI0/XI0_60/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_14 XI11_6/net21_1_ xsel_60_ XI11_6/XI0/XI0_60/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_13 XI11_6/net21_2_ xsel_60_ XI11_6/XI0/XI0_60/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_12 XI11_6/net21_3_ xsel_60_ XI11_6/XI0/XI0_60/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_11 XI11_6/net21_4_ xsel_60_ XI11_6/XI0/XI0_60/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_10 XI11_6/net21_5_ xsel_60_ XI11_6/XI0/XI0_60/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_9 XI11_6/net21_6_ xsel_60_ XI11_6/XI0/XI0_60/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_8 XI11_6/net21_7_ xsel_60_ XI11_6/XI0/XI0_60/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_7 XI11_6/net21_8_ xsel_60_ XI11_6/XI0/XI0_60/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_6 XI11_6/net21_9_ xsel_60_ XI11_6/XI0/XI0_60/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_5 XI11_6/net21_10_ xsel_60_ XI11_6/XI0/XI0_60/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_4 XI11_6/net21_11_ xsel_60_ XI11_6/XI0/XI0_60/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_3 XI11_6/net21_12_ xsel_60_ XI11_6/XI0/XI0_60/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_2 XI11_6/net21_13_ xsel_60_ XI11_6/XI0/XI0_60/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_1 XI11_6/net21_14_ xsel_60_ XI11_6/XI0/XI0_60/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_0 XI11_6/net21_15_ xsel_60_ XI11_6/XI0/XI0_60/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_15 XI11_6/XI0/XI0_60/d__15_ xsel_60_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_14 XI11_6/XI0/XI0_60/d__14_ xsel_60_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_13 XI11_6/XI0/XI0_60/d__13_ xsel_60_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_12 XI11_6/XI0/XI0_60/d__12_ xsel_60_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_11 XI11_6/XI0/XI0_60/d__11_ xsel_60_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_10 XI11_6/XI0/XI0_60/d__10_ xsel_60_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_9 XI11_6/XI0/XI0_60/d__9_ xsel_60_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_8 XI11_6/XI0/XI0_60/d__8_ xsel_60_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_7 XI11_6/XI0/XI0_60/d__7_ xsel_60_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_6 XI11_6/XI0/XI0_60/d__6_ xsel_60_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_5 XI11_6/XI0/XI0_60/d__5_ xsel_60_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_4 XI11_6/XI0/XI0_60/d__4_ xsel_60_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_3 XI11_6/XI0/XI0_60/d__3_ xsel_60_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_2 XI11_6/XI0/XI0_60/d__2_ xsel_60_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_1 XI11_6/XI0/XI0_60/d__1_ xsel_60_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_0 XI11_6/XI0/XI0_60/d__0_ xsel_60_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_15 XI11_6/net21_0_ xsel_59_ XI11_6/XI0/XI0_59/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_14 XI11_6/net21_1_ xsel_59_ XI11_6/XI0/XI0_59/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_13 XI11_6/net21_2_ xsel_59_ XI11_6/XI0/XI0_59/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_12 XI11_6/net21_3_ xsel_59_ XI11_6/XI0/XI0_59/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_11 XI11_6/net21_4_ xsel_59_ XI11_6/XI0/XI0_59/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_10 XI11_6/net21_5_ xsel_59_ XI11_6/XI0/XI0_59/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_9 XI11_6/net21_6_ xsel_59_ XI11_6/XI0/XI0_59/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_8 XI11_6/net21_7_ xsel_59_ XI11_6/XI0/XI0_59/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_7 XI11_6/net21_8_ xsel_59_ XI11_6/XI0/XI0_59/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_6 XI11_6/net21_9_ xsel_59_ XI11_6/XI0/XI0_59/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_5 XI11_6/net21_10_ xsel_59_ XI11_6/XI0/XI0_59/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_4 XI11_6/net21_11_ xsel_59_ XI11_6/XI0/XI0_59/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_3 XI11_6/net21_12_ xsel_59_ XI11_6/XI0/XI0_59/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_2 XI11_6/net21_13_ xsel_59_ XI11_6/XI0/XI0_59/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_1 XI11_6/net21_14_ xsel_59_ XI11_6/XI0/XI0_59/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_0 XI11_6/net21_15_ xsel_59_ XI11_6/XI0/XI0_59/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_15 XI11_6/XI0/XI0_59/d__15_ xsel_59_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_14 XI11_6/XI0/XI0_59/d__14_ xsel_59_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_13 XI11_6/XI0/XI0_59/d__13_ xsel_59_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_12 XI11_6/XI0/XI0_59/d__12_ xsel_59_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_11 XI11_6/XI0/XI0_59/d__11_ xsel_59_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_10 XI11_6/XI0/XI0_59/d__10_ xsel_59_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_9 XI11_6/XI0/XI0_59/d__9_ xsel_59_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_8 XI11_6/XI0/XI0_59/d__8_ xsel_59_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_7 XI11_6/XI0/XI0_59/d__7_ xsel_59_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_6 XI11_6/XI0/XI0_59/d__6_ xsel_59_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_5 XI11_6/XI0/XI0_59/d__5_ xsel_59_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_4 XI11_6/XI0/XI0_59/d__4_ xsel_59_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_3 XI11_6/XI0/XI0_59/d__3_ xsel_59_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_2 XI11_6/XI0/XI0_59/d__2_ xsel_59_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_1 XI11_6/XI0/XI0_59/d__1_ xsel_59_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_0 XI11_6/XI0/XI0_59/d__0_ xsel_59_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_15 XI11_6/net21_0_ xsel_58_ XI11_6/XI0/XI0_58/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_14 XI11_6/net21_1_ xsel_58_ XI11_6/XI0/XI0_58/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_13 XI11_6/net21_2_ xsel_58_ XI11_6/XI0/XI0_58/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_12 XI11_6/net21_3_ xsel_58_ XI11_6/XI0/XI0_58/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_11 XI11_6/net21_4_ xsel_58_ XI11_6/XI0/XI0_58/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_10 XI11_6/net21_5_ xsel_58_ XI11_6/XI0/XI0_58/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_9 XI11_6/net21_6_ xsel_58_ XI11_6/XI0/XI0_58/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_8 XI11_6/net21_7_ xsel_58_ XI11_6/XI0/XI0_58/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_7 XI11_6/net21_8_ xsel_58_ XI11_6/XI0/XI0_58/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_6 XI11_6/net21_9_ xsel_58_ XI11_6/XI0/XI0_58/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_5 XI11_6/net21_10_ xsel_58_ XI11_6/XI0/XI0_58/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_4 XI11_6/net21_11_ xsel_58_ XI11_6/XI0/XI0_58/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_3 XI11_6/net21_12_ xsel_58_ XI11_6/XI0/XI0_58/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_2 XI11_6/net21_13_ xsel_58_ XI11_6/XI0/XI0_58/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_1 XI11_6/net21_14_ xsel_58_ XI11_6/XI0/XI0_58/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_0 XI11_6/net21_15_ xsel_58_ XI11_6/XI0/XI0_58/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_15 XI11_6/XI0/XI0_58/d__15_ xsel_58_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_14 XI11_6/XI0/XI0_58/d__14_ xsel_58_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_13 XI11_6/XI0/XI0_58/d__13_ xsel_58_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_12 XI11_6/XI0/XI0_58/d__12_ xsel_58_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_11 XI11_6/XI0/XI0_58/d__11_ xsel_58_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_10 XI11_6/XI0/XI0_58/d__10_ xsel_58_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_9 XI11_6/XI0/XI0_58/d__9_ xsel_58_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_8 XI11_6/XI0/XI0_58/d__8_ xsel_58_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_7 XI11_6/XI0/XI0_58/d__7_ xsel_58_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_6 XI11_6/XI0/XI0_58/d__6_ xsel_58_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_5 XI11_6/XI0/XI0_58/d__5_ xsel_58_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_4 XI11_6/XI0/XI0_58/d__4_ xsel_58_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_3 XI11_6/XI0/XI0_58/d__3_ xsel_58_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_2 XI11_6/XI0/XI0_58/d__2_ xsel_58_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_1 XI11_6/XI0/XI0_58/d__1_ xsel_58_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_0 XI11_6/XI0/XI0_58/d__0_ xsel_58_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_15 XI11_6/net21_0_ xsel_57_ XI11_6/XI0/XI0_57/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_14 XI11_6/net21_1_ xsel_57_ XI11_6/XI0/XI0_57/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_13 XI11_6/net21_2_ xsel_57_ XI11_6/XI0/XI0_57/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_12 XI11_6/net21_3_ xsel_57_ XI11_6/XI0/XI0_57/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_11 XI11_6/net21_4_ xsel_57_ XI11_6/XI0/XI0_57/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_10 XI11_6/net21_5_ xsel_57_ XI11_6/XI0/XI0_57/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_9 XI11_6/net21_6_ xsel_57_ XI11_6/XI0/XI0_57/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_8 XI11_6/net21_7_ xsel_57_ XI11_6/XI0/XI0_57/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_7 XI11_6/net21_8_ xsel_57_ XI11_6/XI0/XI0_57/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_6 XI11_6/net21_9_ xsel_57_ XI11_6/XI0/XI0_57/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_5 XI11_6/net21_10_ xsel_57_ XI11_6/XI0/XI0_57/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_4 XI11_6/net21_11_ xsel_57_ XI11_6/XI0/XI0_57/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_3 XI11_6/net21_12_ xsel_57_ XI11_6/XI0/XI0_57/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_2 XI11_6/net21_13_ xsel_57_ XI11_6/XI0/XI0_57/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_1 XI11_6/net21_14_ xsel_57_ XI11_6/XI0/XI0_57/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_0 XI11_6/net21_15_ xsel_57_ XI11_6/XI0/XI0_57/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_15 XI11_6/XI0/XI0_57/d__15_ xsel_57_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_14 XI11_6/XI0/XI0_57/d__14_ xsel_57_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_13 XI11_6/XI0/XI0_57/d__13_ xsel_57_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_12 XI11_6/XI0/XI0_57/d__12_ xsel_57_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_11 XI11_6/XI0/XI0_57/d__11_ xsel_57_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_10 XI11_6/XI0/XI0_57/d__10_ xsel_57_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_9 XI11_6/XI0/XI0_57/d__9_ xsel_57_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_8 XI11_6/XI0/XI0_57/d__8_ xsel_57_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_7 XI11_6/XI0/XI0_57/d__7_ xsel_57_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_6 XI11_6/XI0/XI0_57/d__6_ xsel_57_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_5 XI11_6/XI0/XI0_57/d__5_ xsel_57_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_4 XI11_6/XI0/XI0_57/d__4_ xsel_57_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_3 XI11_6/XI0/XI0_57/d__3_ xsel_57_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_2 XI11_6/XI0/XI0_57/d__2_ xsel_57_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_1 XI11_6/XI0/XI0_57/d__1_ xsel_57_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_0 XI11_6/XI0/XI0_57/d__0_ xsel_57_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_15 XI11_6/net21_0_ xsel_56_ XI11_6/XI0/XI0_56/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_14 XI11_6/net21_1_ xsel_56_ XI11_6/XI0/XI0_56/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_13 XI11_6/net21_2_ xsel_56_ XI11_6/XI0/XI0_56/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_12 XI11_6/net21_3_ xsel_56_ XI11_6/XI0/XI0_56/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_11 XI11_6/net21_4_ xsel_56_ XI11_6/XI0/XI0_56/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_10 XI11_6/net21_5_ xsel_56_ XI11_6/XI0/XI0_56/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_9 XI11_6/net21_6_ xsel_56_ XI11_6/XI0/XI0_56/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_8 XI11_6/net21_7_ xsel_56_ XI11_6/XI0/XI0_56/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_7 XI11_6/net21_8_ xsel_56_ XI11_6/XI0/XI0_56/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_6 XI11_6/net21_9_ xsel_56_ XI11_6/XI0/XI0_56/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_5 XI11_6/net21_10_ xsel_56_ XI11_6/XI0/XI0_56/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_4 XI11_6/net21_11_ xsel_56_ XI11_6/XI0/XI0_56/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_3 XI11_6/net21_12_ xsel_56_ XI11_6/XI0/XI0_56/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_2 XI11_6/net21_13_ xsel_56_ XI11_6/XI0/XI0_56/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_1 XI11_6/net21_14_ xsel_56_ XI11_6/XI0/XI0_56/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_0 XI11_6/net21_15_ xsel_56_ XI11_6/XI0/XI0_56/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_15 XI11_6/XI0/XI0_56/d__15_ xsel_56_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_14 XI11_6/XI0/XI0_56/d__14_ xsel_56_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_13 XI11_6/XI0/XI0_56/d__13_ xsel_56_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_12 XI11_6/XI0/XI0_56/d__12_ xsel_56_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_11 XI11_6/XI0/XI0_56/d__11_ xsel_56_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_10 XI11_6/XI0/XI0_56/d__10_ xsel_56_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_9 XI11_6/XI0/XI0_56/d__9_ xsel_56_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_8 XI11_6/XI0/XI0_56/d__8_ xsel_56_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_7 XI11_6/XI0/XI0_56/d__7_ xsel_56_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_6 XI11_6/XI0/XI0_56/d__6_ xsel_56_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_5 XI11_6/XI0/XI0_56/d__5_ xsel_56_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_4 XI11_6/XI0/XI0_56/d__4_ xsel_56_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_3 XI11_6/XI0/XI0_56/d__3_ xsel_56_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_2 XI11_6/XI0/XI0_56/d__2_ xsel_56_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_1 XI11_6/XI0/XI0_56/d__1_ xsel_56_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_0 XI11_6/XI0/XI0_56/d__0_ xsel_56_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_15 XI11_6/net21_0_ xsel_55_ XI11_6/XI0/XI0_55/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_14 XI11_6/net21_1_ xsel_55_ XI11_6/XI0/XI0_55/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_13 XI11_6/net21_2_ xsel_55_ XI11_6/XI0/XI0_55/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_12 XI11_6/net21_3_ xsel_55_ XI11_6/XI0/XI0_55/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_11 XI11_6/net21_4_ xsel_55_ XI11_6/XI0/XI0_55/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_10 XI11_6/net21_5_ xsel_55_ XI11_6/XI0/XI0_55/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_9 XI11_6/net21_6_ xsel_55_ XI11_6/XI0/XI0_55/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_8 XI11_6/net21_7_ xsel_55_ XI11_6/XI0/XI0_55/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_7 XI11_6/net21_8_ xsel_55_ XI11_6/XI0/XI0_55/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_6 XI11_6/net21_9_ xsel_55_ XI11_6/XI0/XI0_55/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_5 XI11_6/net21_10_ xsel_55_ XI11_6/XI0/XI0_55/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_4 XI11_6/net21_11_ xsel_55_ XI11_6/XI0/XI0_55/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_3 XI11_6/net21_12_ xsel_55_ XI11_6/XI0/XI0_55/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_2 XI11_6/net21_13_ xsel_55_ XI11_6/XI0/XI0_55/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_1 XI11_6/net21_14_ xsel_55_ XI11_6/XI0/XI0_55/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_0 XI11_6/net21_15_ xsel_55_ XI11_6/XI0/XI0_55/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_15 XI11_6/XI0/XI0_55/d__15_ xsel_55_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_14 XI11_6/XI0/XI0_55/d__14_ xsel_55_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_13 XI11_6/XI0/XI0_55/d__13_ xsel_55_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_12 XI11_6/XI0/XI0_55/d__12_ xsel_55_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_11 XI11_6/XI0/XI0_55/d__11_ xsel_55_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_10 XI11_6/XI0/XI0_55/d__10_ xsel_55_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_9 XI11_6/XI0/XI0_55/d__9_ xsel_55_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_8 XI11_6/XI0/XI0_55/d__8_ xsel_55_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_7 XI11_6/XI0/XI0_55/d__7_ xsel_55_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_6 XI11_6/XI0/XI0_55/d__6_ xsel_55_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_5 XI11_6/XI0/XI0_55/d__5_ xsel_55_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_4 XI11_6/XI0/XI0_55/d__4_ xsel_55_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_3 XI11_6/XI0/XI0_55/d__3_ xsel_55_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_2 XI11_6/XI0/XI0_55/d__2_ xsel_55_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_1 XI11_6/XI0/XI0_55/d__1_ xsel_55_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_0 XI11_6/XI0/XI0_55/d__0_ xsel_55_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_15 XI11_6/net21_0_ xsel_54_ XI11_6/XI0/XI0_54/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_14 XI11_6/net21_1_ xsel_54_ XI11_6/XI0/XI0_54/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_13 XI11_6/net21_2_ xsel_54_ XI11_6/XI0/XI0_54/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_12 XI11_6/net21_3_ xsel_54_ XI11_6/XI0/XI0_54/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_11 XI11_6/net21_4_ xsel_54_ XI11_6/XI0/XI0_54/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_10 XI11_6/net21_5_ xsel_54_ XI11_6/XI0/XI0_54/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_9 XI11_6/net21_6_ xsel_54_ XI11_6/XI0/XI0_54/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_8 XI11_6/net21_7_ xsel_54_ XI11_6/XI0/XI0_54/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_7 XI11_6/net21_8_ xsel_54_ XI11_6/XI0/XI0_54/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_6 XI11_6/net21_9_ xsel_54_ XI11_6/XI0/XI0_54/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_5 XI11_6/net21_10_ xsel_54_ XI11_6/XI0/XI0_54/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_4 XI11_6/net21_11_ xsel_54_ XI11_6/XI0/XI0_54/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_3 XI11_6/net21_12_ xsel_54_ XI11_6/XI0/XI0_54/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_2 XI11_6/net21_13_ xsel_54_ XI11_6/XI0/XI0_54/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_1 XI11_6/net21_14_ xsel_54_ XI11_6/XI0/XI0_54/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_0 XI11_6/net21_15_ xsel_54_ XI11_6/XI0/XI0_54/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_15 XI11_6/XI0/XI0_54/d__15_ xsel_54_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_14 XI11_6/XI0/XI0_54/d__14_ xsel_54_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_13 XI11_6/XI0/XI0_54/d__13_ xsel_54_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_12 XI11_6/XI0/XI0_54/d__12_ xsel_54_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_11 XI11_6/XI0/XI0_54/d__11_ xsel_54_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_10 XI11_6/XI0/XI0_54/d__10_ xsel_54_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_9 XI11_6/XI0/XI0_54/d__9_ xsel_54_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_8 XI11_6/XI0/XI0_54/d__8_ xsel_54_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_7 XI11_6/XI0/XI0_54/d__7_ xsel_54_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_6 XI11_6/XI0/XI0_54/d__6_ xsel_54_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_5 XI11_6/XI0/XI0_54/d__5_ xsel_54_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_4 XI11_6/XI0/XI0_54/d__4_ xsel_54_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_3 XI11_6/XI0/XI0_54/d__3_ xsel_54_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_2 XI11_6/XI0/XI0_54/d__2_ xsel_54_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_1 XI11_6/XI0/XI0_54/d__1_ xsel_54_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_0 XI11_6/XI0/XI0_54/d__0_ xsel_54_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_15 XI11_6/net21_0_ xsel_53_ XI11_6/XI0/XI0_53/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_14 XI11_6/net21_1_ xsel_53_ XI11_6/XI0/XI0_53/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_13 XI11_6/net21_2_ xsel_53_ XI11_6/XI0/XI0_53/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_12 XI11_6/net21_3_ xsel_53_ XI11_6/XI0/XI0_53/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_11 XI11_6/net21_4_ xsel_53_ XI11_6/XI0/XI0_53/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_10 XI11_6/net21_5_ xsel_53_ XI11_6/XI0/XI0_53/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_9 XI11_6/net21_6_ xsel_53_ XI11_6/XI0/XI0_53/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_8 XI11_6/net21_7_ xsel_53_ XI11_6/XI0/XI0_53/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_7 XI11_6/net21_8_ xsel_53_ XI11_6/XI0/XI0_53/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_6 XI11_6/net21_9_ xsel_53_ XI11_6/XI0/XI0_53/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_5 XI11_6/net21_10_ xsel_53_ XI11_6/XI0/XI0_53/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_4 XI11_6/net21_11_ xsel_53_ XI11_6/XI0/XI0_53/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_3 XI11_6/net21_12_ xsel_53_ XI11_6/XI0/XI0_53/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_2 XI11_6/net21_13_ xsel_53_ XI11_6/XI0/XI0_53/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_1 XI11_6/net21_14_ xsel_53_ XI11_6/XI0/XI0_53/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_0 XI11_6/net21_15_ xsel_53_ XI11_6/XI0/XI0_53/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_15 XI11_6/XI0/XI0_53/d__15_ xsel_53_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_14 XI11_6/XI0/XI0_53/d__14_ xsel_53_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_13 XI11_6/XI0/XI0_53/d__13_ xsel_53_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_12 XI11_6/XI0/XI0_53/d__12_ xsel_53_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_11 XI11_6/XI0/XI0_53/d__11_ xsel_53_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_10 XI11_6/XI0/XI0_53/d__10_ xsel_53_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_9 XI11_6/XI0/XI0_53/d__9_ xsel_53_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_8 XI11_6/XI0/XI0_53/d__8_ xsel_53_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_7 XI11_6/XI0/XI0_53/d__7_ xsel_53_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_6 XI11_6/XI0/XI0_53/d__6_ xsel_53_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_5 XI11_6/XI0/XI0_53/d__5_ xsel_53_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_4 XI11_6/XI0/XI0_53/d__4_ xsel_53_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_3 XI11_6/XI0/XI0_53/d__3_ xsel_53_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_2 XI11_6/XI0/XI0_53/d__2_ xsel_53_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_1 XI11_6/XI0/XI0_53/d__1_ xsel_53_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_0 XI11_6/XI0/XI0_53/d__0_ xsel_53_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_15 XI11_6/net21_0_ xsel_52_ XI11_6/XI0/XI0_52/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_14 XI11_6/net21_1_ xsel_52_ XI11_6/XI0/XI0_52/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_13 XI11_6/net21_2_ xsel_52_ XI11_6/XI0/XI0_52/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_12 XI11_6/net21_3_ xsel_52_ XI11_6/XI0/XI0_52/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_11 XI11_6/net21_4_ xsel_52_ XI11_6/XI0/XI0_52/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_10 XI11_6/net21_5_ xsel_52_ XI11_6/XI0/XI0_52/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_9 XI11_6/net21_6_ xsel_52_ XI11_6/XI0/XI0_52/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_8 XI11_6/net21_7_ xsel_52_ XI11_6/XI0/XI0_52/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_7 XI11_6/net21_8_ xsel_52_ XI11_6/XI0/XI0_52/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_6 XI11_6/net21_9_ xsel_52_ XI11_6/XI0/XI0_52/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_5 XI11_6/net21_10_ xsel_52_ XI11_6/XI0/XI0_52/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_4 XI11_6/net21_11_ xsel_52_ XI11_6/XI0/XI0_52/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_3 XI11_6/net21_12_ xsel_52_ XI11_6/XI0/XI0_52/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_2 XI11_6/net21_13_ xsel_52_ XI11_6/XI0/XI0_52/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_1 XI11_6/net21_14_ xsel_52_ XI11_6/XI0/XI0_52/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_0 XI11_6/net21_15_ xsel_52_ XI11_6/XI0/XI0_52/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_15 XI11_6/XI0/XI0_52/d__15_ xsel_52_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_14 XI11_6/XI0/XI0_52/d__14_ xsel_52_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_13 XI11_6/XI0/XI0_52/d__13_ xsel_52_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_12 XI11_6/XI0/XI0_52/d__12_ xsel_52_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_11 XI11_6/XI0/XI0_52/d__11_ xsel_52_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_10 XI11_6/XI0/XI0_52/d__10_ xsel_52_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_9 XI11_6/XI0/XI0_52/d__9_ xsel_52_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_8 XI11_6/XI0/XI0_52/d__8_ xsel_52_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_7 XI11_6/XI0/XI0_52/d__7_ xsel_52_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_6 XI11_6/XI0/XI0_52/d__6_ xsel_52_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_5 XI11_6/XI0/XI0_52/d__5_ xsel_52_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_4 XI11_6/XI0/XI0_52/d__4_ xsel_52_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_3 XI11_6/XI0/XI0_52/d__3_ xsel_52_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_2 XI11_6/XI0/XI0_52/d__2_ xsel_52_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_1 XI11_6/XI0/XI0_52/d__1_ xsel_52_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_0 XI11_6/XI0/XI0_52/d__0_ xsel_52_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_15 XI11_6/net21_0_ xsel_51_ XI11_6/XI0/XI0_51/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_14 XI11_6/net21_1_ xsel_51_ XI11_6/XI0/XI0_51/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_13 XI11_6/net21_2_ xsel_51_ XI11_6/XI0/XI0_51/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_12 XI11_6/net21_3_ xsel_51_ XI11_6/XI0/XI0_51/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_11 XI11_6/net21_4_ xsel_51_ XI11_6/XI0/XI0_51/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_10 XI11_6/net21_5_ xsel_51_ XI11_6/XI0/XI0_51/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_9 XI11_6/net21_6_ xsel_51_ XI11_6/XI0/XI0_51/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_8 XI11_6/net21_7_ xsel_51_ XI11_6/XI0/XI0_51/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_7 XI11_6/net21_8_ xsel_51_ XI11_6/XI0/XI0_51/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_6 XI11_6/net21_9_ xsel_51_ XI11_6/XI0/XI0_51/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_5 XI11_6/net21_10_ xsel_51_ XI11_6/XI0/XI0_51/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_4 XI11_6/net21_11_ xsel_51_ XI11_6/XI0/XI0_51/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_3 XI11_6/net21_12_ xsel_51_ XI11_6/XI0/XI0_51/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_2 XI11_6/net21_13_ xsel_51_ XI11_6/XI0/XI0_51/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_1 XI11_6/net21_14_ xsel_51_ XI11_6/XI0/XI0_51/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_0 XI11_6/net21_15_ xsel_51_ XI11_6/XI0/XI0_51/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_15 XI11_6/XI0/XI0_51/d__15_ xsel_51_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_14 XI11_6/XI0/XI0_51/d__14_ xsel_51_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_13 XI11_6/XI0/XI0_51/d__13_ xsel_51_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_12 XI11_6/XI0/XI0_51/d__12_ xsel_51_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_11 XI11_6/XI0/XI0_51/d__11_ xsel_51_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_10 XI11_6/XI0/XI0_51/d__10_ xsel_51_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_9 XI11_6/XI0/XI0_51/d__9_ xsel_51_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_8 XI11_6/XI0/XI0_51/d__8_ xsel_51_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_7 XI11_6/XI0/XI0_51/d__7_ xsel_51_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_6 XI11_6/XI0/XI0_51/d__6_ xsel_51_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_5 XI11_6/XI0/XI0_51/d__5_ xsel_51_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_4 XI11_6/XI0/XI0_51/d__4_ xsel_51_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_3 XI11_6/XI0/XI0_51/d__3_ xsel_51_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_2 XI11_6/XI0/XI0_51/d__2_ xsel_51_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_1 XI11_6/XI0/XI0_51/d__1_ xsel_51_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_0 XI11_6/XI0/XI0_51/d__0_ xsel_51_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_15 XI11_6/net21_0_ xsel_50_ XI11_6/XI0/XI0_50/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_14 XI11_6/net21_1_ xsel_50_ XI11_6/XI0/XI0_50/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_13 XI11_6/net21_2_ xsel_50_ XI11_6/XI0/XI0_50/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_12 XI11_6/net21_3_ xsel_50_ XI11_6/XI0/XI0_50/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_11 XI11_6/net21_4_ xsel_50_ XI11_6/XI0/XI0_50/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_10 XI11_6/net21_5_ xsel_50_ XI11_6/XI0/XI0_50/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_9 XI11_6/net21_6_ xsel_50_ XI11_6/XI0/XI0_50/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_8 XI11_6/net21_7_ xsel_50_ XI11_6/XI0/XI0_50/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_7 XI11_6/net21_8_ xsel_50_ XI11_6/XI0/XI0_50/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_6 XI11_6/net21_9_ xsel_50_ XI11_6/XI0/XI0_50/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_5 XI11_6/net21_10_ xsel_50_ XI11_6/XI0/XI0_50/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_4 XI11_6/net21_11_ xsel_50_ XI11_6/XI0/XI0_50/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_3 XI11_6/net21_12_ xsel_50_ XI11_6/XI0/XI0_50/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_2 XI11_6/net21_13_ xsel_50_ XI11_6/XI0/XI0_50/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_1 XI11_6/net21_14_ xsel_50_ XI11_6/XI0/XI0_50/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_0 XI11_6/net21_15_ xsel_50_ XI11_6/XI0/XI0_50/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_15 XI11_6/XI0/XI0_50/d__15_ xsel_50_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_14 XI11_6/XI0/XI0_50/d__14_ xsel_50_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_13 XI11_6/XI0/XI0_50/d__13_ xsel_50_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_12 XI11_6/XI0/XI0_50/d__12_ xsel_50_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_11 XI11_6/XI0/XI0_50/d__11_ xsel_50_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_10 XI11_6/XI0/XI0_50/d__10_ xsel_50_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_9 XI11_6/XI0/XI0_50/d__9_ xsel_50_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_8 XI11_6/XI0/XI0_50/d__8_ xsel_50_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_7 XI11_6/XI0/XI0_50/d__7_ xsel_50_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_6 XI11_6/XI0/XI0_50/d__6_ xsel_50_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_5 XI11_6/XI0/XI0_50/d__5_ xsel_50_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_4 XI11_6/XI0/XI0_50/d__4_ xsel_50_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_3 XI11_6/XI0/XI0_50/d__3_ xsel_50_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_2 XI11_6/XI0/XI0_50/d__2_ xsel_50_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_1 XI11_6/XI0/XI0_50/d__1_ xsel_50_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_0 XI11_6/XI0/XI0_50/d__0_ xsel_50_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_15 XI11_6/net21_0_ xsel_49_ XI11_6/XI0/XI0_49/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_14 XI11_6/net21_1_ xsel_49_ XI11_6/XI0/XI0_49/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_13 XI11_6/net21_2_ xsel_49_ XI11_6/XI0/XI0_49/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_12 XI11_6/net21_3_ xsel_49_ XI11_6/XI0/XI0_49/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_11 XI11_6/net21_4_ xsel_49_ XI11_6/XI0/XI0_49/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_10 XI11_6/net21_5_ xsel_49_ XI11_6/XI0/XI0_49/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_9 XI11_6/net21_6_ xsel_49_ XI11_6/XI0/XI0_49/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_8 XI11_6/net21_7_ xsel_49_ XI11_6/XI0/XI0_49/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_7 XI11_6/net21_8_ xsel_49_ XI11_6/XI0/XI0_49/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_6 XI11_6/net21_9_ xsel_49_ XI11_6/XI0/XI0_49/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_5 XI11_6/net21_10_ xsel_49_ XI11_6/XI0/XI0_49/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_4 XI11_6/net21_11_ xsel_49_ XI11_6/XI0/XI0_49/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_3 XI11_6/net21_12_ xsel_49_ XI11_6/XI0/XI0_49/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_2 XI11_6/net21_13_ xsel_49_ XI11_6/XI0/XI0_49/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_1 XI11_6/net21_14_ xsel_49_ XI11_6/XI0/XI0_49/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_0 XI11_6/net21_15_ xsel_49_ XI11_6/XI0/XI0_49/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_15 XI11_6/XI0/XI0_49/d__15_ xsel_49_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_14 XI11_6/XI0/XI0_49/d__14_ xsel_49_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_13 XI11_6/XI0/XI0_49/d__13_ xsel_49_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_12 XI11_6/XI0/XI0_49/d__12_ xsel_49_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_11 XI11_6/XI0/XI0_49/d__11_ xsel_49_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_10 XI11_6/XI0/XI0_49/d__10_ xsel_49_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_9 XI11_6/XI0/XI0_49/d__9_ xsel_49_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_8 XI11_6/XI0/XI0_49/d__8_ xsel_49_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_7 XI11_6/XI0/XI0_49/d__7_ xsel_49_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_6 XI11_6/XI0/XI0_49/d__6_ xsel_49_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_5 XI11_6/XI0/XI0_49/d__5_ xsel_49_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_4 XI11_6/XI0/XI0_49/d__4_ xsel_49_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_3 XI11_6/XI0/XI0_49/d__3_ xsel_49_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_2 XI11_6/XI0/XI0_49/d__2_ xsel_49_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_1 XI11_6/XI0/XI0_49/d__1_ xsel_49_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_0 XI11_6/XI0/XI0_49/d__0_ xsel_49_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_15 XI11_6/net21_0_ xsel_48_ XI11_6/XI0/XI0_48/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_14 XI11_6/net21_1_ xsel_48_ XI11_6/XI0/XI0_48/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_13 XI11_6/net21_2_ xsel_48_ XI11_6/XI0/XI0_48/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_12 XI11_6/net21_3_ xsel_48_ XI11_6/XI0/XI0_48/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_11 XI11_6/net21_4_ xsel_48_ XI11_6/XI0/XI0_48/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_10 XI11_6/net21_5_ xsel_48_ XI11_6/XI0/XI0_48/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_9 XI11_6/net21_6_ xsel_48_ XI11_6/XI0/XI0_48/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_8 XI11_6/net21_7_ xsel_48_ XI11_6/XI0/XI0_48/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_7 XI11_6/net21_8_ xsel_48_ XI11_6/XI0/XI0_48/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_6 XI11_6/net21_9_ xsel_48_ XI11_6/XI0/XI0_48/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_5 XI11_6/net21_10_ xsel_48_ XI11_6/XI0/XI0_48/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_4 XI11_6/net21_11_ xsel_48_ XI11_6/XI0/XI0_48/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_3 XI11_6/net21_12_ xsel_48_ XI11_6/XI0/XI0_48/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_2 XI11_6/net21_13_ xsel_48_ XI11_6/XI0/XI0_48/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_1 XI11_6/net21_14_ xsel_48_ XI11_6/XI0/XI0_48/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_0 XI11_6/net21_15_ xsel_48_ XI11_6/XI0/XI0_48/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_15 XI11_6/XI0/XI0_48/d__15_ xsel_48_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_14 XI11_6/XI0/XI0_48/d__14_ xsel_48_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_13 XI11_6/XI0/XI0_48/d__13_ xsel_48_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_12 XI11_6/XI0/XI0_48/d__12_ xsel_48_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_11 XI11_6/XI0/XI0_48/d__11_ xsel_48_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_10 XI11_6/XI0/XI0_48/d__10_ xsel_48_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_9 XI11_6/XI0/XI0_48/d__9_ xsel_48_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_8 XI11_6/XI0/XI0_48/d__8_ xsel_48_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_7 XI11_6/XI0/XI0_48/d__7_ xsel_48_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_6 XI11_6/XI0/XI0_48/d__6_ xsel_48_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_5 XI11_6/XI0/XI0_48/d__5_ xsel_48_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_4 XI11_6/XI0/XI0_48/d__4_ xsel_48_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_3 XI11_6/XI0/XI0_48/d__3_ xsel_48_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_2 XI11_6/XI0/XI0_48/d__2_ xsel_48_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_1 XI11_6/XI0/XI0_48/d__1_ xsel_48_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_0 XI11_6/XI0/XI0_48/d__0_ xsel_48_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_15 XI11_6/net21_0_ xsel_47_ XI11_6/XI0/XI0_47/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_14 XI11_6/net21_1_ xsel_47_ XI11_6/XI0/XI0_47/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_13 XI11_6/net21_2_ xsel_47_ XI11_6/XI0/XI0_47/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_12 XI11_6/net21_3_ xsel_47_ XI11_6/XI0/XI0_47/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_11 XI11_6/net21_4_ xsel_47_ XI11_6/XI0/XI0_47/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_10 XI11_6/net21_5_ xsel_47_ XI11_6/XI0/XI0_47/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_9 XI11_6/net21_6_ xsel_47_ XI11_6/XI0/XI0_47/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_8 XI11_6/net21_7_ xsel_47_ XI11_6/XI0/XI0_47/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_7 XI11_6/net21_8_ xsel_47_ XI11_6/XI0/XI0_47/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_6 XI11_6/net21_9_ xsel_47_ XI11_6/XI0/XI0_47/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_5 XI11_6/net21_10_ xsel_47_ XI11_6/XI0/XI0_47/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_4 XI11_6/net21_11_ xsel_47_ XI11_6/XI0/XI0_47/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_3 XI11_6/net21_12_ xsel_47_ XI11_6/XI0/XI0_47/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_2 XI11_6/net21_13_ xsel_47_ XI11_6/XI0/XI0_47/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_1 XI11_6/net21_14_ xsel_47_ XI11_6/XI0/XI0_47/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_0 XI11_6/net21_15_ xsel_47_ XI11_6/XI0/XI0_47/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_15 XI11_6/XI0/XI0_47/d__15_ xsel_47_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_14 XI11_6/XI0/XI0_47/d__14_ xsel_47_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_13 XI11_6/XI0/XI0_47/d__13_ xsel_47_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_12 XI11_6/XI0/XI0_47/d__12_ xsel_47_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_11 XI11_6/XI0/XI0_47/d__11_ xsel_47_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_10 XI11_6/XI0/XI0_47/d__10_ xsel_47_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_9 XI11_6/XI0/XI0_47/d__9_ xsel_47_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_8 XI11_6/XI0/XI0_47/d__8_ xsel_47_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_7 XI11_6/XI0/XI0_47/d__7_ xsel_47_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_6 XI11_6/XI0/XI0_47/d__6_ xsel_47_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_5 XI11_6/XI0/XI0_47/d__5_ xsel_47_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_4 XI11_6/XI0/XI0_47/d__4_ xsel_47_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_3 XI11_6/XI0/XI0_47/d__3_ xsel_47_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_2 XI11_6/XI0/XI0_47/d__2_ xsel_47_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_1 XI11_6/XI0/XI0_47/d__1_ xsel_47_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_0 XI11_6/XI0/XI0_47/d__0_ xsel_47_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_15 XI11_6/net21_0_ xsel_46_ XI11_6/XI0/XI0_46/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_14 XI11_6/net21_1_ xsel_46_ XI11_6/XI0/XI0_46/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_13 XI11_6/net21_2_ xsel_46_ XI11_6/XI0/XI0_46/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_12 XI11_6/net21_3_ xsel_46_ XI11_6/XI0/XI0_46/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_11 XI11_6/net21_4_ xsel_46_ XI11_6/XI0/XI0_46/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_10 XI11_6/net21_5_ xsel_46_ XI11_6/XI0/XI0_46/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_9 XI11_6/net21_6_ xsel_46_ XI11_6/XI0/XI0_46/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_8 XI11_6/net21_7_ xsel_46_ XI11_6/XI0/XI0_46/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_7 XI11_6/net21_8_ xsel_46_ XI11_6/XI0/XI0_46/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_6 XI11_6/net21_9_ xsel_46_ XI11_6/XI0/XI0_46/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_5 XI11_6/net21_10_ xsel_46_ XI11_6/XI0/XI0_46/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_4 XI11_6/net21_11_ xsel_46_ XI11_6/XI0/XI0_46/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_3 XI11_6/net21_12_ xsel_46_ XI11_6/XI0/XI0_46/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_2 XI11_6/net21_13_ xsel_46_ XI11_6/XI0/XI0_46/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_1 XI11_6/net21_14_ xsel_46_ XI11_6/XI0/XI0_46/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_0 XI11_6/net21_15_ xsel_46_ XI11_6/XI0/XI0_46/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_15 XI11_6/XI0/XI0_46/d__15_ xsel_46_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_14 XI11_6/XI0/XI0_46/d__14_ xsel_46_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_13 XI11_6/XI0/XI0_46/d__13_ xsel_46_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_12 XI11_6/XI0/XI0_46/d__12_ xsel_46_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_11 XI11_6/XI0/XI0_46/d__11_ xsel_46_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_10 XI11_6/XI0/XI0_46/d__10_ xsel_46_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_9 XI11_6/XI0/XI0_46/d__9_ xsel_46_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_8 XI11_6/XI0/XI0_46/d__8_ xsel_46_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_7 XI11_6/XI0/XI0_46/d__7_ xsel_46_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_6 XI11_6/XI0/XI0_46/d__6_ xsel_46_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_5 XI11_6/XI0/XI0_46/d__5_ xsel_46_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_4 XI11_6/XI0/XI0_46/d__4_ xsel_46_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_3 XI11_6/XI0/XI0_46/d__3_ xsel_46_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_2 XI11_6/XI0/XI0_46/d__2_ xsel_46_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_1 XI11_6/XI0/XI0_46/d__1_ xsel_46_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_0 XI11_6/XI0/XI0_46/d__0_ xsel_46_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_15 XI11_6/net21_0_ xsel_45_ XI11_6/XI0/XI0_45/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_14 XI11_6/net21_1_ xsel_45_ XI11_6/XI0/XI0_45/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_13 XI11_6/net21_2_ xsel_45_ XI11_6/XI0/XI0_45/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_12 XI11_6/net21_3_ xsel_45_ XI11_6/XI0/XI0_45/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_11 XI11_6/net21_4_ xsel_45_ XI11_6/XI0/XI0_45/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_10 XI11_6/net21_5_ xsel_45_ XI11_6/XI0/XI0_45/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_9 XI11_6/net21_6_ xsel_45_ XI11_6/XI0/XI0_45/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_8 XI11_6/net21_7_ xsel_45_ XI11_6/XI0/XI0_45/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_7 XI11_6/net21_8_ xsel_45_ XI11_6/XI0/XI0_45/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_6 XI11_6/net21_9_ xsel_45_ XI11_6/XI0/XI0_45/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_5 XI11_6/net21_10_ xsel_45_ XI11_6/XI0/XI0_45/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_4 XI11_6/net21_11_ xsel_45_ XI11_6/XI0/XI0_45/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_3 XI11_6/net21_12_ xsel_45_ XI11_6/XI0/XI0_45/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_2 XI11_6/net21_13_ xsel_45_ XI11_6/XI0/XI0_45/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_1 XI11_6/net21_14_ xsel_45_ XI11_6/XI0/XI0_45/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_0 XI11_6/net21_15_ xsel_45_ XI11_6/XI0/XI0_45/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_15 XI11_6/XI0/XI0_45/d__15_ xsel_45_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_14 XI11_6/XI0/XI0_45/d__14_ xsel_45_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_13 XI11_6/XI0/XI0_45/d__13_ xsel_45_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_12 XI11_6/XI0/XI0_45/d__12_ xsel_45_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_11 XI11_6/XI0/XI0_45/d__11_ xsel_45_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_10 XI11_6/XI0/XI0_45/d__10_ xsel_45_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_9 XI11_6/XI0/XI0_45/d__9_ xsel_45_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_8 XI11_6/XI0/XI0_45/d__8_ xsel_45_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_7 XI11_6/XI0/XI0_45/d__7_ xsel_45_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_6 XI11_6/XI0/XI0_45/d__6_ xsel_45_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_5 XI11_6/XI0/XI0_45/d__5_ xsel_45_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_4 XI11_6/XI0/XI0_45/d__4_ xsel_45_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_3 XI11_6/XI0/XI0_45/d__3_ xsel_45_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_2 XI11_6/XI0/XI0_45/d__2_ xsel_45_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_1 XI11_6/XI0/XI0_45/d__1_ xsel_45_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_0 XI11_6/XI0/XI0_45/d__0_ xsel_45_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_15 XI11_6/net21_0_ xsel_44_ XI11_6/XI0/XI0_44/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_14 XI11_6/net21_1_ xsel_44_ XI11_6/XI0/XI0_44/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_13 XI11_6/net21_2_ xsel_44_ XI11_6/XI0/XI0_44/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_12 XI11_6/net21_3_ xsel_44_ XI11_6/XI0/XI0_44/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_11 XI11_6/net21_4_ xsel_44_ XI11_6/XI0/XI0_44/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_10 XI11_6/net21_5_ xsel_44_ XI11_6/XI0/XI0_44/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_9 XI11_6/net21_6_ xsel_44_ XI11_6/XI0/XI0_44/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_8 XI11_6/net21_7_ xsel_44_ XI11_6/XI0/XI0_44/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_7 XI11_6/net21_8_ xsel_44_ XI11_6/XI0/XI0_44/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_6 XI11_6/net21_9_ xsel_44_ XI11_6/XI0/XI0_44/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_5 XI11_6/net21_10_ xsel_44_ XI11_6/XI0/XI0_44/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_4 XI11_6/net21_11_ xsel_44_ XI11_6/XI0/XI0_44/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_3 XI11_6/net21_12_ xsel_44_ XI11_6/XI0/XI0_44/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_2 XI11_6/net21_13_ xsel_44_ XI11_6/XI0/XI0_44/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_1 XI11_6/net21_14_ xsel_44_ XI11_6/XI0/XI0_44/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_0 XI11_6/net21_15_ xsel_44_ XI11_6/XI0/XI0_44/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_15 XI11_6/XI0/XI0_44/d__15_ xsel_44_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_14 XI11_6/XI0/XI0_44/d__14_ xsel_44_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_13 XI11_6/XI0/XI0_44/d__13_ xsel_44_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_12 XI11_6/XI0/XI0_44/d__12_ xsel_44_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_11 XI11_6/XI0/XI0_44/d__11_ xsel_44_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_10 XI11_6/XI0/XI0_44/d__10_ xsel_44_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_9 XI11_6/XI0/XI0_44/d__9_ xsel_44_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_8 XI11_6/XI0/XI0_44/d__8_ xsel_44_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_7 XI11_6/XI0/XI0_44/d__7_ xsel_44_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_6 XI11_6/XI0/XI0_44/d__6_ xsel_44_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_5 XI11_6/XI0/XI0_44/d__5_ xsel_44_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_4 XI11_6/XI0/XI0_44/d__4_ xsel_44_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_3 XI11_6/XI0/XI0_44/d__3_ xsel_44_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_2 XI11_6/XI0/XI0_44/d__2_ xsel_44_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_1 XI11_6/XI0/XI0_44/d__1_ xsel_44_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_0 XI11_6/XI0/XI0_44/d__0_ xsel_44_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_15 XI11_6/net21_0_ xsel_43_ XI11_6/XI0/XI0_43/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_14 XI11_6/net21_1_ xsel_43_ XI11_6/XI0/XI0_43/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_13 XI11_6/net21_2_ xsel_43_ XI11_6/XI0/XI0_43/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_12 XI11_6/net21_3_ xsel_43_ XI11_6/XI0/XI0_43/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_11 XI11_6/net21_4_ xsel_43_ XI11_6/XI0/XI0_43/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_10 XI11_6/net21_5_ xsel_43_ XI11_6/XI0/XI0_43/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_9 XI11_6/net21_6_ xsel_43_ XI11_6/XI0/XI0_43/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_8 XI11_6/net21_7_ xsel_43_ XI11_6/XI0/XI0_43/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_7 XI11_6/net21_8_ xsel_43_ XI11_6/XI0/XI0_43/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_6 XI11_6/net21_9_ xsel_43_ XI11_6/XI0/XI0_43/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_5 XI11_6/net21_10_ xsel_43_ XI11_6/XI0/XI0_43/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_4 XI11_6/net21_11_ xsel_43_ XI11_6/XI0/XI0_43/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_3 XI11_6/net21_12_ xsel_43_ XI11_6/XI0/XI0_43/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_2 XI11_6/net21_13_ xsel_43_ XI11_6/XI0/XI0_43/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_1 XI11_6/net21_14_ xsel_43_ XI11_6/XI0/XI0_43/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_0 XI11_6/net21_15_ xsel_43_ XI11_6/XI0/XI0_43/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_15 XI11_6/XI0/XI0_43/d__15_ xsel_43_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_14 XI11_6/XI0/XI0_43/d__14_ xsel_43_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_13 XI11_6/XI0/XI0_43/d__13_ xsel_43_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_12 XI11_6/XI0/XI0_43/d__12_ xsel_43_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_11 XI11_6/XI0/XI0_43/d__11_ xsel_43_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_10 XI11_6/XI0/XI0_43/d__10_ xsel_43_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_9 XI11_6/XI0/XI0_43/d__9_ xsel_43_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_8 XI11_6/XI0/XI0_43/d__8_ xsel_43_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_7 XI11_6/XI0/XI0_43/d__7_ xsel_43_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_6 XI11_6/XI0/XI0_43/d__6_ xsel_43_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_5 XI11_6/XI0/XI0_43/d__5_ xsel_43_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_4 XI11_6/XI0/XI0_43/d__4_ xsel_43_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_3 XI11_6/XI0/XI0_43/d__3_ xsel_43_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_2 XI11_6/XI0/XI0_43/d__2_ xsel_43_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_1 XI11_6/XI0/XI0_43/d__1_ xsel_43_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_0 XI11_6/XI0/XI0_43/d__0_ xsel_43_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_15 XI11_6/net21_0_ xsel_42_ XI11_6/XI0/XI0_42/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_14 XI11_6/net21_1_ xsel_42_ XI11_6/XI0/XI0_42/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_13 XI11_6/net21_2_ xsel_42_ XI11_6/XI0/XI0_42/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_12 XI11_6/net21_3_ xsel_42_ XI11_6/XI0/XI0_42/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_11 XI11_6/net21_4_ xsel_42_ XI11_6/XI0/XI0_42/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_10 XI11_6/net21_5_ xsel_42_ XI11_6/XI0/XI0_42/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_9 XI11_6/net21_6_ xsel_42_ XI11_6/XI0/XI0_42/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_8 XI11_6/net21_7_ xsel_42_ XI11_6/XI0/XI0_42/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_7 XI11_6/net21_8_ xsel_42_ XI11_6/XI0/XI0_42/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_6 XI11_6/net21_9_ xsel_42_ XI11_6/XI0/XI0_42/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_5 XI11_6/net21_10_ xsel_42_ XI11_6/XI0/XI0_42/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_4 XI11_6/net21_11_ xsel_42_ XI11_6/XI0/XI0_42/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_3 XI11_6/net21_12_ xsel_42_ XI11_6/XI0/XI0_42/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_2 XI11_6/net21_13_ xsel_42_ XI11_6/XI0/XI0_42/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_1 XI11_6/net21_14_ xsel_42_ XI11_6/XI0/XI0_42/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_0 XI11_6/net21_15_ xsel_42_ XI11_6/XI0/XI0_42/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_15 XI11_6/XI0/XI0_42/d__15_ xsel_42_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_14 XI11_6/XI0/XI0_42/d__14_ xsel_42_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_13 XI11_6/XI0/XI0_42/d__13_ xsel_42_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_12 XI11_6/XI0/XI0_42/d__12_ xsel_42_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_11 XI11_6/XI0/XI0_42/d__11_ xsel_42_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_10 XI11_6/XI0/XI0_42/d__10_ xsel_42_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_9 XI11_6/XI0/XI0_42/d__9_ xsel_42_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_8 XI11_6/XI0/XI0_42/d__8_ xsel_42_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_7 XI11_6/XI0/XI0_42/d__7_ xsel_42_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_6 XI11_6/XI0/XI0_42/d__6_ xsel_42_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_5 XI11_6/XI0/XI0_42/d__5_ xsel_42_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_4 XI11_6/XI0/XI0_42/d__4_ xsel_42_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_3 XI11_6/XI0/XI0_42/d__3_ xsel_42_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_2 XI11_6/XI0/XI0_42/d__2_ xsel_42_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_1 XI11_6/XI0/XI0_42/d__1_ xsel_42_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_0 XI11_6/XI0/XI0_42/d__0_ xsel_42_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_15 XI11_6/net21_0_ xsel_41_ XI11_6/XI0/XI0_41/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_14 XI11_6/net21_1_ xsel_41_ XI11_6/XI0/XI0_41/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_13 XI11_6/net21_2_ xsel_41_ XI11_6/XI0/XI0_41/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_12 XI11_6/net21_3_ xsel_41_ XI11_6/XI0/XI0_41/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_11 XI11_6/net21_4_ xsel_41_ XI11_6/XI0/XI0_41/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_10 XI11_6/net21_5_ xsel_41_ XI11_6/XI0/XI0_41/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_9 XI11_6/net21_6_ xsel_41_ XI11_6/XI0/XI0_41/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_8 XI11_6/net21_7_ xsel_41_ XI11_6/XI0/XI0_41/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_7 XI11_6/net21_8_ xsel_41_ XI11_6/XI0/XI0_41/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_6 XI11_6/net21_9_ xsel_41_ XI11_6/XI0/XI0_41/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_5 XI11_6/net21_10_ xsel_41_ XI11_6/XI0/XI0_41/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_4 XI11_6/net21_11_ xsel_41_ XI11_6/XI0/XI0_41/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_3 XI11_6/net21_12_ xsel_41_ XI11_6/XI0/XI0_41/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_2 XI11_6/net21_13_ xsel_41_ XI11_6/XI0/XI0_41/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_1 XI11_6/net21_14_ xsel_41_ XI11_6/XI0/XI0_41/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_0 XI11_6/net21_15_ xsel_41_ XI11_6/XI0/XI0_41/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_15 XI11_6/XI0/XI0_41/d__15_ xsel_41_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_14 XI11_6/XI0/XI0_41/d__14_ xsel_41_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_13 XI11_6/XI0/XI0_41/d__13_ xsel_41_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_12 XI11_6/XI0/XI0_41/d__12_ xsel_41_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_11 XI11_6/XI0/XI0_41/d__11_ xsel_41_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_10 XI11_6/XI0/XI0_41/d__10_ xsel_41_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_9 XI11_6/XI0/XI0_41/d__9_ xsel_41_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_8 XI11_6/XI0/XI0_41/d__8_ xsel_41_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_7 XI11_6/XI0/XI0_41/d__7_ xsel_41_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_6 XI11_6/XI0/XI0_41/d__6_ xsel_41_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_5 XI11_6/XI0/XI0_41/d__5_ xsel_41_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_4 XI11_6/XI0/XI0_41/d__4_ xsel_41_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_3 XI11_6/XI0/XI0_41/d__3_ xsel_41_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_2 XI11_6/XI0/XI0_41/d__2_ xsel_41_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_1 XI11_6/XI0/XI0_41/d__1_ xsel_41_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_0 XI11_6/XI0/XI0_41/d__0_ xsel_41_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_15 XI11_6/net21_0_ xsel_40_ XI11_6/XI0/XI0_40/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_14 XI11_6/net21_1_ xsel_40_ XI11_6/XI0/XI0_40/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_13 XI11_6/net21_2_ xsel_40_ XI11_6/XI0/XI0_40/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_12 XI11_6/net21_3_ xsel_40_ XI11_6/XI0/XI0_40/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_11 XI11_6/net21_4_ xsel_40_ XI11_6/XI0/XI0_40/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_10 XI11_6/net21_5_ xsel_40_ XI11_6/XI0/XI0_40/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_9 XI11_6/net21_6_ xsel_40_ XI11_6/XI0/XI0_40/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_8 XI11_6/net21_7_ xsel_40_ XI11_6/XI0/XI0_40/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_7 XI11_6/net21_8_ xsel_40_ XI11_6/XI0/XI0_40/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_6 XI11_6/net21_9_ xsel_40_ XI11_6/XI0/XI0_40/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_5 XI11_6/net21_10_ xsel_40_ XI11_6/XI0/XI0_40/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_4 XI11_6/net21_11_ xsel_40_ XI11_6/XI0/XI0_40/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_3 XI11_6/net21_12_ xsel_40_ XI11_6/XI0/XI0_40/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_2 XI11_6/net21_13_ xsel_40_ XI11_6/XI0/XI0_40/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_1 XI11_6/net21_14_ xsel_40_ XI11_6/XI0/XI0_40/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_0 XI11_6/net21_15_ xsel_40_ XI11_6/XI0/XI0_40/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_15 XI11_6/XI0/XI0_40/d__15_ xsel_40_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_14 XI11_6/XI0/XI0_40/d__14_ xsel_40_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_13 XI11_6/XI0/XI0_40/d__13_ xsel_40_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_12 XI11_6/XI0/XI0_40/d__12_ xsel_40_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_11 XI11_6/XI0/XI0_40/d__11_ xsel_40_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_10 XI11_6/XI0/XI0_40/d__10_ xsel_40_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_9 XI11_6/XI0/XI0_40/d__9_ xsel_40_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_8 XI11_6/XI0/XI0_40/d__8_ xsel_40_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_7 XI11_6/XI0/XI0_40/d__7_ xsel_40_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_6 XI11_6/XI0/XI0_40/d__6_ xsel_40_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_5 XI11_6/XI0/XI0_40/d__5_ xsel_40_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_4 XI11_6/XI0/XI0_40/d__4_ xsel_40_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_3 XI11_6/XI0/XI0_40/d__3_ xsel_40_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_2 XI11_6/XI0/XI0_40/d__2_ xsel_40_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_1 XI11_6/XI0/XI0_40/d__1_ xsel_40_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_0 XI11_6/XI0/XI0_40/d__0_ xsel_40_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_15 XI11_6/net21_0_ xsel_39_ XI11_6/XI0/XI0_39/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_14 XI11_6/net21_1_ xsel_39_ XI11_6/XI0/XI0_39/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_13 XI11_6/net21_2_ xsel_39_ XI11_6/XI0/XI0_39/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_12 XI11_6/net21_3_ xsel_39_ XI11_6/XI0/XI0_39/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_11 XI11_6/net21_4_ xsel_39_ XI11_6/XI0/XI0_39/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_10 XI11_6/net21_5_ xsel_39_ XI11_6/XI0/XI0_39/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_9 XI11_6/net21_6_ xsel_39_ XI11_6/XI0/XI0_39/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_8 XI11_6/net21_7_ xsel_39_ XI11_6/XI0/XI0_39/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_7 XI11_6/net21_8_ xsel_39_ XI11_6/XI0/XI0_39/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_6 XI11_6/net21_9_ xsel_39_ XI11_6/XI0/XI0_39/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_5 XI11_6/net21_10_ xsel_39_ XI11_6/XI0/XI0_39/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_4 XI11_6/net21_11_ xsel_39_ XI11_6/XI0/XI0_39/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_3 XI11_6/net21_12_ xsel_39_ XI11_6/XI0/XI0_39/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_2 XI11_6/net21_13_ xsel_39_ XI11_6/XI0/XI0_39/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_1 XI11_6/net21_14_ xsel_39_ XI11_6/XI0/XI0_39/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_0 XI11_6/net21_15_ xsel_39_ XI11_6/XI0/XI0_39/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_15 XI11_6/XI0/XI0_39/d__15_ xsel_39_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_14 XI11_6/XI0/XI0_39/d__14_ xsel_39_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_13 XI11_6/XI0/XI0_39/d__13_ xsel_39_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_12 XI11_6/XI0/XI0_39/d__12_ xsel_39_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_11 XI11_6/XI0/XI0_39/d__11_ xsel_39_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_10 XI11_6/XI0/XI0_39/d__10_ xsel_39_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_9 XI11_6/XI0/XI0_39/d__9_ xsel_39_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_8 XI11_6/XI0/XI0_39/d__8_ xsel_39_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_7 XI11_6/XI0/XI0_39/d__7_ xsel_39_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_6 XI11_6/XI0/XI0_39/d__6_ xsel_39_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_5 XI11_6/XI0/XI0_39/d__5_ xsel_39_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_4 XI11_6/XI0/XI0_39/d__4_ xsel_39_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_3 XI11_6/XI0/XI0_39/d__3_ xsel_39_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_2 XI11_6/XI0/XI0_39/d__2_ xsel_39_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_1 XI11_6/XI0/XI0_39/d__1_ xsel_39_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_0 XI11_6/XI0/XI0_39/d__0_ xsel_39_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_15 XI11_6/net21_0_ xsel_38_ XI11_6/XI0/XI0_38/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_14 XI11_6/net21_1_ xsel_38_ XI11_6/XI0/XI0_38/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_13 XI11_6/net21_2_ xsel_38_ XI11_6/XI0/XI0_38/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_12 XI11_6/net21_3_ xsel_38_ XI11_6/XI0/XI0_38/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_11 XI11_6/net21_4_ xsel_38_ XI11_6/XI0/XI0_38/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_10 XI11_6/net21_5_ xsel_38_ XI11_6/XI0/XI0_38/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_9 XI11_6/net21_6_ xsel_38_ XI11_6/XI0/XI0_38/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_8 XI11_6/net21_7_ xsel_38_ XI11_6/XI0/XI0_38/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_7 XI11_6/net21_8_ xsel_38_ XI11_6/XI0/XI0_38/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_6 XI11_6/net21_9_ xsel_38_ XI11_6/XI0/XI0_38/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_5 XI11_6/net21_10_ xsel_38_ XI11_6/XI0/XI0_38/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_4 XI11_6/net21_11_ xsel_38_ XI11_6/XI0/XI0_38/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_3 XI11_6/net21_12_ xsel_38_ XI11_6/XI0/XI0_38/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_2 XI11_6/net21_13_ xsel_38_ XI11_6/XI0/XI0_38/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_1 XI11_6/net21_14_ xsel_38_ XI11_6/XI0/XI0_38/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_0 XI11_6/net21_15_ xsel_38_ XI11_6/XI0/XI0_38/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_15 XI11_6/XI0/XI0_38/d__15_ xsel_38_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_14 XI11_6/XI0/XI0_38/d__14_ xsel_38_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_13 XI11_6/XI0/XI0_38/d__13_ xsel_38_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_12 XI11_6/XI0/XI0_38/d__12_ xsel_38_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_11 XI11_6/XI0/XI0_38/d__11_ xsel_38_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_10 XI11_6/XI0/XI0_38/d__10_ xsel_38_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_9 XI11_6/XI0/XI0_38/d__9_ xsel_38_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_8 XI11_6/XI0/XI0_38/d__8_ xsel_38_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_7 XI11_6/XI0/XI0_38/d__7_ xsel_38_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_6 XI11_6/XI0/XI0_38/d__6_ xsel_38_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_5 XI11_6/XI0/XI0_38/d__5_ xsel_38_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_4 XI11_6/XI0/XI0_38/d__4_ xsel_38_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_3 XI11_6/XI0/XI0_38/d__3_ xsel_38_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_2 XI11_6/XI0/XI0_38/d__2_ xsel_38_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_1 XI11_6/XI0/XI0_38/d__1_ xsel_38_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_0 XI11_6/XI0/XI0_38/d__0_ xsel_38_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_15 XI11_6/net21_0_ xsel_37_ XI11_6/XI0/XI0_37/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_14 XI11_6/net21_1_ xsel_37_ XI11_6/XI0/XI0_37/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_13 XI11_6/net21_2_ xsel_37_ XI11_6/XI0/XI0_37/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_12 XI11_6/net21_3_ xsel_37_ XI11_6/XI0/XI0_37/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_11 XI11_6/net21_4_ xsel_37_ XI11_6/XI0/XI0_37/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_10 XI11_6/net21_5_ xsel_37_ XI11_6/XI0/XI0_37/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_9 XI11_6/net21_6_ xsel_37_ XI11_6/XI0/XI0_37/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_8 XI11_6/net21_7_ xsel_37_ XI11_6/XI0/XI0_37/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_7 XI11_6/net21_8_ xsel_37_ XI11_6/XI0/XI0_37/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_6 XI11_6/net21_9_ xsel_37_ XI11_6/XI0/XI0_37/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_5 XI11_6/net21_10_ xsel_37_ XI11_6/XI0/XI0_37/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_4 XI11_6/net21_11_ xsel_37_ XI11_6/XI0/XI0_37/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_3 XI11_6/net21_12_ xsel_37_ XI11_6/XI0/XI0_37/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_2 XI11_6/net21_13_ xsel_37_ XI11_6/XI0/XI0_37/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_1 XI11_6/net21_14_ xsel_37_ XI11_6/XI0/XI0_37/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_0 XI11_6/net21_15_ xsel_37_ XI11_6/XI0/XI0_37/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_15 XI11_6/XI0/XI0_37/d__15_ xsel_37_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_14 XI11_6/XI0/XI0_37/d__14_ xsel_37_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_13 XI11_6/XI0/XI0_37/d__13_ xsel_37_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_12 XI11_6/XI0/XI0_37/d__12_ xsel_37_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_11 XI11_6/XI0/XI0_37/d__11_ xsel_37_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_10 XI11_6/XI0/XI0_37/d__10_ xsel_37_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_9 XI11_6/XI0/XI0_37/d__9_ xsel_37_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_8 XI11_6/XI0/XI0_37/d__8_ xsel_37_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_7 XI11_6/XI0/XI0_37/d__7_ xsel_37_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_6 XI11_6/XI0/XI0_37/d__6_ xsel_37_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_5 XI11_6/XI0/XI0_37/d__5_ xsel_37_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_4 XI11_6/XI0/XI0_37/d__4_ xsel_37_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_3 XI11_6/XI0/XI0_37/d__3_ xsel_37_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_2 XI11_6/XI0/XI0_37/d__2_ xsel_37_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_1 XI11_6/XI0/XI0_37/d__1_ xsel_37_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_0 XI11_6/XI0/XI0_37/d__0_ xsel_37_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_15 XI11_6/net21_0_ xsel_36_ XI11_6/XI0/XI0_36/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_14 XI11_6/net21_1_ xsel_36_ XI11_6/XI0/XI0_36/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_13 XI11_6/net21_2_ xsel_36_ XI11_6/XI0/XI0_36/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_12 XI11_6/net21_3_ xsel_36_ XI11_6/XI0/XI0_36/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_11 XI11_6/net21_4_ xsel_36_ XI11_6/XI0/XI0_36/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_10 XI11_6/net21_5_ xsel_36_ XI11_6/XI0/XI0_36/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_9 XI11_6/net21_6_ xsel_36_ XI11_6/XI0/XI0_36/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_8 XI11_6/net21_7_ xsel_36_ XI11_6/XI0/XI0_36/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_7 XI11_6/net21_8_ xsel_36_ XI11_6/XI0/XI0_36/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_6 XI11_6/net21_9_ xsel_36_ XI11_6/XI0/XI0_36/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_5 XI11_6/net21_10_ xsel_36_ XI11_6/XI0/XI0_36/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_4 XI11_6/net21_11_ xsel_36_ XI11_6/XI0/XI0_36/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_3 XI11_6/net21_12_ xsel_36_ XI11_6/XI0/XI0_36/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_2 XI11_6/net21_13_ xsel_36_ XI11_6/XI0/XI0_36/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_1 XI11_6/net21_14_ xsel_36_ XI11_6/XI0/XI0_36/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_0 XI11_6/net21_15_ xsel_36_ XI11_6/XI0/XI0_36/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_15 XI11_6/XI0/XI0_36/d__15_ xsel_36_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_14 XI11_6/XI0/XI0_36/d__14_ xsel_36_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_13 XI11_6/XI0/XI0_36/d__13_ xsel_36_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_12 XI11_6/XI0/XI0_36/d__12_ xsel_36_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_11 XI11_6/XI0/XI0_36/d__11_ xsel_36_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_10 XI11_6/XI0/XI0_36/d__10_ xsel_36_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_9 XI11_6/XI0/XI0_36/d__9_ xsel_36_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_8 XI11_6/XI0/XI0_36/d__8_ xsel_36_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_7 XI11_6/XI0/XI0_36/d__7_ xsel_36_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_6 XI11_6/XI0/XI0_36/d__6_ xsel_36_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_5 XI11_6/XI0/XI0_36/d__5_ xsel_36_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_4 XI11_6/XI0/XI0_36/d__4_ xsel_36_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_3 XI11_6/XI0/XI0_36/d__3_ xsel_36_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_2 XI11_6/XI0/XI0_36/d__2_ xsel_36_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_1 XI11_6/XI0/XI0_36/d__1_ xsel_36_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_0 XI11_6/XI0/XI0_36/d__0_ xsel_36_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_15 XI11_6/net21_0_ xsel_35_ XI11_6/XI0/XI0_35/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_14 XI11_6/net21_1_ xsel_35_ XI11_6/XI0/XI0_35/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_13 XI11_6/net21_2_ xsel_35_ XI11_6/XI0/XI0_35/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_12 XI11_6/net21_3_ xsel_35_ XI11_6/XI0/XI0_35/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_11 XI11_6/net21_4_ xsel_35_ XI11_6/XI0/XI0_35/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_10 XI11_6/net21_5_ xsel_35_ XI11_6/XI0/XI0_35/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_9 XI11_6/net21_6_ xsel_35_ XI11_6/XI0/XI0_35/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_8 XI11_6/net21_7_ xsel_35_ XI11_6/XI0/XI0_35/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_7 XI11_6/net21_8_ xsel_35_ XI11_6/XI0/XI0_35/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_6 XI11_6/net21_9_ xsel_35_ XI11_6/XI0/XI0_35/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_5 XI11_6/net21_10_ xsel_35_ XI11_6/XI0/XI0_35/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_4 XI11_6/net21_11_ xsel_35_ XI11_6/XI0/XI0_35/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_3 XI11_6/net21_12_ xsel_35_ XI11_6/XI0/XI0_35/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_2 XI11_6/net21_13_ xsel_35_ XI11_6/XI0/XI0_35/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_1 XI11_6/net21_14_ xsel_35_ XI11_6/XI0/XI0_35/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_0 XI11_6/net21_15_ xsel_35_ XI11_6/XI0/XI0_35/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_15 XI11_6/XI0/XI0_35/d__15_ xsel_35_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_14 XI11_6/XI0/XI0_35/d__14_ xsel_35_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_13 XI11_6/XI0/XI0_35/d__13_ xsel_35_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_12 XI11_6/XI0/XI0_35/d__12_ xsel_35_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_11 XI11_6/XI0/XI0_35/d__11_ xsel_35_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_10 XI11_6/XI0/XI0_35/d__10_ xsel_35_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_9 XI11_6/XI0/XI0_35/d__9_ xsel_35_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_8 XI11_6/XI0/XI0_35/d__8_ xsel_35_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_7 XI11_6/XI0/XI0_35/d__7_ xsel_35_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_6 XI11_6/XI0/XI0_35/d__6_ xsel_35_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_5 XI11_6/XI0/XI0_35/d__5_ xsel_35_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_4 XI11_6/XI0/XI0_35/d__4_ xsel_35_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_3 XI11_6/XI0/XI0_35/d__3_ xsel_35_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_2 XI11_6/XI0/XI0_35/d__2_ xsel_35_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_1 XI11_6/XI0/XI0_35/d__1_ xsel_35_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_0 XI11_6/XI0/XI0_35/d__0_ xsel_35_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_15 XI11_6/net21_0_ xsel_34_ XI11_6/XI0/XI0_34/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_14 XI11_6/net21_1_ xsel_34_ XI11_6/XI0/XI0_34/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_13 XI11_6/net21_2_ xsel_34_ XI11_6/XI0/XI0_34/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_12 XI11_6/net21_3_ xsel_34_ XI11_6/XI0/XI0_34/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_11 XI11_6/net21_4_ xsel_34_ XI11_6/XI0/XI0_34/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_10 XI11_6/net21_5_ xsel_34_ XI11_6/XI0/XI0_34/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_9 XI11_6/net21_6_ xsel_34_ XI11_6/XI0/XI0_34/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_8 XI11_6/net21_7_ xsel_34_ XI11_6/XI0/XI0_34/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_7 XI11_6/net21_8_ xsel_34_ XI11_6/XI0/XI0_34/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_6 XI11_6/net21_9_ xsel_34_ XI11_6/XI0/XI0_34/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_5 XI11_6/net21_10_ xsel_34_ XI11_6/XI0/XI0_34/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_4 XI11_6/net21_11_ xsel_34_ XI11_6/XI0/XI0_34/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_3 XI11_6/net21_12_ xsel_34_ XI11_6/XI0/XI0_34/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_2 XI11_6/net21_13_ xsel_34_ XI11_6/XI0/XI0_34/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_1 XI11_6/net21_14_ xsel_34_ XI11_6/XI0/XI0_34/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_0 XI11_6/net21_15_ xsel_34_ XI11_6/XI0/XI0_34/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_15 XI11_6/XI0/XI0_34/d__15_ xsel_34_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_14 XI11_6/XI0/XI0_34/d__14_ xsel_34_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_13 XI11_6/XI0/XI0_34/d__13_ xsel_34_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_12 XI11_6/XI0/XI0_34/d__12_ xsel_34_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_11 XI11_6/XI0/XI0_34/d__11_ xsel_34_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_10 XI11_6/XI0/XI0_34/d__10_ xsel_34_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_9 XI11_6/XI0/XI0_34/d__9_ xsel_34_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_8 XI11_6/XI0/XI0_34/d__8_ xsel_34_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_7 XI11_6/XI0/XI0_34/d__7_ xsel_34_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_6 XI11_6/XI0/XI0_34/d__6_ xsel_34_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_5 XI11_6/XI0/XI0_34/d__5_ xsel_34_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_4 XI11_6/XI0/XI0_34/d__4_ xsel_34_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_3 XI11_6/XI0/XI0_34/d__3_ xsel_34_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_2 XI11_6/XI0/XI0_34/d__2_ xsel_34_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_1 XI11_6/XI0/XI0_34/d__1_ xsel_34_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_0 XI11_6/XI0/XI0_34/d__0_ xsel_34_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_15 XI11_6/net21_0_ xsel_33_ XI11_6/XI0/XI0_33/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_14 XI11_6/net21_1_ xsel_33_ XI11_6/XI0/XI0_33/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_13 XI11_6/net21_2_ xsel_33_ XI11_6/XI0/XI0_33/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_12 XI11_6/net21_3_ xsel_33_ XI11_6/XI0/XI0_33/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_11 XI11_6/net21_4_ xsel_33_ XI11_6/XI0/XI0_33/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_10 XI11_6/net21_5_ xsel_33_ XI11_6/XI0/XI0_33/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_9 XI11_6/net21_6_ xsel_33_ XI11_6/XI0/XI0_33/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_8 XI11_6/net21_7_ xsel_33_ XI11_6/XI0/XI0_33/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_7 XI11_6/net21_8_ xsel_33_ XI11_6/XI0/XI0_33/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_6 XI11_6/net21_9_ xsel_33_ XI11_6/XI0/XI0_33/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_5 XI11_6/net21_10_ xsel_33_ XI11_6/XI0/XI0_33/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_4 XI11_6/net21_11_ xsel_33_ XI11_6/XI0/XI0_33/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_3 XI11_6/net21_12_ xsel_33_ XI11_6/XI0/XI0_33/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_2 XI11_6/net21_13_ xsel_33_ XI11_6/XI0/XI0_33/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_1 XI11_6/net21_14_ xsel_33_ XI11_6/XI0/XI0_33/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_0 XI11_6/net21_15_ xsel_33_ XI11_6/XI0/XI0_33/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_15 XI11_6/XI0/XI0_33/d__15_ xsel_33_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_14 XI11_6/XI0/XI0_33/d__14_ xsel_33_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_13 XI11_6/XI0/XI0_33/d__13_ xsel_33_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_12 XI11_6/XI0/XI0_33/d__12_ xsel_33_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_11 XI11_6/XI0/XI0_33/d__11_ xsel_33_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_10 XI11_6/XI0/XI0_33/d__10_ xsel_33_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_9 XI11_6/XI0/XI0_33/d__9_ xsel_33_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_8 XI11_6/XI0/XI0_33/d__8_ xsel_33_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_7 XI11_6/XI0/XI0_33/d__7_ xsel_33_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_6 XI11_6/XI0/XI0_33/d__6_ xsel_33_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_5 XI11_6/XI0/XI0_33/d__5_ xsel_33_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_4 XI11_6/XI0/XI0_33/d__4_ xsel_33_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_3 XI11_6/XI0/XI0_33/d__3_ xsel_33_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_2 XI11_6/XI0/XI0_33/d__2_ xsel_33_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_1 XI11_6/XI0/XI0_33/d__1_ xsel_33_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_0 XI11_6/XI0/XI0_33/d__0_ xsel_33_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_15 XI11_6/net21_0_ xsel_32_ XI11_6/XI0/XI0_32/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_14 XI11_6/net21_1_ xsel_32_ XI11_6/XI0/XI0_32/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_13 XI11_6/net21_2_ xsel_32_ XI11_6/XI0/XI0_32/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_12 XI11_6/net21_3_ xsel_32_ XI11_6/XI0/XI0_32/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_11 XI11_6/net21_4_ xsel_32_ XI11_6/XI0/XI0_32/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_10 XI11_6/net21_5_ xsel_32_ XI11_6/XI0/XI0_32/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_9 XI11_6/net21_6_ xsel_32_ XI11_6/XI0/XI0_32/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_8 XI11_6/net21_7_ xsel_32_ XI11_6/XI0/XI0_32/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_7 XI11_6/net21_8_ xsel_32_ XI11_6/XI0/XI0_32/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_6 XI11_6/net21_9_ xsel_32_ XI11_6/XI0/XI0_32/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_5 XI11_6/net21_10_ xsel_32_ XI11_6/XI0/XI0_32/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_4 XI11_6/net21_11_ xsel_32_ XI11_6/XI0/XI0_32/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_3 XI11_6/net21_12_ xsel_32_ XI11_6/XI0/XI0_32/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_2 XI11_6/net21_13_ xsel_32_ XI11_6/XI0/XI0_32/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_1 XI11_6/net21_14_ xsel_32_ XI11_6/XI0/XI0_32/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_0 XI11_6/net21_15_ xsel_32_ XI11_6/XI0/XI0_32/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_15 XI11_6/XI0/XI0_32/d__15_ xsel_32_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_14 XI11_6/XI0/XI0_32/d__14_ xsel_32_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_13 XI11_6/XI0/XI0_32/d__13_ xsel_32_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_12 XI11_6/XI0/XI0_32/d__12_ xsel_32_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_11 XI11_6/XI0/XI0_32/d__11_ xsel_32_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_10 XI11_6/XI0/XI0_32/d__10_ xsel_32_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_9 XI11_6/XI0/XI0_32/d__9_ xsel_32_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_8 XI11_6/XI0/XI0_32/d__8_ xsel_32_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_7 XI11_6/XI0/XI0_32/d__7_ xsel_32_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_6 XI11_6/XI0/XI0_32/d__6_ xsel_32_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_5 XI11_6/XI0/XI0_32/d__5_ xsel_32_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_4 XI11_6/XI0/XI0_32/d__4_ xsel_32_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_3 XI11_6/XI0/XI0_32/d__3_ xsel_32_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_2 XI11_6/XI0/XI0_32/d__2_ xsel_32_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_1 XI11_6/XI0/XI0_32/d__1_ xsel_32_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_0 XI11_6/XI0/XI0_32/d__0_ xsel_32_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_15 XI11_6/net21_0_ xsel_31_ XI11_6/XI0/XI0_31/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_14 XI11_6/net21_1_ xsel_31_ XI11_6/XI0/XI0_31/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_13 XI11_6/net21_2_ xsel_31_ XI11_6/XI0/XI0_31/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_12 XI11_6/net21_3_ xsel_31_ XI11_6/XI0/XI0_31/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_11 XI11_6/net21_4_ xsel_31_ XI11_6/XI0/XI0_31/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_10 XI11_6/net21_5_ xsel_31_ XI11_6/XI0/XI0_31/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_9 XI11_6/net21_6_ xsel_31_ XI11_6/XI0/XI0_31/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_8 XI11_6/net21_7_ xsel_31_ XI11_6/XI0/XI0_31/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_7 XI11_6/net21_8_ xsel_31_ XI11_6/XI0/XI0_31/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_6 XI11_6/net21_9_ xsel_31_ XI11_6/XI0/XI0_31/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_5 XI11_6/net21_10_ xsel_31_ XI11_6/XI0/XI0_31/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_4 XI11_6/net21_11_ xsel_31_ XI11_6/XI0/XI0_31/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_3 XI11_6/net21_12_ xsel_31_ XI11_6/XI0/XI0_31/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_2 XI11_6/net21_13_ xsel_31_ XI11_6/XI0/XI0_31/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_1 XI11_6/net21_14_ xsel_31_ XI11_6/XI0/XI0_31/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_0 XI11_6/net21_15_ xsel_31_ XI11_6/XI0/XI0_31/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_15 XI11_6/XI0/XI0_31/d__15_ xsel_31_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_14 XI11_6/XI0/XI0_31/d__14_ xsel_31_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_13 XI11_6/XI0/XI0_31/d__13_ xsel_31_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_12 XI11_6/XI0/XI0_31/d__12_ xsel_31_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_11 XI11_6/XI0/XI0_31/d__11_ xsel_31_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_10 XI11_6/XI0/XI0_31/d__10_ xsel_31_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_9 XI11_6/XI0/XI0_31/d__9_ xsel_31_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_8 XI11_6/XI0/XI0_31/d__8_ xsel_31_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_7 XI11_6/XI0/XI0_31/d__7_ xsel_31_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_6 XI11_6/XI0/XI0_31/d__6_ xsel_31_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_5 XI11_6/XI0/XI0_31/d__5_ xsel_31_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_4 XI11_6/XI0/XI0_31/d__4_ xsel_31_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_3 XI11_6/XI0/XI0_31/d__3_ xsel_31_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_2 XI11_6/XI0/XI0_31/d__2_ xsel_31_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_1 XI11_6/XI0/XI0_31/d__1_ xsel_31_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_0 XI11_6/XI0/XI0_31/d__0_ xsel_31_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_15 XI11_6/net21_0_ xsel_30_ XI11_6/XI0/XI0_30/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_14 XI11_6/net21_1_ xsel_30_ XI11_6/XI0/XI0_30/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_13 XI11_6/net21_2_ xsel_30_ XI11_6/XI0/XI0_30/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_12 XI11_6/net21_3_ xsel_30_ XI11_6/XI0/XI0_30/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_11 XI11_6/net21_4_ xsel_30_ XI11_6/XI0/XI0_30/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_10 XI11_6/net21_5_ xsel_30_ XI11_6/XI0/XI0_30/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_9 XI11_6/net21_6_ xsel_30_ XI11_6/XI0/XI0_30/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_8 XI11_6/net21_7_ xsel_30_ XI11_6/XI0/XI0_30/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_7 XI11_6/net21_8_ xsel_30_ XI11_6/XI0/XI0_30/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_6 XI11_6/net21_9_ xsel_30_ XI11_6/XI0/XI0_30/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_5 XI11_6/net21_10_ xsel_30_ XI11_6/XI0/XI0_30/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_4 XI11_6/net21_11_ xsel_30_ XI11_6/XI0/XI0_30/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_3 XI11_6/net21_12_ xsel_30_ XI11_6/XI0/XI0_30/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_2 XI11_6/net21_13_ xsel_30_ XI11_6/XI0/XI0_30/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_1 XI11_6/net21_14_ xsel_30_ XI11_6/XI0/XI0_30/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_0 XI11_6/net21_15_ xsel_30_ XI11_6/XI0/XI0_30/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_15 XI11_6/XI0/XI0_30/d__15_ xsel_30_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_14 XI11_6/XI0/XI0_30/d__14_ xsel_30_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_13 XI11_6/XI0/XI0_30/d__13_ xsel_30_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_12 XI11_6/XI0/XI0_30/d__12_ xsel_30_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_11 XI11_6/XI0/XI0_30/d__11_ xsel_30_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_10 XI11_6/XI0/XI0_30/d__10_ xsel_30_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_9 XI11_6/XI0/XI0_30/d__9_ xsel_30_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_8 XI11_6/XI0/XI0_30/d__8_ xsel_30_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_7 XI11_6/XI0/XI0_30/d__7_ xsel_30_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_6 XI11_6/XI0/XI0_30/d__6_ xsel_30_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_5 XI11_6/XI0/XI0_30/d__5_ xsel_30_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_4 XI11_6/XI0/XI0_30/d__4_ xsel_30_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_3 XI11_6/XI0/XI0_30/d__3_ xsel_30_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_2 XI11_6/XI0/XI0_30/d__2_ xsel_30_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_1 XI11_6/XI0/XI0_30/d__1_ xsel_30_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_0 XI11_6/XI0/XI0_30/d__0_ xsel_30_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_15 XI11_6/net21_0_ xsel_29_ XI11_6/XI0/XI0_29/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_14 XI11_6/net21_1_ xsel_29_ XI11_6/XI0/XI0_29/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_13 XI11_6/net21_2_ xsel_29_ XI11_6/XI0/XI0_29/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_12 XI11_6/net21_3_ xsel_29_ XI11_6/XI0/XI0_29/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_11 XI11_6/net21_4_ xsel_29_ XI11_6/XI0/XI0_29/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_10 XI11_6/net21_5_ xsel_29_ XI11_6/XI0/XI0_29/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_9 XI11_6/net21_6_ xsel_29_ XI11_6/XI0/XI0_29/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_8 XI11_6/net21_7_ xsel_29_ XI11_6/XI0/XI0_29/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_7 XI11_6/net21_8_ xsel_29_ XI11_6/XI0/XI0_29/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_6 XI11_6/net21_9_ xsel_29_ XI11_6/XI0/XI0_29/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_5 XI11_6/net21_10_ xsel_29_ XI11_6/XI0/XI0_29/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_4 XI11_6/net21_11_ xsel_29_ XI11_6/XI0/XI0_29/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_3 XI11_6/net21_12_ xsel_29_ XI11_6/XI0/XI0_29/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_2 XI11_6/net21_13_ xsel_29_ XI11_6/XI0/XI0_29/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_1 XI11_6/net21_14_ xsel_29_ XI11_6/XI0/XI0_29/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_0 XI11_6/net21_15_ xsel_29_ XI11_6/XI0/XI0_29/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_15 XI11_6/XI0/XI0_29/d__15_ xsel_29_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_14 XI11_6/XI0/XI0_29/d__14_ xsel_29_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_13 XI11_6/XI0/XI0_29/d__13_ xsel_29_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_12 XI11_6/XI0/XI0_29/d__12_ xsel_29_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_11 XI11_6/XI0/XI0_29/d__11_ xsel_29_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_10 XI11_6/XI0/XI0_29/d__10_ xsel_29_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_9 XI11_6/XI0/XI0_29/d__9_ xsel_29_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_8 XI11_6/XI0/XI0_29/d__8_ xsel_29_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_7 XI11_6/XI0/XI0_29/d__7_ xsel_29_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_6 XI11_6/XI0/XI0_29/d__6_ xsel_29_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_5 XI11_6/XI0/XI0_29/d__5_ xsel_29_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_4 XI11_6/XI0/XI0_29/d__4_ xsel_29_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_3 XI11_6/XI0/XI0_29/d__3_ xsel_29_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_2 XI11_6/XI0/XI0_29/d__2_ xsel_29_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_1 XI11_6/XI0/XI0_29/d__1_ xsel_29_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_0 XI11_6/XI0/XI0_29/d__0_ xsel_29_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_15 XI11_6/net21_0_ xsel_28_ XI11_6/XI0/XI0_28/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_14 XI11_6/net21_1_ xsel_28_ XI11_6/XI0/XI0_28/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_13 XI11_6/net21_2_ xsel_28_ XI11_6/XI0/XI0_28/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_12 XI11_6/net21_3_ xsel_28_ XI11_6/XI0/XI0_28/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_11 XI11_6/net21_4_ xsel_28_ XI11_6/XI0/XI0_28/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_10 XI11_6/net21_5_ xsel_28_ XI11_6/XI0/XI0_28/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_9 XI11_6/net21_6_ xsel_28_ XI11_6/XI0/XI0_28/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_8 XI11_6/net21_7_ xsel_28_ XI11_6/XI0/XI0_28/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_7 XI11_6/net21_8_ xsel_28_ XI11_6/XI0/XI0_28/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_6 XI11_6/net21_9_ xsel_28_ XI11_6/XI0/XI0_28/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_5 XI11_6/net21_10_ xsel_28_ XI11_6/XI0/XI0_28/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_4 XI11_6/net21_11_ xsel_28_ XI11_6/XI0/XI0_28/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_3 XI11_6/net21_12_ xsel_28_ XI11_6/XI0/XI0_28/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_2 XI11_6/net21_13_ xsel_28_ XI11_6/XI0/XI0_28/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_1 XI11_6/net21_14_ xsel_28_ XI11_6/XI0/XI0_28/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_0 XI11_6/net21_15_ xsel_28_ XI11_6/XI0/XI0_28/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_15 XI11_6/XI0/XI0_28/d__15_ xsel_28_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_14 XI11_6/XI0/XI0_28/d__14_ xsel_28_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_13 XI11_6/XI0/XI0_28/d__13_ xsel_28_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_12 XI11_6/XI0/XI0_28/d__12_ xsel_28_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_11 XI11_6/XI0/XI0_28/d__11_ xsel_28_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_10 XI11_6/XI0/XI0_28/d__10_ xsel_28_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_9 XI11_6/XI0/XI0_28/d__9_ xsel_28_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_8 XI11_6/XI0/XI0_28/d__8_ xsel_28_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_7 XI11_6/XI0/XI0_28/d__7_ xsel_28_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_6 XI11_6/XI0/XI0_28/d__6_ xsel_28_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_5 XI11_6/XI0/XI0_28/d__5_ xsel_28_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_4 XI11_6/XI0/XI0_28/d__4_ xsel_28_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_3 XI11_6/XI0/XI0_28/d__3_ xsel_28_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_2 XI11_6/XI0/XI0_28/d__2_ xsel_28_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_1 XI11_6/XI0/XI0_28/d__1_ xsel_28_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_0 XI11_6/XI0/XI0_28/d__0_ xsel_28_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_15 XI11_6/net21_0_ xsel_27_ XI11_6/XI0/XI0_27/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_14 XI11_6/net21_1_ xsel_27_ XI11_6/XI0/XI0_27/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_13 XI11_6/net21_2_ xsel_27_ XI11_6/XI0/XI0_27/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_12 XI11_6/net21_3_ xsel_27_ XI11_6/XI0/XI0_27/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_11 XI11_6/net21_4_ xsel_27_ XI11_6/XI0/XI0_27/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_10 XI11_6/net21_5_ xsel_27_ XI11_6/XI0/XI0_27/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_9 XI11_6/net21_6_ xsel_27_ XI11_6/XI0/XI0_27/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_8 XI11_6/net21_7_ xsel_27_ XI11_6/XI0/XI0_27/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_7 XI11_6/net21_8_ xsel_27_ XI11_6/XI0/XI0_27/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_6 XI11_6/net21_9_ xsel_27_ XI11_6/XI0/XI0_27/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_5 XI11_6/net21_10_ xsel_27_ XI11_6/XI0/XI0_27/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_4 XI11_6/net21_11_ xsel_27_ XI11_6/XI0/XI0_27/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_3 XI11_6/net21_12_ xsel_27_ XI11_6/XI0/XI0_27/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_2 XI11_6/net21_13_ xsel_27_ XI11_6/XI0/XI0_27/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_1 XI11_6/net21_14_ xsel_27_ XI11_6/XI0/XI0_27/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_0 XI11_6/net21_15_ xsel_27_ XI11_6/XI0/XI0_27/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_15 XI11_6/XI0/XI0_27/d__15_ xsel_27_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_14 XI11_6/XI0/XI0_27/d__14_ xsel_27_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_13 XI11_6/XI0/XI0_27/d__13_ xsel_27_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_12 XI11_6/XI0/XI0_27/d__12_ xsel_27_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_11 XI11_6/XI0/XI0_27/d__11_ xsel_27_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_10 XI11_6/XI0/XI0_27/d__10_ xsel_27_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_9 XI11_6/XI0/XI0_27/d__9_ xsel_27_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_8 XI11_6/XI0/XI0_27/d__8_ xsel_27_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_7 XI11_6/XI0/XI0_27/d__7_ xsel_27_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_6 XI11_6/XI0/XI0_27/d__6_ xsel_27_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_5 XI11_6/XI0/XI0_27/d__5_ xsel_27_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_4 XI11_6/XI0/XI0_27/d__4_ xsel_27_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_3 XI11_6/XI0/XI0_27/d__3_ xsel_27_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_2 XI11_6/XI0/XI0_27/d__2_ xsel_27_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_1 XI11_6/XI0/XI0_27/d__1_ xsel_27_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_0 XI11_6/XI0/XI0_27/d__0_ xsel_27_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_15 XI11_6/net21_0_ xsel_26_ XI11_6/XI0/XI0_26/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_14 XI11_6/net21_1_ xsel_26_ XI11_6/XI0/XI0_26/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_13 XI11_6/net21_2_ xsel_26_ XI11_6/XI0/XI0_26/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_12 XI11_6/net21_3_ xsel_26_ XI11_6/XI0/XI0_26/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_11 XI11_6/net21_4_ xsel_26_ XI11_6/XI0/XI0_26/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_10 XI11_6/net21_5_ xsel_26_ XI11_6/XI0/XI0_26/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_9 XI11_6/net21_6_ xsel_26_ XI11_6/XI0/XI0_26/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_8 XI11_6/net21_7_ xsel_26_ XI11_6/XI0/XI0_26/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_7 XI11_6/net21_8_ xsel_26_ XI11_6/XI0/XI0_26/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_6 XI11_6/net21_9_ xsel_26_ XI11_6/XI0/XI0_26/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_5 XI11_6/net21_10_ xsel_26_ XI11_6/XI0/XI0_26/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_4 XI11_6/net21_11_ xsel_26_ XI11_6/XI0/XI0_26/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_3 XI11_6/net21_12_ xsel_26_ XI11_6/XI0/XI0_26/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_2 XI11_6/net21_13_ xsel_26_ XI11_6/XI0/XI0_26/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_1 XI11_6/net21_14_ xsel_26_ XI11_6/XI0/XI0_26/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_0 XI11_6/net21_15_ xsel_26_ XI11_6/XI0/XI0_26/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_15 XI11_6/XI0/XI0_26/d__15_ xsel_26_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_14 XI11_6/XI0/XI0_26/d__14_ xsel_26_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_13 XI11_6/XI0/XI0_26/d__13_ xsel_26_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_12 XI11_6/XI0/XI0_26/d__12_ xsel_26_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_11 XI11_6/XI0/XI0_26/d__11_ xsel_26_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_10 XI11_6/XI0/XI0_26/d__10_ xsel_26_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_9 XI11_6/XI0/XI0_26/d__9_ xsel_26_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_8 XI11_6/XI0/XI0_26/d__8_ xsel_26_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_7 XI11_6/XI0/XI0_26/d__7_ xsel_26_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_6 XI11_6/XI0/XI0_26/d__6_ xsel_26_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_5 XI11_6/XI0/XI0_26/d__5_ xsel_26_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_4 XI11_6/XI0/XI0_26/d__4_ xsel_26_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_3 XI11_6/XI0/XI0_26/d__3_ xsel_26_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_2 XI11_6/XI0/XI0_26/d__2_ xsel_26_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_1 XI11_6/XI0/XI0_26/d__1_ xsel_26_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_0 XI11_6/XI0/XI0_26/d__0_ xsel_26_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_15 XI11_6/net21_0_ xsel_25_ XI11_6/XI0/XI0_25/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_14 XI11_6/net21_1_ xsel_25_ XI11_6/XI0/XI0_25/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_13 XI11_6/net21_2_ xsel_25_ XI11_6/XI0/XI0_25/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_12 XI11_6/net21_3_ xsel_25_ XI11_6/XI0/XI0_25/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_11 XI11_6/net21_4_ xsel_25_ XI11_6/XI0/XI0_25/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_10 XI11_6/net21_5_ xsel_25_ XI11_6/XI0/XI0_25/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_9 XI11_6/net21_6_ xsel_25_ XI11_6/XI0/XI0_25/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_8 XI11_6/net21_7_ xsel_25_ XI11_6/XI0/XI0_25/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_7 XI11_6/net21_8_ xsel_25_ XI11_6/XI0/XI0_25/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_6 XI11_6/net21_9_ xsel_25_ XI11_6/XI0/XI0_25/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_5 XI11_6/net21_10_ xsel_25_ XI11_6/XI0/XI0_25/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_4 XI11_6/net21_11_ xsel_25_ XI11_6/XI0/XI0_25/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_3 XI11_6/net21_12_ xsel_25_ XI11_6/XI0/XI0_25/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_2 XI11_6/net21_13_ xsel_25_ XI11_6/XI0/XI0_25/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_1 XI11_6/net21_14_ xsel_25_ XI11_6/XI0/XI0_25/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_0 XI11_6/net21_15_ xsel_25_ XI11_6/XI0/XI0_25/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_15 XI11_6/XI0/XI0_25/d__15_ xsel_25_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_14 XI11_6/XI0/XI0_25/d__14_ xsel_25_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_13 XI11_6/XI0/XI0_25/d__13_ xsel_25_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_12 XI11_6/XI0/XI0_25/d__12_ xsel_25_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_11 XI11_6/XI0/XI0_25/d__11_ xsel_25_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_10 XI11_6/XI0/XI0_25/d__10_ xsel_25_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_9 XI11_6/XI0/XI0_25/d__9_ xsel_25_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_8 XI11_6/XI0/XI0_25/d__8_ xsel_25_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_7 XI11_6/XI0/XI0_25/d__7_ xsel_25_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_6 XI11_6/XI0/XI0_25/d__6_ xsel_25_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_5 XI11_6/XI0/XI0_25/d__5_ xsel_25_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_4 XI11_6/XI0/XI0_25/d__4_ xsel_25_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_3 XI11_6/XI0/XI0_25/d__3_ xsel_25_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_2 XI11_6/XI0/XI0_25/d__2_ xsel_25_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_1 XI11_6/XI0/XI0_25/d__1_ xsel_25_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_0 XI11_6/XI0/XI0_25/d__0_ xsel_25_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_15 XI11_6/net21_0_ xsel_24_ XI11_6/XI0/XI0_24/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_14 XI11_6/net21_1_ xsel_24_ XI11_6/XI0/XI0_24/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_13 XI11_6/net21_2_ xsel_24_ XI11_6/XI0/XI0_24/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_12 XI11_6/net21_3_ xsel_24_ XI11_6/XI0/XI0_24/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_11 XI11_6/net21_4_ xsel_24_ XI11_6/XI0/XI0_24/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_10 XI11_6/net21_5_ xsel_24_ XI11_6/XI0/XI0_24/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_9 XI11_6/net21_6_ xsel_24_ XI11_6/XI0/XI0_24/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_8 XI11_6/net21_7_ xsel_24_ XI11_6/XI0/XI0_24/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_7 XI11_6/net21_8_ xsel_24_ XI11_6/XI0/XI0_24/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_6 XI11_6/net21_9_ xsel_24_ XI11_6/XI0/XI0_24/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_5 XI11_6/net21_10_ xsel_24_ XI11_6/XI0/XI0_24/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_4 XI11_6/net21_11_ xsel_24_ XI11_6/XI0/XI0_24/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_3 XI11_6/net21_12_ xsel_24_ XI11_6/XI0/XI0_24/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_2 XI11_6/net21_13_ xsel_24_ XI11_6/XI0/XI0_24/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_1 XI11_6/net21_14_ xsel_24_ XI11_6/XI0/XI0_24/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_0 XI11_6/net21_15_ xsel_24_ XI11_6/XI0/XI0_24/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_15 XI11_6/XI0/XI0_24/d__15_ xsel_24_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_14 XI11_6/XI0/XI0_24/d__14_ xsel_24_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_13 XI11_6/XI0/XI0_24/d__13_ xsel_24_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_12 XI11_6/XI0/XI0_24/d__12_ xsel_24_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_11 XI11_6/XI0/XI0_24/d__11_ xsel_24_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_10 XI11_6/XI0/XI0_24/d__10_ xsel_24_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_9 XI11_6/XI0/XI0_24/d__9_ xsel_24_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_8 XI11_6/XI0/XI0_24/d__8_ xsel_24_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_7 XI11_6/XI0/XI0_24/d__7_ xsel_24_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_6 XI11_6/XI0/XI0_24/d__6_ xsel_24_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_5 XI11_6/XI0/XI0_24/d__5_ xsel_24_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_4 XI11_6/XI0/XI0_24/d__4_ xsel_24_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_3 XI11_6/XI0/XI0_24/d__3_ xsel_24_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_2 XI11_6/XI0/XI0_24/d__2_ xsel_24_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_1 XI11_6/XI0/XI0_24/d__1_ xsel_24_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_0 XI11_6/XI0/XI0_24/d__0_ xsel_24_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_15 XI11_6/net21_0_ xsel_23_ XI11_6/XI0/XI0_23/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_14 XI11_6/net21_1_ xsel_23_ XI11_6/XI0/XI0_23/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_13 XI11_6/net21_2_ xsel_23_ XI11_6/XI0/XI0_23/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_12 XI11_6/net21_3_ xsel_23_ XI11_6/XI0/XI0_23/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_11 XI11_6/net21_4_ xsel_23_ XI11_6/XI0/XI0_23/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_10 XI11_6/net21_5_ xsel_23_ XI11_6/XI0/XI0_23/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_9 XI11_6/net21_6_ xsel_23_ XI11_6/XI0/XI0_23/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_8 XI11_6/net21_7_ xsel_23_ XI11_6/XI0/XI0_23/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_7 XI11_6/net21_8_ xsel_23_ XI11_6/XI0/XI0_23/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_6 XI11_6/net21_9_ xsel_23_ XI11_6/XI0/XI0_23/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_5 XI11_6/net21_10_ xsel_23_ XI11_6/XI0/XI0_23/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_4 XI11_6/net21_11_ xsel_23_ XI11_6/XI0/XI0_23/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_3 XI11_6/net21_12_ xsel_23_ XI11_6/XI0/XI0_23/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_2 XI11_6/net21_13_ xsel_23_ XI11_6/XI0/XI0_23/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_1 XI11_6/net21_14_ xsel_23_ XI11_6/XI0/XI0_23/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_0 XI11_6/net21_15_ xsel_23_ XI11_6/XI0/XI0_23/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_15 XI11_6/XI0/XI0_23/d__15_ xsel_23_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_14 XI11_6/XI0/XI0_23/d__14_ xsel_23_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_13 XI11_6/XI0/XI0_23/d__13_ xsel_23_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_12 XI11_6/XI0/XI0_23/d__12_ xsel_23_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_11 XI11_6/XI0/XI0_23/d__11_ xsel_23_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_10 XI11_6/XI0/XI0_23/d__10_ xsel_23_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_9 XI11_6/XI0/XI0_23/d__9_ xsel_23_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_8 XI11_6/XI0/XI0_23/d__8_ xsel_23_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_7 XI11_6/XI0/XI0_23/d__7_ xsel_23_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_6 XI11_6/XI0/XI0_23/d__6_ xsel_23_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_5 XI11_6/XI0/XI0_23/d__5_ xsel_23_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_4 XI11_6/XI0/XI0_23/d__4_ xsel_23_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_3 XI11_6/XI0/XI0_23/d__3_ xsel_23_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_2 XI11_6/XI0/XI0_23/d__2_ xsel_23_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_1 XI11_6/XI0/XI0_23/d__1_ xsel_23_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_0 XI11_6/XI0/XI0_23/d__0_ xsel_23_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_15 XI11_6/net21_0_ xsel_22_ XI11_6/XI0/XI0_22/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_14 XI11_6/net21_1_ xsel_22_ XI11_6/XI0/XI0_22/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_13 XI11_6/net21_2_ xsel_22_ XI11_6/XI0/XI0_22/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_12 XI11_6/net21_3_ xsel_22_ XI11_6/XI0/XI0_22/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_11 XI11_6/net21_4_ xsel_22_ XI11_6/XI0/XI0_22/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_10 XI11_6/net21_5_ xsel_22_ XI11_6/XI0/XI0_22/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_9 XI11_6/net21_6_ xsel_22_ XI11_6/XI0/XI0_22/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_8 XI11_6/net21_7_ xsel_22_ XI11_6/XI0/XI0_22/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_7 XI11_6/net21_8_ xsel_22_ XI11_6/XI0/XI0_22/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_6 XI11_6/net21_9_ xsel_22_ XI11_6/XI0/XI0_22/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_5 XI11_6/net21_10_ xsel_22_ XI11_6/XI0/XI0_22/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_4 XI11_6/net21_11_ xsel_22_ XI11_6/XI0/XI0_22/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_3 XI11_6/net21_12_ xsel_22_ XI11_6/XI0/XI0_22/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_2 XI11_6/net21_13_ xsel_22_ XI11_6/XI0/XI0_22/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_1 XI11_6/net21_14_ xsel_22_ XI11_6/XI0/XI0_22/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_0 XI11_6/net21_15_ xsel_22_ XI11_6/XI0/XI0_22/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_15 XI11_6/XI0/XI0_22/d__15_ xsel_22_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_14 XI11_6/XI0/XI0_22/d__14_ xsel_22_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_13 XI11_6/XI0/XI0_22/d__13_ xsel_22_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_12 XI11_6/XI0/XI0_22/d__12_ xsel_22_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_11 XI11_6/XI0/XI0_22/d__11_ xsel_22_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_10 XI11_6/XI0/XI0_22/d__10_ xsel_22_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_9 XI11_6/XI0/XI0_22/d__9_ xsel_22_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_8 XI11_6/XI0/XI0_22/d__8_ xsel_22_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_7 XI11_6/XI0/XI0_22/d__7_ xsel_22_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_6 XI11_6/XI0/XI0_22/d__6_ xsel_22_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_5 XI11_6/XI0/XI0_22/d__5_ xsel_22_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_4 XI11_6/XI0/XI0_22/d__4_ xsel_22_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_3 XI11_6/XI0/XI0_22/d__3_ xsel_22_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_2 XI11_6/XI0/XI0_22/d__2_ xsel_22_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_1 XI11_6/XI0/XI0_22/d__1_ xsel_22_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_0 XI11_6/XI0/XI0_22/d__0_ xsel_22_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_15 XI11_6/net21_0_ xsel_21_ XI11_6/XI0/XI0_21/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_14 XI11_6/net21_1_ xsel_21_ XI11_6/XI0/XI0_21/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_13 XI11_6/net21_2_ xsel_21_ XI11_6/XI0/XI0_21/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_12 XI11_6/net21_3_ xsel_21_ XI11_6/XI0/XI0_21/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_11 XI11_6/net21_4_ xsel_21_ XI11_6/XI0/XI0_21/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_10 XI11_6/net21_5_ xsel_21_ XI11_6/XI0/XI0_21/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_9 XI11_6/net21_6_ xsel_21_ XI11_6/XI0/XI0_21/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_8 XI11_6/net21_7_ xsel_21_ XI11_6/XI0/XI0_21/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_7 XI11_6/net21_8_ xsel_21_ XI11_6/XI0/XI0_21/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_6 XI11_6/net21_9_ xsel_21_ XI11_6/XI0/XI0_21/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_5 XI11_6/net21_10_ xsel_21_ XI11_6/XI0/XI0_21/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_4 XI11_6/net21_11_ xsel_21_ XI11_6/XI0/XI0_21/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_3 XI11_6/net21_12_ xsel_21_ XI11_6/XI0/XI0_21/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_2 XI11_6/net21_13_ xsel_21_ XI11_6/XI0/XI0_21/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_1 XI11_6/net21_14_ xsel_21_ XI11_6/XI0/XI0_21/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_0 XI11_6/net21_15_ xsel_21_ XI11_6/XI0/XI0_21/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_15 XI11_6/XI0/XI0_21/d__15_ xsel_21_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_14 XI11_6/XI0/XI0_21/d__14_ xsel_21_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_13 XI11_6/XI0/XI0_21/d__13_ xsel_21_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_12 XI11_6/XI0/XI0_21/d__12_ xsel_21_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_11 XI11_6/XI0/XI0_21/d__11_ xsel_21_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_10 XI11_6/XI0/XI0_21/d__10_ xsel_21_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_9 XI11_6/XI0/XI0_21/d__9_ xsel_21_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_8 XI11_6/XI0/XI0_21/d__8_ xsel_21_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_7 XI11_6/XI0/XI0_21/d__7_ xsel_21_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_6 XI11_6/XI0/XI0_21/d__6_ xsel_21_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_5 XI11_6/XI0/XI0_21/d__5_ xsel_21_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_4 XI11_6/XI0/XI0_21/d__4_ xsel_21_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_3 XI11_6/XI0/XI0_21/d__3_ xsel_21_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_2 XI11_6/XI0/XI0_21/d__2_ xsel_21_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_1 XI11_6/XI0/XI0_21/d__1_ xsel_21_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_0 XI11_6/XI0/XI0_21/d__0_ xsel_21_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_15 XI11_6/net21_0_ xsel_20_ XI11_6/XI0/XI0_20/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_14 XI11_6/net21_1_ xsel_20_ XI11_6/XI0/XI0_20/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_13 XI11_6/net21_2_ xsel_20_ XI11_6/XI0/XI0_20/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_12 XI11_6/net21_3_ xsel_20_ XI11_6/XI0/XI0_20/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_11 XI11_6/net21_4_ xsel_20_ XI11_6/XI0/XI0_20/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_10 XI11_6/net21_5_ xsel_20_ XI11_6/XI0/XI0_20/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_9 XI11_6/net21_6_ xsel_20_ XI11_6/XI0/XI0_20/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_8 XI11_6/net21_7_ xsel_20_ XI11_6/XI0/XI0_20/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_7 XI11_6/net21_8_ xsel_20_ XI11_6/XI0/XI0_20/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_6 XI11_6/net21_9_ xsel_20_ XI11_6/XI0/XI0_20/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_5 XI11_6/net21_10_ xsel_20_ XI11_6/XI0/XI0_20/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_4 XI11_6/net21_11_ xsel_20_ XI11_6/XI0/XI0_20/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_3 XI11_6/net21_12_ xsel_20_ XI11_6/XI0/XI0_20/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_2 XI11_6/net21_13_ xsel_20_ XI11_6/XI0/XI0_20/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_1 XI11_6/net21_14_ xsel_20_ XI11_6/XI0/XI0_20/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_0 XI11_6/net21_15_ xsel_20_ XI11_6/XI0/XI0_20/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_15 XI11_6/XI0/XI0_20/d__15_ xsel_20_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_14 XI11_6/XI0/XI0_20/d__14_ xsel_20_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_13 XI11_6/XI0/XI0_20/d__13_ xsel_20_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_12 XI11_6/XI0/XI0_20/d__12_ xsel_20_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_11 XI11_6/XI0/XI0_20/d__11_ xsel_20_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_10 XI11_6/XI0/XI0_20/d__10_ xsel_20_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_9 XI11_6/XI0/XI0_20/d__9_ xsel_20_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_8 XI11_6/XI0/XI0_20/d__8_ xsel_20_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_7 XI11_6/XI0/XI0_20/d__7_ xsel_20_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_6 XI11_6/XI0/XI0_20/d__6_ xsel_20_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_5 XI11_6/XI0/XI0_20/d__5_ xsel_20_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_4 XI11_6/XI0/XI0_20/d__4_ xsel_20_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_3 XI11_6/XI0/XI0_20/d__3_ xsel_20_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_2 XI11_6/XI0/XI0_20/d__2_ xsel_20_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_1 XI11_6/XI0/XI0_20/d__1_ xsel_20_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_0 XI11_6/XI0/XI0_20/d__0_ xsel_20_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_15 XI11_6/net21_0_ xsel_19_ XI11_6/XI0/XI0_19/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_14 XI11_6/net21_1_ xsel_19_ XI11_6/XI0/XI0_19/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_13 XI11_6/net21_2_ xsel_19_ XI11_6/XI0/XI0_19/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_12 XI11_6/net21_3_ xsel_19_ XI11_6/XI0/XI0_19/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_11 XI11_6/net21_4_ xsel_19_ XI11_6/XI0/XI0_19/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_10 XI11_6/net21_5_ xsel_19_ XI11_6/XI0/XI0_19/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_9 XI11_6/net21_6_ xsel_19_ XI11_6/XI0/XI0_19/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_8 XI11_6/net21_7_ xsel_19_ XI11_6/XI0/XI0_19/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_7 XI11_6/net21_8_ xsel_19_ XI11_6/XI0/XI0_19/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_6 XI11_6/net21_9_ xsel_19_ XI11_6/XI0/XI0_19/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_5 XI11_6/net21_10_ xsel_19_ XI11_6/XI0/XI0_19/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_4 XI11_6/net21_11_ xsel_19_ XI11_6/XI0/XI0_19/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_3 XI11_6/net21_12_ xsel_19_ XI11_6/XI0/XI0_19/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_2 XI11_6/net21_13_ xsel_19_ XI11_6/XI0/XI0_19/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_1 XI11_6/net21_14_ xsel_19_ XI11_6/XI0/XI0_19/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_0 XI11_6/net21_15_ xsel_19_ XI11_6/XI0/XI0_19/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_15 XI11_6/XI0/XI0_19/d__15_ xsel_19_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_14 XI11_6/XI0/XI0_19/d__14_ xsel_19_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_13 XI11_6/XI0/XI0_19/d__13_ xsel_19_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_12 XI11_6/XI0/XI0_19/d__12_ xsel_19_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_11 XI11_6/XI0/XI0_19/d__11_ xsel_19_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_10 XI11_6/XI0/XI0_19/d__10_ xsel_19_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_9 XI11_6/XI0/XI0_19/d__9_ xsel_19_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_8 XI11_6/XI0/XI0_19/d__8_ xsel_19_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_7 XI11_6/XI0/XI0_19/d__7_ xsel_19_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_6 XI11_6/XI0/XI0_19/d__6_ xsel_19_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_5 XI11_6/XI0/XI0_19/d__5_ xsel_19_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_4 XI11_6/XI0/XI0_19/d__4_ xsel_19_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_3 XI11_6/XI0/XI0_19/d__3_ xsel_19_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_2 XI11_6/XI0/XI0_19/d__2_ xsel_19_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_1 XI11_6/XI0/XI0_19/d__1_ xsel_19_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_0 XI11_6/XI0/XI0_19/d__0_ xsel_19_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_15 XI11_6/net21_0_ xsel_18_ XI11_6/XI0/XI0_18/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_14 XI11_6/net21_1_ xsel_18_ XI11_6/XI0/XI0_18/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_13 XI11_6/net21_2_ xsel_18_ XI11_6/XI0/XI0_18/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_12 XI11_6/net21_3_ xsel_18_ XI11_6/XI0/XI0_18/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_11 XI11_6/net21_4_ xsel_18_ XI11_6/XI0/XI0_18/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_10 XI11_6/net21_5_ xsel_18_ XI11_6/XI0/XI0_18/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_9 XI11_6/net21_6_ xsel_18_ XI11_6/XI0/XI0_18/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_8 XI11_6/net21_7_ xsel_18_ XI11_6/XI0/XI0_18/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_7 XI11_6/net21_8_ xsel_18_ XI11_6/XI0/XI0_18/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_6 XI11_6/net21_9_ xsel_18_ XI11_6/XI0/XI0_18/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_5 XI11_6/net21_10_ xsel_18_ XI11_6/XI0/XI0_18/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_4 XI11_6/net21_11_ xsel_18_ XI11_6/XI0/XI0_18/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_3 XI11_6/net21_12_ xsel_18_ XI11_6/XI0/XI0_18/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_2 XI11_6/net21_13_ xsel_18_ XI11_6/XI0/XI0_18/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_1 XI11_6/net21_14_ xsel_18_ XI11_6/XI0/XI0_18/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_0 XI11_6/net21_15_ xsel_18_ XI11_6/XI0/XI0_18/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_15 XI11_6/XI0/XI0_18/d__15_ xsel_18_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_14 XI11_6/XI0/XI0_18/d__14_ xsel_18_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_13 XI11_6/XI0/XI0_18/d__13_ xsel_18_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_12 XI11_6/XI0/XI0_18/d__12_ xsel_18_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_11 XI11_6/XI0/XI0_18/d__11_ xsel_18_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_10 XI11_6/XI0/XI0_18/d__10_ xsel_18_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_9 XI11_6/XI0/XI0_18/d__9_ xsel_18_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_8 XI11_6/XI0/XI0_18/d__8_ xsel_18_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_7 XI11_6/XI0/XI0_18/d__7_ xsel_18_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_6 XI11_6/XI0/XI0_18/d__6_ xsel_18_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_5 XI11_6/XI0/XI0_18/d__5_ xsel_18_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_4 XI11_6/XI0/XI0_18/d__4_ xsel_18_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_3 XI11_6/XI0/XI0_18/d__3_ xsel_18_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_2 XI11_6/XI0/XI0_18/d__2_ xsel_18_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_1 XI11_6/XI0/XI0_18/d__1_ xsel_18_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_0 XI11_6/XI0/XI0_18/d__0_ xsel_18_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_15 XI11_6/net21_0_ xsel_17_ XI11_6/XI0/XI0_17/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_14 XI11_6/net21_1_ xsel_17_ XI11_6/XI0/XI0_17/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_13 XI11_6/net21_2_ xsel_17_ XI11_6/XI0/XI0_17/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_12 XI11_6/net21_3_ xsel_17_ XI11_6/XI0/XI0_17/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_11 XI11_6/net21_4_ xsel_17_ XI11_6/XI0/XI0_17/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_10 XI11_6/net21_5_ xsel_17_ XI11_6/XI0/XI0_17/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_9 XI11_6/net21_6_ xsel_17_ XI11_6/XI0/XI0_17/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_8 XI11_6/net21_7_ xsel_17_ XI11_6/XI0/XI0_17/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_7 XI11_6/net21_8_ xsel_17_ XI11_6/XI0/XI0_17/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_6 XI11_6/net21_9_ xsel_17_ XI11_6/XI0/XI0_17/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_5 XI11_6/net21_10_ xsel_17_ XI11_6/XI0/XI0_17/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_4 XI11_6/net21_11_ xsel_17_ XI11_6/XI0/XI0_17/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_3 XI11_6/net21_12_ xsel_17_ XI11_6/XI0/XI0_17/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_2 XI11_6/net21_13_ xsel_17_ XI11_6/XI0/XI0_17/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_1 XI11_6/net21_14_ xsel_17_ XI11_6/XI0/XI0_17/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_0 XI11_6/net21_15_ xsel_17_ XI11_6/XI0/XI0_17/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_15 XI11_6/XI0/XI0_17/d__15_ xsel_17_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_14 XI11_6/XI0/XI0_17/d__14_ xsel_17_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_13 XI11_6/XI0/XI0_17/d__13_ xsel_17_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_12 XI11_6/XI0/XI0_17/d__12_ xsel_17_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_11 XI11_6/XI0/XI0_17/d__11_ xsel_17_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_10 XI11_6/XI0/XI0_17/d__10_ xsel_17_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_9 XI11_6/XI0/XI0_17/d__9_ xsel_17_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_8 XI11_6/XI0/XI0_17/d__8_ xsel_17_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_7 XI11_6/XI0/XI0_17/d__7_ xsel_17_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_6 XI11_6/XI0/XI0_17/d__6_ xsel_17_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_5 XI11_6/XI0/XI0_17/d__5_ xsel_17_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_4 XI11_6/XI0/XI0_17/d__4_ xsel_17_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_3 XI11_6/XI0/XI0_17/d__3_ xsel_17_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_2 XI11_6/XI0/XI0_17/d__2_ xsel_17_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_1 XI11_6/XI0/XI0_17/d__1_ xsel_17_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_0 XI11_6/XI0/XI0_17/d__0_ xsel_17_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_15 XI11_6/net21_0_ xsel_16_ XI11_6/XI0/XI0_16/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_14 XI11_6/net21_1_ xsel_16_ XI11_6/XI0/XI0_16/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_13 XI11_6/net21_2_ xsel_16_ XI11_6/XI0/XI0_16/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_12 XI11_6/net21_3_ xsel_16_ XI11_6/XI0/XI0_16/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_11 XI11_6/net21_4_ xsel_16_ XI11_6/XI0/XI0_16/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_10 XI11_6/net21_5_ xsel_16_ XI11_6/XI0/XI0_16/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_9 XI11_6/net21_6_ xsel_16_ XI11_6/XI0/XI0_16/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_8 XI11_6/net21_7_ xsel_16_ XI11_6/XI0/XI0_16/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_7 XI11_6/net21_8_ xsel_16_ XI11_6/XI0/XI0_16/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_6 XI11_6/net21_9_ xsel_16_ XI11_6/XI0/XI0_16/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_5 XI11_6/net21_10_ xsel_16_ XI11_6/XI0/XI0_16/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_4 XI11_6/net21_11_ xsel_16_ XI11_6/XI0/XI0_16/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_3 XI11_6/net21_12_ xsel_16_ XI11_6/XI0/XI0_16/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_2 XI11_6/net21_13_ xsel_16_ XI11_6/XI0/XI0_16/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_1 XI11_6/net21_14_ xsel_16_ XI11_6/XI0/XI0_16/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_0 XI11_6/net21_15_ xsel_16_ XI11_6/XI0/XI0_16/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_15 XI11_6/XI0/XI0_16/d__15_ xsel_16_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_14 XI11_6/XI0/XI0_16/d__14_ xsel_16_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_13 XI11_6/XI0/XI0_16/d__13_ xsel_16_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_12 XI11_6/XI0/XI0_16/d__12_ xsel_16_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_11 XI11_6/XI0/XI0_16/d__11_ xsel_16_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_10 XI11_6/XI0/XI0_16/d__10_ xsel_16_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_9 XI11_6/XI0/XI0_16/d__9_ xsel_16_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_8 XI11_6/XI0/XI0_16/d__8_ xsel_16_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_7 XI11_6/XI0/XI0_16/d__7_ xsel_16_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_6 XI11_6/XI0/XI0_16/d__6_ xsel_16_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_5 XI11_6/XI0/XI0_16/d__5_ xsel_16_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_4 XI11_6/XI0/XI0_16/d__4_ xsel_16_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_3 XI11_6/XI0/XI0_16/d__3_ xsel_16_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_2 XI11_6/XI0/XI0_16/d__2_ xsel_16_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_1 XI11_6/XI0/XI0_16/d__1_ xsel_16_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_0 XI11_6/XI0/XI0_16/d__0_ xsel_16_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_15 XI11_6/net21_0_ xsel_15_ XI11_6/XI0/XI0_15/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_14 XI11_6/net21_1_ xsel_15_ XI11_6/XI0/XI0_15/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_13 XI11_6/net21_2_ xsel_15_ XI11_6/XI0/XI0_15/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_12 XI11_6/net21_3_ xsel_15_ XI11_6/XI0/XI0_15/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_11 XI11_6/net21_4_ xsel_15_ XI11_6/XI0/XI0_15/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_10 XI11_6/net21_5_ xsel_15_ XI11_6/XI0/XI0_15/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_9 XI11_6/net21_6_ xsel_15_ XI11_6/XI0/XI0_15/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_8 XI11_6/net21_7_ xsel_15_ XI11_6/XI0/XI0_15/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_7 XI11_6/net21_8_ xsel_15_ XI11_6/XI0/XI0_15/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_6 XI11_6/net21_9_ xsel_15_ XI11_6/XI0/XI0_15/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_5 XI11_6/net21_10_ xsel_15_ XI11_6/XI0/XI0_15/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_4 XI11_6/net21_11_ xsel_15_ XI11_6/XI0/XI0_15/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_3 XI11_6/net21_12_ xsel_15_ XI11_6/XI0/XI0_15/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_2 XI11_6/net21_13_ xsel_15_ XI11_6/XI0/XI0_15/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_1 XI11_6/net21_14_ xsel_15_ XI11_6/XI0/XI0_15/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_0 XI11_6/net21_15_ xsel_15_ XI11_6/XI0/XI0_15/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_15 XI11_6/XI0/XI0_15/d__15_ xsel_15_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_14 XI11_6/XI0/XI0_15/d__14_ xsel_15_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_13 XI11_6/XI0/XI0_15/d__13_ xsel_15_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_12 XI11_6/XI0/XI0_15/d__12_ xsel_15_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_11 XI11_6/XI0/XI0_15/d__11_ xsel_15_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_10 XI11_6/XI0/XI0_15/d__10_ xsel_15_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_9 XI11_6/XI0/XI0_15/d__9_ xsel_15_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_8 XI11_6/XI0/XI0_15/d__8_ xsel_15_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_7 XI11_6/XI0/XI0_15/d__7_ xsel_15_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_6 XI11_6/XI0/XI0_15/d__6_ xsel_15_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_5 XI11_6/XI0/XI0_15/d__5_ xsel_15_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_4 XI11_6/XI0/XI0_15/d__4_ xsel_15_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_3 XI11_6/XI0/XI0_15/d__3_ xsel_15_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_2 XI11_6/XI0/XI0_15/d__2_ xsel_15_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_1 XI11_6/XI0/XI0_15/d__1_ xsel_15_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_0 XI11_6/XI0/XI0_15/d__0_ xsel_15_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_15 XI11_6/net21_0_ xsel_14_ XI11_6/XI0/XI0_14/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_14 XI11_6/net21_1_ xsel_14_ XI11_6/XI0/XI0_14/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_13 XI11_6/net21_2_ xsel_14_ XI11_6/XI0/XI0_14/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_12 XI11_6/net21_3_ xsel_14_ XI11_6/XI0/XI0_14/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_11 XI11_6/net21_4_ xsel_14_ XI11_6/XI0/XI0_14/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_10 XI11_6/net21_5_ xsel_14_ XI11_6/XI0/XI0_14/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_9 XI11_6/net21_6_ xsel_14_ XI11_6/XI0/XI0_14/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_8 XI11_6/net21_7_ xsel_14_ XI11_6/XI0/XI0_14/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_7 XI11_6/net21_8_ xsel_14_ XI11_6/XI0/XI0_14/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_6 XI11_6/net21_9_ xsel_14_ XI11_6/XI0/XI0_14/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_5 XI11_6/net21_10_ xsel_14_ XI11_6/XI0/XI0_14/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_4 XI11_6/net21_11_ xsel_14_ XI11_6/XI0/XI0_14/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_3 XI11_6/net21_12_ xsel_14_ XI11_6/XI0/XI0_14/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_2 XI11_6/net21_13_ xsel_14_ XI11_6/XI0/XI0_14/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_1 XI11_6/net21_14_ xsel_14_ XI11_6/XI0/XI0_14/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_0 XI11_6/net21_15_ xsel_14_ XI11_6/XI0/XI0_14/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_15 XI11_6/XI0/XI0_14/d__15_ xsel_14_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_14 XI11_6/XI0/XI0_14/d__14_ xsel_14_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_13 XI11_6/XI0/XI0_14/d__13_ xsel_14_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_12 XI11_6/XI0/XI0_14/d__12_ xsel_14_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_11 XI11_6/XI0/XI0_14/d__11_ xsel_14_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_10 XI11_6/XI0/XI0_14/d__10_ xsel_14_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_9 XI11_6/XI0/XI0_14/d__9_ xsel_14_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_8 XI11_6/XI0/XI0_14/d__8_ xsel_14_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_7 XI11_6/XI0/XI0_14/d__7_ xsel_14_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_6 XI11_6/XI0/XI0_14/d__6_ xsel_14_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_5 XI11_6/XI0/XI0_14/d__5_ xsel_14_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_4 XI11_6/XI0/XI0_14/d__4_ xsel_14_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_3 XI11_6/XI0/XI0_14/d__3_ xsel_14_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_2 XI11_6/XI0/XI0_14/d__2_ xsel_14_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_1 XI11_6/XI0/XI0_14/d__1_ xsel_14_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_0 XI11_6/XI0/XI0_14/d__0_ xsel_14_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_15 XI11_6/net21_0_ xsel_13_ XI11_6/XI0/XI0_13/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_14 XI11_6/net21_1_ xsel_13_ XI11_6/XI0/XI0_13/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_13 XI11_6/net21_2_ xsel_13_ XI11_6/XI0/XI0_13/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_12 XI11_6/net21_3_ xsel_13_ XI11_6/XI0/XI0_13/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_11 XI11_6/net21_4_ xsel_13_ XI11_6/XI0/XI0_13/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_10 XI11_6/net21_5_ xsel_13_ XI11_6/XI0/XI0_13/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_9 XI11_6/net21_6_ xsel_13_ XI11_6/XI0/XI0_13/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_8 XI11_6/net21_7_ xsel_13_ XI11_6/XI0/XI0_13/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_7 XI11_6/net21_8_ xsel_13_ XI11_6/XI0/XI0_13/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_6 XI11_6/net21_9_ xsel_13_ XI11_6/XI0/XI0_13/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_5 XI11_6/net21_10_ xsel_13_ XI11_6/XI0/XI0_13/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_4 XI11_6/net21_11_ xsel_13_ XI11_6/XI0/XI0_13/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_3 XI11_6/net21_12_ xsel_13_ XI11_6/XI0/XI0_13/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_2 XI11_6/net21_13_ xsel_13_ XI11_6/XI0/XI0_13/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_1 XI11_6/net21_14_ xsel_13_ XI11_6/XI0/XI0_13/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_0 XI11_6/net21_15_ xsel_13_ XI11_6/XI0/XI0_13/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_15 XI11_6/XI0/XI0_13/d__15_ xsel_13_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_14 XI11_6/XI0/XI0_13/d__14_ xsel_13_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_13 XI11_6/XI0/XI0_13/d__13_ xsel_13_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_12 XI11_6/XI0/XI0_13/d__12_ xsel_13_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_11 XI11_6/XI0/XI0_13/d__11_ xsel_13_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_10 XI11_6/XI0/XI0_13/d__10_ xsel_13_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_9 XI11_6/XI0/XI0_13/d__9_ xsel_13_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_8 XI11_6/XI0/XI0_13/d__8_ xsel_13_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_7 XI11_6/XI0/XI0_13/d__7_ xsel_13_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_6 XI11_6/XI0/XI0_13/d__6_ xsel_13_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_5 XI11_6/XI0/XI0_13/d__5_ xsel_13_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_4 XI11_6/XI0/XI0_13/d__4_ xsel_13_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_3 XI11_6/XI0/XI0_13/d__3_ xsel_13_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_2 XI11_6/XI0/XI0_13/d__2_ xsel_13_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_1 XI11_6/XI0/XI0_13/d__1_ xsel_13_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_0 XI11_6/XI0/XI0_13/d__0_ xsel_13_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_15 XI11_6/net21_0_ xsel_12_ XI11_6/XI0/XI0_12/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_14 XI11_6/net21_1_ xsel_12_ XI11_6/XI0/XI0_12/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_13 XI11_6/net21_2_ xsel_12_ XI11_6/XI0/XI0_12/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_12 XI11_6/net21_3_ xsel_12_ XI11_6/XI0/XI0_12/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_11 XI11_6/net21_4_ xsel_12_ XI11_6/XI0/XI0_12/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_10 XI11_6/net21_5_ xsel_12_ XI11_6/XI0/XI0_12/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_9 XI11_6/net21_6_ xsel_12_ XI11_6/XI0/XI0_12/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_8 XI11_6/net21_7_ xsel_12_ XI11_6/XI0/XI0_12/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_7 XI11_6/net21_8_ xsel_12_ XI11_6/XI0/XI0_12/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_6 XI11_6/net21_9_ xsel_12_ XI11_6/XI0/XI0_12/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_5 XI11_6/net21_10_ xsel_12_ XI11_6/XI0/XI0_12/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_4 XI11_6/net21_11_ xsel_12_ XI11_6/XI0/XI0_12/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_3 XI11_6/net21_12_ xsel_12_ XI11_6/XI0/XI0_12/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_2 XI11_6/net21_13_ xsel_12_ XI11_6/XI0/XI0_12/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_1 XI11_6/net21_14_ xsel_12_ XI11_6/XI0/XI0_12/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_0 XI11_6/net21_15_ xsel_12_ XI11_6/XI0/XI0_12/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_15 XI11_6/XI0/XI0_12/d__15_ xsel_12_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_14 XI11_6/XI0/XI0_12/d__14_ xsel_12_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_13 XI11_6/XI0/XI0_12/d__13_ xsel_12_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_12 XI11_6/XI0/XI0_12/d__12_ xsel_12_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_11 XI11_6/XI0/XI0_12/d__11_ xsel_12_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_10 XI11_6/XI0/XI0_12/d__10_ xsel_12_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_9 XI11_6/XI0/XI0_12/d__9_ xsel_12_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_8 XI11_6/XI0/XI0_12/d__8_ xsel_12_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_7 XI11_6/XI0/XI0_12/d__7_ xsel_12_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_6 XI11_6/XI0/XI0_12/d__6_ xsel_12_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_5 XI11_6/XI0/XI0_12/d__5_ xsel_12_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_4 XI11_6/XI0/XI0_12/d__4_ xsel_12_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_3 XI11_6/XI0/XI0_12/d__3_ xsel_12_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_2 XI11_6/XI0/XI0_12/d__2_ xsel_12_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_1 XI11_6/XI0/XI0_12/d__1_ xsel_12_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_0 XI11_6/XI0/XI0_12/d__0_ xsel_12_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_15 XI11_6/net21_0_ xsel_11_ XI11_6/XI0/XI0_11/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_14 XI11_6/net21_1_ xsel_11_ XI11_6/XI0/XI0_11/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_13 XI11_6/net21_2_ xsel_11_ XI11_6/XI0/XI0_11/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_12 XI11_6/net21_3_ xsel_11_ XI11_6/XI0/XI0_11/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_11 XI11_6/net21_4_ xsel_11_ XI11_6/XI0/XI0_11/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_10 XI11_6/net21_5_ xsel_11_ XI11_6/XI0/XI0_11/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_9 XI11_6/net21_6_ xsel_11_ XI11_6/XI0/XI0_11/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_8 XI11_6/net21_7_ xsel_11_ XI11_6/XI0/XI0_11/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_7 XI11_6/net21_8_ xsel_11_ XI11_6/XI0/XI0_11/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_6 XI11_6/net21_9_ xsel_11_ XI11_6/XI0/XI0_11/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_5 XI11_6/net21_10_ xsel_11_ XI11_6/XI0/XI0_11/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_4 XI11_6/net21_11_ xsel_11_ XI11_6/XI0/XI0_11/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_3 XI11_6/net21_12_ xsel_11_ XI11_6/XI0/XI0_11/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_2 XI11_6/net21_13_ xsel_11_ XI11_6/XI0/XI0_11/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_1 XI11_6/net21_14_ xsel_11_ XI11_6/XI0/XI0_11/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_0 XI11_6/net21_15_ xsel_11_ XI11_6/XI0/XI0_11/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_15 XI11_6/XI0/XI0_11/d__15_ xsel_11_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_14 XI11_6/XI0/XI0_11/d__14_ xsel_11_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_13 XI11_6/XI0/XI0_11/d__13_ xsel_11_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_12 XI11_6/XI0/XI0_11/d__12_ xsel_11_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_11 XI11_6/XI0/XI0_11/d__11_ xsel_11_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_10 XI11_6/XI0/XI0_11/d__10_ xsel_11_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_9 XI11_6/XI0/XI0_11/d__9_ xsel_11_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_8 XI11_6/XI0/XI0_11/d__8_ xsel_11_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_7 XI11_6/XI0/XI0_11/d__7_ xsel_11_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_6 XI11_6/XI0/XI0_11/d__6_ xsel_11_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_5 XI11_6/XI0/XI0_11/d__5_ xsel_11_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_4 XI11_6/XI0/XI0_11/d__4_ xsel_11_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_3 XI11_6/XI0/XI0_11/d__3_ xsel_11_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_2 XI11_6/XI0/XI0_11/d__2_ xsel_11_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_1 XI11_6/XI0/XI0_11/d__1_ xsel_11_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_0 XI11_6/XI0/XI0_11/d__0_ xsel_11_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_15 XI11_6/net21_0_ xsel_10_ XI11_6/XI0/XI0_10/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_14 XI11_6/net21_1_ xsel_10_ XI11_6/XI0/XI0_10/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_13 XI11_6/net21_2_ xsel_10_ XI11_6/XI0/XI0_10/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_12 XI11_6/net21_3_ xsel_10_ XI11_6/XI0/XI0_10/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_11 XI11_6/net21_4_ xsel_10_ XI11_6/XI0/XI0_10/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_10 XI11_6/net21_5_ xsel_10_ XI11_6/XI0/XI0_10/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_9 XI11_6/net21_6_ xsel_10_ XI11_6/XI0/XI0_10/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_8 XI11_6/net21_7_ xsel_10_ XI11_6/XI0/XI0_10/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_7 XI11_6/net21_8_ xsel_10_ XI11_6/XI0/XI0_10/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_6 XI11_6/net21_9_ xsel_10_ XI11_6/XI0/XI0_10/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_5 XI11_6/net21_10_ xsel_10_ XI11_6/XI0/XI0_10/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_4 XI11_6/net21_11_ xsel_10_ XI11_6/XI0/XI0_10/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_3 XI11_6/net21_12_ xsel_10_ XI11_6/XI0/XI0_10/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_2 XI11_6/net21_13_ xsel_10_ XI11_6/XI0/XI0_10/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_1 XI11_6/net21_14_ xsel_10_ XI11_6/XI0/XI0_10/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_0 XI11_6/net21_15_ xsel_10_ XI11_6/XI0/XI0_10/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_15 XI11_6/XI0/XI0_10/d__15_ xsel_10_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_14 XI11_6/XI0/XI0_10/d__14_ xsel_10_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_13 XI11_6/XI0/XI0_10/d__13_ xsel_10_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_12 XI11_6/XI0/XI0_10/d__12_ xsel_10_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_11 XI11_6/XI0/XI0_10/d__11_ xsel_10_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_10 XI11_6/XI0/XI0_10/d__10_ xsel_10_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_9 XI11_6/XI0/XI0_10/d__9_ xsel_10_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_8 XI11_6/XI0/XI0_10/d__8_ xsel_10_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_7 XI11_6/XI0/XI0_10/d__7_ xsel_10_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_6 XI11_6/XI0/XI0_10/d__6_ xsel_10_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_5 XI11_6/XI0/XI0_10/d__5_ xsel_10_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_4 XI11_6/XI0/XI0_10/d__4_ xsel_10_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_3 XI11_6/XI0/XI0_10/d__3_ xsel_10_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_2 XI11_6/XI0/XI0_10/d__2_ xsel_10_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_1 XI11_6/XI0/XI0_10/d__1_ xsel_10_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_0 XI11_6/XI0/XI0_10/d__0_ xsel_10_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_15 XI11_6/net21_0_ xsel_9_ XI11_6/XI0/XI0_9/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_14 XI11_6/net21_1_ xsel_9_ XI11_6/XI0/XI0_9/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_13 XI11_6/net21_2_ xsel_9_ XI11_6/XI0/XI0_9/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_12 XI11_6/net21_3_ xsel_9_ XI11_6/XI0/XI0_9/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_11 XI11_6/net21_4_ xsel_9_ XI11_6/XI0/XI0_9/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_10 XI11_6/net21_5_ xsel_9_ XI11_6/XI0/XI0_9/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_9 XI11_6/net21_6_ xsel_9_ XI11_6/XI0/XI0_9/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_8 XI11_6/net21_7_ xsel_9_ XI11_6/XI0/XI0_9/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_7 XI11_6/net21_8_ xsel_9_ XI11_6/XI0/XI0_9/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_6 XI11_6/net21_9_ xsel_9_ XI11_6/XI0/XI0_9/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_5 XI11_6/net21_10_ xsel_9_ XI11_6/XI0/XI0_9/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_4 XI11_6/net21_11_ xsel_9_ XI11_6/XI0/XI0_9/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_3 XI11_6/net21_12_ xsel_9_ XI11_6/XI0/XI0_9/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_2 XI11_6/net21_13_ xsel_9_ XI11_6/XI0/XI0_9/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_1 XI11_6/net21_14_ xsel_9_ XI11_6/XI0/XI0_9/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_0 XI11_6/net21_15_ xsel_9_ XI11_6/XI0/XI0_9/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_15 XI11_6/XI0/XI0_9/d__15_ xsel_9_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_14 XI11_6/XI0/XI0_9/d__14_ xsel_9_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_13 XI11_6/XI0/XI0_9/d__13_ xsel_9_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_12 XI11_6/XI0/XI0_9/d__12_ xsel_9_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_11 XI11_6/XI0/XI0_9/d__11_ xsel_9_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_10 XI11_6/XI0/XI0_9/d__10_ xsel_9_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_9 XI11_6/XI0/XI0_9/d__9_ xsel_9_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_8 XI11_6/XI0/XI0_9/d__8_ xsel_9_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_7 XI11_6/XI0/XI0_9/d__7_ xsel_9_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_6 XI11_6/XI0/XI0_9/d__6_ xsel_9_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_5 XI11_6/XI0/XI0_9/d__5_ xsel_9_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_4 XI11_6/XI0/XI0_9/d__4_ xsel_9_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_3 XI11_6/XI0/XI0_9/d__3_ xsel_9_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_2 XI11_6/XI0/XI0_9/d__2_ xsel_9_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_1 XI11_6/XI0/XI0_9/d__1_ xsel_9_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_0 XI11_6/XI0/XI0_9/d__0_ xsel_9_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_15 XI11_6/net21_0_ xsel_8_ XI11_6/XI0/XI0_8/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_14 XI11_6/net21_1_ xsel_8_ XI11_6/XI0/XI0_8/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_13 XI11_6/net21_2_ xsel_8_ XI11_6/XI0/XI0_8/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_12 XI11_6/net21_3_ xsel_8_ XI11_6/XI0/XI0_8/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_11 XI11_6/net21_4_ xsel_8_ XI11_6/XI0/XI0_8/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_10 XI11_6/net21_5_ xsel_8_ XI11_6/XI0/XI0_8/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_9 XI11_6/net21_6_ xsel_8_ XI11_6/XI0/XI0_8/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_8 XI11_6/net21_7_ xsel_8_ XI11_6/XI0/XI0_8/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_7 XI11_6/net21_8_ xsel_8_ XI11_6/XI0/XI0_8/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_6 XI11_6/net21_9_ xsel_8_ XI11_6/XI0/XI0_8/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_5 XI11_6/net21_10_ xsel_8_ XI11_6/XI0/XI0_8/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_4 XI11_6/net21_11_ xsel_8_ XI11_6/XI0/XI0_8/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_3 XI11_6/net21_12_ xsel_8_ XI11_6/XI0/XI0_8/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_2 XI11_6/net21_13_ xsel_8_ XI11_6/XI0/XI0_8/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_1 XI11_6/net21_14_ xsel_8_ XI11_6/XI0/XI0_8/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_0 XI11_6/net21_15_ xsel_8_ XI11_6/XI0/XI0_8/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_15 XI11_6/XI0/XI0_8/d__15_ xsel_8_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_14 XI11_6/XI0/XI0_8/d__14_ xsel_8_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_13 XI11_6/XI0/XI0_8/d__13_ xsel_8_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_12 XI11_6/XI0/XI0_8/d__12_ xsel_8_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_11 XI11_6/XI0/XI0_8/d__11_ xsel_8_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_10 XI11_6/XI0/XI0_8/d__10_ xsel_8_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_9 XI11_6/XI0/XI0_8/d__9_ xsel_8_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_8 XI11_6/XI0/XI0_8/d__8_ xsel_8_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_7 XI11_6/XI0/XI0_8/d__7_ xsel_8_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_6 XI11_6/XI0/XI0_8/d__6_ xsel_8_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_5 XI11_6/XI0/XI0_8/d__5_ xsel_8_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_4 XI11_6/XI0/XI0_8/d__4_ xsel_8_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_3 XI11_6/XI0/XI0_8/d__3_ xsel_8_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_2 XI11_6/XI0/XI0_8/d__2_ xsel_8_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_1 XI11_6/XI0/XI0_8/d__1_ xsel_8_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_0 XI11_6/XI0/XI0_8/d__0_ xsel_8_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_15 XI11_6/net21_0_ xsel_7_ XI11_6/XI0/XI0_7/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_14 XI11_6/net21_1_ xsel_7_ XI11_6/XI0/XI0_7/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_13 XI11_6/net21_2_ xsel_7_ XI11_6/XI0/XI0_7/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_12 XI11_6/net21_3_ xsel_7_ XI11_6/XI0/XI0_7/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_11 XI11_6/net21_4_ xsel_7_ XI11_6/XI0/XI0_7/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_10 XI11_6/net21_5_ xsel_7_ XI11_6/XI0/XI0_7/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_9 XI11_6/net21_6_ xsel_7_ XI11_6/XI0/XI0_7/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_8 XI11_6/net21_7_ xsel_7_ XI11_6/XI0/XI0_7/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_7 XI11_6/net21_8_ xsel_7_ XI11_6/XI0/XI0_7/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_6 XI11_6/net21_9_ xsel_7_ XI11_6/XI0/XI0_7/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_5 XI11_6/net21_10_ xsel_7_ XI11_6/XI0/XI0_7/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_4 XI11_6/net21_11_ xsel_7_ XI11_6/XI0/XI0_7/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_3 XI11_6/net21_12_ xsel_7_ XI11_6/XI0/XI0_7/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_2 XI11_6/net21_13_ xsel_7_ XI11_6/XI0/XI0_7/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_1 XI11_6/net21_14_ xsel_7_ XI11_6/XI0/XI0_7/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_0 XI11_6/net21_15_ xsel_7_ XI11_6/XI0/XI0_7/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_15 XI11_6/XI0/XI0_7/d__15_ xsel_7_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_14 XI11_6/XI0/XI0_7/d__14_ xsel_7_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_13 XI11_6/XI0/XI0_7/d__13_ xsel_7_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_12 XI11_6/XI0/XI0_7/d__12_ xsel_7_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_11 XI11_6/XI0/XI0_7/d__11_ xsel_7_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_10 XI11_6/XI0/XI0_7/d__10_ xsel_7_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_9 XI11_6/XI0/XI0_7/d__9_ xsel_7_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_8 XI11_6/XI0/XI0_7/d__8_ xsel_7_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_7 XI11_6/XI0/XI0_7/d__7_ xsel_7_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_6 XI11_6/XI0/XI0_7/d__6_ xsel_7_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_5 XI11_6/XI0/XI0_7/d__5_ xsel_7_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_4 XI11_6/XI0/XI0_7/d__4_ xsel_7_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_3 XI11_6/XI0/XI0_7/d__3_ xsel_7_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_2 XI11_6/XI0/XI0_7/d__2_ xsel_7_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_1 XI11_6/XI0/XI0_7/d__1_ xsel_7_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_0 XI11_6/XI0/XI0_7/d__0_ xsel_7_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_15 XI11_6/net21_0_ xsel_6_ XI11_6/XI0/XI0_6/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_14 XI11_6/net21_1_ xsel_6_ XI11_6/XI0/XI0_6/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_13 XI11_6/net21_2_ xsel_6_ XI11_6/XI0/XI0_6/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_12 XI11_6/net21_3_ xsel_6_ XI11_6/XI0/XI0_6/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_11 XI11_6/net21_4_ xsel_6_ XI11_6/XI0/XI0_6/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_10 XI11_6/net21_5_ xsel_6_ XI11_6/XI0/XI0_6/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_9 XI11_6/net21_6_ xsel_6_ XI11_6/XI0/XI0_6/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_8 XI11_6/net21_7_ xsel_6_ XI11_6/XI0/XI0_6/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_7 XI11_6/net21_8_ xsel_6_ XI11_6/XI0/XI0_6/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_6 XI11_6/net21_9_ xsel_6_ XI11_6/XI0/XI0_6/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_5 XI11_6/net21_10_ xsel_6_ XI11_6/XI0/XI0_6/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_4 XI11_6/net21_11_ xsel_6_ XI11_6/XI0/XI0_6/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_3 XI11_6/net21_12_ xsel_6_ XI11_6/XI0/XI0_6/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_2 XI11_6/net21_13_ xsel_6_ XI11_6/XI0/XI0_6/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_1 XI11_6/net21_14_ xsel_6_ XI11_6/XI0/XI0_6/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_0 XI11_6/net21_15_ xsel_6_ XI11_6/XI0/XI0_6/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_15 XI11_6/XI0/XI0_6/d__15_ xsel_6_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_14 XI11_6/XI0/XI0_6/d__14_ xsel_6_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_13 XI11_6/XI0/XI0_6/d__13_ xsel_6_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_12 XI11_6/XI0/XI0_6/d__12_ xsel_6_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_11 XI11_6/XI0/XI0_6/d__11_ xsel_6_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_10 XI11_6/XI0/XI0_6/d__10_ xsel_6_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_9 XI11_6/XI0/XI0_6/d__9_ xsel_6_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_8 XI11_6/XI0/XI0_6/d__8_ xsel_6_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_7 XI11_6/XI0/XI0_6/d__7_ xsel_6_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_6 XI11_6/XI0/XI0_6/d__6_ xsel_6_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_5 XI11_6/XI0/XI0_6/d__5_ xsel_6_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_4 XI11_6/XI0/XI0_6/d__4_ xsel_6_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_3 XI11_6/XI0/XI0_6/d__3_ xsel_6_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_2 XI11_6/XI0/XI0_6/d__2_ xsel_6_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_1 XI11_6/XI0/XI0_6/d__1_ xsel_6_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_0 XI11_6/XI0/XI0_6/d__0_ xsel_6_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_15 XI11_6/net21_0_ xsel_5_ XI11_6/XI0/XI0_5/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_14 XI11_6/net21_1_ xsel_5_ XI11_6/XI0/XI0_5/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_13 XI11_6/net21_2_ xsel_5_ XI11_6/XI0/XI0_5/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_12 XI11_6/net21_3_ xsel_5_ XI11_6/XI0/XI0_5/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_11 XI11_6/net21_4_ xsel_5_ XI11_6/XI0/XI0_5/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_10 XI11_6/net21_5_ xsel_5_ XI11_6/XI0/XI0_5/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_9 XI11_6/net21_6_ xsel_5_ XI11_6/XI0/XI0_5/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_8 XI11_6/net21_7_ xsel_5_ XI11_6/XI0/XI0_5/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_7 XI11_6/net21_8_ xsel_5_ XI11_6/XI0/XI0_5/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_6 XI11_6/net21_9_ xsel_5_ XI11_6/XI0/XI0_5/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_5 XI11_6/net21_10_ xsel_5_ XI11_6/XI0/XI0_5/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_4 XI11_6/net21_11_ xsel_5_ XI11_6/XI0/XI0_5/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_3 XI11_6/net21_12_ xsel_5_ XI11_6/XI0/XI0_5/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_2 XI11_6/net21_13_ xsel_5_ XI11_6/XI0/XI0_5/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_1 XI11_6/net21_14_ xsel_5_ XI11_6/XI0/XI0_5/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_0 XI11_6/net21_15_ xsel_5_ XI11_6/XI0/XI0_5/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_15 XI11_6/XI0/XI0_5/d__15_ xsel_5_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_14 XI11_6/XI0/XI0_5/d__14_ xsel_5_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_13 XI11_6/XI0/XI0_5/d__13_ xsel_5_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_12 XI11_6/XI0/XI0_5/d__12_ xsel_5_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_11 XI11_6/XI0/XI0_5/d__11_ xsel_5_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_10 XI11_6/XI0/XI0_5/d__10_ xsel_5_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_9 XI11_6/XI0/XI0_5/d__9_ xsel_5_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_8 XI11_6/XI0/XI0_5/d__8_ xsel_5_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_7 XI11_6/XI0/XI0_5/d__7_ xsel_5_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_6 XI11_6/XI0/XI0_5/d__6_ xsel_5_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_5 XI11_6/XI0/XI0_5/d__5_ xsel_5_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_4 XI11_6/XI0/XI0_5/d__4_ xsel_5_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_3 XI11_6/XI0/XI0_5/d__3_ xsel_5_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_2 XI11_6/XI0/XI0_5/d__2_ xsel_5_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_1 XI11_6/XI0/XI0_5/d__1_ xsel_5_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_0 XI11_6/XI0/XI0_5/d__0_ xsel_5_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_15 XI11_6/net21_0_ xsel_4_ XI11_6/XI0/XI0_4/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_14 XI11_6/net21_1_ xsel_4_ XI11_6/XI0/XI0_4/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_13 XI11_6/net21_2_ xsel_4_ XI11_6/XI0/XI0_4/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_12 XI11_6/net21_3_ xsel_4_ XI11_6/XI0/XI0_4/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_11 XI11_6/net21_4_ xsel_4_ XI11_6/XI0/XI0_4/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_10 XI11_6/net21_5_ xsel_4_ XI11_6/XI0/XI0_4/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_9 XI11_6/net21_6_ xsel_4_ XI11_6/XI0/XI0_4/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_8 XI11_6/net21_7_ xsel_4_ XI11_6/XI0/XI0_4/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_7 XI11_6/net21_8_ xsel_4_ XI11_6/XI0/XI0_4/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_6 XI11_6/net21_9_ xsel_4_ XI11_6/XI0/XI0_4/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_5 XI11_6/net21_10_ xsel_4_ XI11_6/XI0/XI0_4/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_4 XI11_6/net21_11_ xsel_4_ XI11_6/XI0/XI0_4/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_3 XI11_6/net21_12_ xsel_4_ XI11_6/XI0/XI0_4/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_2 XI11_6/net21_13_ xsel_4_ XI11_6/XI0/XI0_4/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_1 XI11_6/net21_14_ xsel_4_ XI11_6/XI0/XI0_4/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_0 XI11_6/net21_15_ xsel_4_ XI11_6/XI0/XI0_4/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_15 XI11_6/XI0/XI0_4/d__15_ xsel_4_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_14 XI11_6/XI0/XI0_4/d__14_ xsel_4_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_13 XI11_6/XI0/XI0_4/d__13_ xsel_4_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_12 XI11_6/XI0/XI0_4/d__12_ xsel_4_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_11 XI11_6/XI0/XI0_4/d__11_ xsel_4_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_10 XI11_6/XI0/XI0_4/d__10_ xsel_4_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_9 XI11_6/XI0/XI0_4/d__9_ xsel_4_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_8 XI11_6/XI0/XI0_4/d__8_ xsel_4_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_7 XI11_6/XI0/XI0_4/d__7_ xsel_4_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_6 XI11_6/XI0/XI0_4/d__6_ xsel_4_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_5 XI11_6/XI0/XI0_4/d__5_ xsel_4_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_4 XI11_6/XI0/XI0_4/d__4_ xsel_4_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_3 XI11_6/XI0/XI0_4/d__3_ xsel_4_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_2 XI11_6/XI0/XI0_4/d__2_ xsel_4_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_1 XI11_6/XI0/XI0_4/d__1_ xsel_4_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_0 XI11_6/XI0/XI0_4/d__0_ xsel_4_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_15 XI11_6/net21_0_ xsel_3_ XI11_6/XI0/XI0_3/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_14 XI11_6/net21_1_ xsel_3_ XI11_6/XI0/XI0_3/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_13 XI11_6/net21_2_ xsel_3_ XI11_6/XI0/XI0_3/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_12 XI11_6/net21_3_ xsel_3_ XI11_6/XI0/XI0_3/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_11 XI11_6/net21_4_ xsel_3_ XI11_6/XI0/XI0_3/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_10 XI11_6/net21_5_ xsel_3_ XI11_6/XI0/XI0_3/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_9 XI11_6/net21_6_ xsel_3_ XI11_6/XI0/XI0_3/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_8 XI11_6/net21_7_ xsel_3_ XI11_6/XI0/XI0_3/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_7 XI11_6/net21_8_ xsel_3_ XI11_6/XI0/XI0_3/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_6 XI11_6/net21_9_ xsel_3_ XI11_6/XI0/XI0_3/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_5 XI11_6/net21_10_ xsel_3_ XI11_6/XI0/XI0_3/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_4 XI11_6/net21_11_ xsel_3_ XI11_6/XI0/XI0_3/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_3 XI11_6/net21_12_ xsel_3_ XI11_6/XI0/XI0_3/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_2 XI11_6/net21_13_ xsel_3_ XI11_6/XI0/XI0_3/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_1 XI11_6/net21_14_ xsel_3_ XI11_6/XI0/XI0_3/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_0 XI11_6/net21_15_ xsel_3_ XI11_6/XI0/XI0_3/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_15 XI11_6/XI0/XI0_3/d__15_ xsel_3_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_14 XI11_6/XI0/XI0_3/d__14_ xsel_3_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_13 XI11_6/XI0/XI0_3/d__13_ xsel_3_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_12 XI11_6/XI0/XI0_3/d__12_ xsel_3_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_11 XI11_6/XI0/XI0_3/d__11_ xsel_3_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_10 XI11_6/XI0/XI0_3/d__10_ xsel_3_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_9 XI11_6/XI0/XI0_3/d__9_ xsel_3_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_8 XI11_6/XI0/XI0_3/d__8_ xsel_3_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_7 XI11_6/XI0/XI0_3/d__7_ xsel_3_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_6 XI11_6/XI0/XI0_3/d__6_ xsel_3_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_5 XI11_6/XI0/XI0_3/d__5_ xsel_3_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_4 XI11_6/XI0/XI0_3/d__4_ xsel_3_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_3 XI11_6/XI0/XI0_3/d__3_ xsel_3_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_2 XI11_6/XI0/XI0_3/d__2_ xsel_3_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_1 XI11_6/XI0/XI0_3/d__1_ xsel_3_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_0 XI11_6/XI0/XI0_3/d__0_ xsel_3_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_15 XI11_6/net21_0_ xsel_2_ XI11_6/XI0/XI0_2/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_14 XI11_6/net21_1_ xsel_2_ XI11_6/XI0/XI0_2/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_13 XI11_6/net21_2_ xsel_2_ XI11_6/XI0/XI0_2/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_12 XI11_6/net21_3_ xsel_2_ XI11_6/XI0/XI0_2/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_11 XI11_6/net21_4_ xsel_2_ XI11_6/XI0/XI0_2/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_10 XI11_6/net21_5_ xsel_2_ XI11_6/XI0/XI0_2/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_9 XI11_6/net21_6_ xsel_2_ XI11_6/XI0/XI0_2/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_8 XI11_6/net21_7_ xsel_2_ XI11_6/XI0/XI0_2/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_7 XI11_6/net21_8_ xsel_2_ XI11_6/XI0/XI0_2/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_6 XI11_6/net21_9_ xsel_2_ XI11_6/XI0/XI0_2/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_5 XI11_6/net21_10_ xsel_2_ XI11_6/XI0/XI0_2/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_4 XI11_6/net21_11_ xsel_2_ XI11_6/XI0/XI0_2/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_3 XI11_6/net21_12_ xsel_2_ XI11_6/XI0/XI0_2/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_2 XI11_6/net21_13_ xsel_2_ XI11_6/XI0/XI0_2/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_1 XI11_6/net21_14_ xsel_2_ XI11_6/XI0/XI0_2/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_0 XI11_6/net21_15_ xsel_2_ XI11_6/XI0/XI0_2/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_15 XI11_6/XI0/XI0_2/d__15_ xsel_2_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_14 XI11_6/XI0/XI0_2/d__14_ xsel_2_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_13 XI11_6/XI0/XI0_2/d__13_ xsel_2_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_12 XI11_6/XI0/XI0_2/d__12_ xsel_2_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_11 XI11_6/XI0/XI0_2/d__11_ xsel_2_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_10 XI11_6/XI0/XI0_2/d__10_ xsel_2_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_9 XI11_6/XI0/XI0_2/d__9_ xsel_2_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_8 XI11_6/XI0/XI0_2/d__8_ xsel_2_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_7 XI11_6/XI0/XI0_2/d__7_ xsel_2_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_6 XI11_6/XI0/XI0_2/d__6_ xsel_2_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_5 XI11_6/XI0/XI0_2/d__5_ xsel_2_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_4 XI11_6/XI0/XI0_2/d__4_ xsel_2_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_3 XI11_6/XI0/XI0_2/d__3_ xsel_2_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_2 XI11_6/XI0/XI0_2/d__2_ xsel_2_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_1 XI11_6/XI0/XI0_2/d__1_ xsel_2_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_0 XI11_6/XI0/XI0_2/d__0_ xsel_2_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_15 XI11_6/net21_0_ xsel_1_ XI11_6/XI0/XI0_1/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_14 XI11_6/net21_1_ xsel_1_ XI11_6/XI0/XI0_1/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_13 XI11_6/net21_2_ xsel_1_ XI11_6/XI0/XI0_1/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_12 XI11_6/net21_3_ xsel_1_ XI11_6/XI0/XI0_1/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_11 XI11_6/net21_4_ xsel_1_ XI11_6/XI0/XI0_1/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_10 XI11_6/net21_5_ xsel_1_ XI11_6/XI0/XI0_1/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_9 XI11_6/net21_6_ xsel_1_ XI11_6/XI0/XI0_1/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_8 XI11_6/net21_7_ xsel_1_ XI11_6/XI0/XI0_1/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_7 XI11_6/net21_8_ xsel_1_ XI11_6/XI0/XI0_1/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_6 XI11_6/net21_9_ xsel_1_ XI11_6/XI0/XI0_1/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_5 XI11_6/net21_10_ xsel_1_ XI11_6/XI0/XI0_1/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_4 XI11_6/net21_11_ xsel_1_ XI11_6/XI0/XI0_1/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_3 XI11_6/net21_12_ xsel_1_ XI11_6/XI0/XI0_1/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_2 XI11_6/net21_13_ xsel_1_ XI11_6/XI0/XI0_1/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_1 XI11_6/net21_14_ xsel_1_ XI11_6/XI0/XI0_1/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_0 XI11_6/net21_15_ xsel_1_ XI11_6/XI0/XI0_1/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_15 XI11_6/XI0/XI0_1/d__15_ xsel_1_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_14 XI11_6/XI0/XI0_1/d__14_ xsel_1_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_13 XI11_6/XI0/XI0_1/d__13_ xsel_1_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_12 XI11_6/XI0/XI0_1/d__12_ xsel_1_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_11 XI11_6/XI0/XI0_1/d__11_ xsel_1_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_10 XI11_6/XI0/XI0_1/d__10_ xsel_1_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_9 XI11_6/XI0/XI0_1/d__9_ xsel_1_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_8 XI11_6/XI0/XI0_1/d__8_ xsel_1_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_7 XI11_6/XI0/XI0_1/d__7_ xsel_1_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_6 XI11_6/XI0/XI0_1/d__6_ xsel_1_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_5 XI11_6/XI0/XI0_1/d__5_ xsel_1_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_4 XI11_6/XI0/XI0_1/d__4_ xsel_1_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_3 XI11_6/XI0/XI0_1/d__3_ xsel_1_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_2 XI11_6/XI0/XI0_1/d__2_ xsel_1_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_1 XI11_6/XI0/XI0_1/d__1_ xsel_1_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_0 XI11_6/XI0/XI0_1/d__0_ xsel_1_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_15 XI11_6/net21_0_ xsel_0_ XI11_6/XI0/XI0_0/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_14 XI11_6/net21_1_ xsel_0_ XI11_6/XI0/XI0_0/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_13 XI11_6/net21_2_ xsel_0_ XI11_6/XI0/XI0_0/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_12 XI11_6/net21_3_ xsel_0_ XI11_6/XI0/XI0_0/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_11 XI11_6/net21_4_ xsel_0_ XI11_6/XI0/XI0_0/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_10 XI11_6/net21_5_ xsel_0_ XI11_6/XI0/XI0_0/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_9 XI11_6/net21_6_ xsel_0_ XI11_6/XI0/XI0_0/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_8 XI11_6/net21_7_ xsel_0_ XI11_6/XI0/XI0_0/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_7 XI11_6/net21_8_ xsel_0_ XI11_6/XI0/XI0_0/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_6 XI11_6/net21_9_ xsel_0_ XI11_6/XI0/XI0_0/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_5 XI11_6/net21_10_ xsel_0_ XI11_6/XI0/XI0_0/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_4 XI11_6/net21_11_ xsel_0_ XI11_6/XI0/XI0_0/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_3 XI11_6/net21_12_ xsel_0_ XI11_6/XI0/XI0_0/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_2 XI11_6/net21_13_ xsel_0_ XI11_6/XI0/XI0_0/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_1 XI11_6/net21_14_ xsel_0_ XI11_6/XI0/XI0_0/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_0 XI11_6/net21_15_ xsel_0_ XI11_6/XI0/XI0_0/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_15 XI11_6/XI0/XI0_0/d__15_ xsel_0_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_14 XI11_6/XI0/XI0_0/d__14_ xsel_0_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_13 XI11_6/XI0/XI0_0/d__13_ xsel_0_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_12 XI11_6/XI0/XI0_0/d__12_ xsel_0_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_11 XI11_6/XI0/XI0_0/d__11_ xsel_0_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_10 XI11_6/XI0/XI0_0/d__10_ xsel_0_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_9 XI11_6/XI0/XI0_0/d__9_ xsel_0_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_8 XI11_6/XI0/XI0_0/d__8_ xsel_0_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_7 XI11_6/XI0/XI0_0/d__7_ xsel_0_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_6 XI11_6/XI0/XI0_0/d__6_ xsel_0_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_5 XI11_6/XI0/XI0_0/d__5_ xsel_0_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_4 XI11_6/XI0/XI0_0/d__4_ xsel_0_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_3 XI11_6/XI0/XI0_0/d__3_ xsel_0_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_2 XI11_6/XI0/XI0_0/d__2_ xsel_0_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_1 XI11_6/XI0/XI0_0/d__1_ xsel_0_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_0 XI11_6/XI0/XI0_0/d__0_ xsel_0_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI2/MN0_15 XI11_5/net21_0_ ysel_15_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_14 XI11_5/net21_1_ ysel_14_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_13 XI11_5/net21_2_ ysel_13_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_12 XI11_5/net21_3_ ysel_12_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_11 XI11_5/net21_4_ ysel_11_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_10 XI11_5/net21_5_ ysel_10_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_9 XI11_5/net21_6_ ysel_9_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_8 XI11_5/net21_7_ ysel_8_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_7 XI11_5/net21_8_ ysel_7_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_6 XI11_5/net21_9_ ysel_6_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_5 XI11_5/net21_10_ ysel_5_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_4 XI11_5/net21_11_ ysel_4_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_3 XI11_5/net21_12_ ysel_3_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_2 XI11_5/net21_13_ ysel_2_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_1 XI11_5/net21_14_ ysel_1_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_0 XI11_5/net21_15_ ysel_0_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_15 XI11_5/net20_0_ ysel_15_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_14 XI11_5/net20_1_ ysel_14_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_13 XI11_5/net20_2_ ysel_13_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_12 XI11_5/net20_3_ ysel_12_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_11 XI11_5/net20_4_ ysel_11_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_10 XI11_5/net20_5_ ysel_10_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_9 XI11_5/net20_6_ ysel_9_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_8 XI11_5/net20_7_ ysel_8_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_7 XI11_5/net20_8_ ysel_7_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_6 XI11_5/net20_9_ ysel_6_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_5 XI11_5/net20_10_ ysel_5_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_4 XI11_5/net20_11_ ysel_4_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_3 XI11_5/net20_12_ ysel_3_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_2 XI11_5/net20_13_ ysel_2_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_1 XI11_5/net20_14_ ysel_1_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_0 XI11_5/net20_15_ ysel_0_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI4/MN8 vdd XI11_5/XI4/net8 XI11_5/net12 vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_5/XI4/MP0 XI11_5/net9 XI11_5/XI4/net23 vdd vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_5/XI4/MP4 XI11_5/net12 XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI4/MP1 XI11_5/net9 XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI4/MP5 XI11_5/net12 XI11_5/preck XI11_5/net9 vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI4/MN7 vdd XI11_5/XI4/net090 DOUT_5_ vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_5/XI4/MP3 gnd XI11_5/XI4/net089 XI11_5/net12 gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_5/XI4/MN5 XI11_5/net9 XI11_5/XI4/net0103 gnd gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_5/XI4/MN4 XI11_5/XI4/data_out_ XI11_5/XI4/net32 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_5/XI4/MN0 XI11_5/XI4/data_out XI11_5/XI4/net52 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_5/XI4/MN9 gnd XI11_5/XI4/net0112 DOUT_5_ gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_5/XI1_15/MP2 XI11_5/net20_0_ XI11_5/preck XI11_5/net21_0_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_15/MP1 XI11_5/net20_0_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_15/MP0 XI11_5/net21_0_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_14/MP2 XI11_5/net20_1_ XI11_5/preck XI11_5/net21_1_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_14/MP1 XI11_5/net20_1_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_14/MP0 XI11_5/net21_1_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_13/MP2 XI11_5/net20_2_ XI11_5/preck XI11_5/net21_2_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_13/MP1 XI11_5/net20_2_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_13/MP0 XI11_5/net21_2_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_12/MP2 XI11_5/net20_3_ XI11_5/preck XI11_5/net21_3_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_12/MP1 XI11_5/net20_3_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_12/MP0 XI11_5/net21_3_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_11/MP2 XI11_5/net20_4_ XI11_5/preck XI11_5/net21_4_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_11/MP1 XI11_5/net20_4_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_11/MP0 XI11_5/net21_4_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_10/MP2 XI11_5/net20_5_ XI11_5/preck XI11_5/net21_5_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_10/MP1 XI11_5/net20_5_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_10/MP0 XI11_5/net21_5_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_9/MP2 XI11_5/net20_6_ XI11_5/preck XI11_5/net21_6_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_9/MP1 XI11_5/net20_6_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_9/MP0 XI11_5/net21_6_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_8/MP2 XI11_5/net20_7_ XI11_5/preck XI11_5/net21_7_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_8/MP1 XI11_5/net20_7_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_8/MP0 XI11_5/net21_7_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_7/MP2 XI11_5/net20_8_ XI11_5/preck XI11_5/net21_8_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_7/MP1 XI11_5/net20_8_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_7/MP0 XI11_5/net21_8_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_6/MP2 XI11_5/net20_9_ XI11_5/preck XI11_5/net21_9_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_6/MP1 XI11_5/net20_9_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_6/MP0 XI11_5/net21_9_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_5/MP2 XI11_5/net20_10_ XI11_5/preck XI11_5/net21_10_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_5/MP1 XI11_5/net20_10_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_5/MP0 XI11_5/net21_10_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_4/MP2 XI11_5/net20_11_ XI11_5/preck XI11_5/net21_11_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_4/MP1 XI11_5/net20_11_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_4/MP0 XI11_5/net21_11_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_3/MP2 XI11_5/net20_12_ XI11_5/preck XI11_5/net21_12_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_3/MP1 XI11_5/net20_12_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_3/MP0 XI11_5/net21_12_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_2/MP2 XI11_5/net20_13_ XI11_5/preck XI11_5/net21_13_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_2/MP1 XI11_5/net20_13_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_2/MP0 XI11_5/net21_13_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_1/MP2 XI11_5/net20_14_ XI11_5/preck XI11_5/net21_14_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_1/MP1 XI11_5/net20_14_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_1/MP0 XI11_5/net21_14_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_0/MP2 XI11_5/net20_15_ XI11_5/preck XI11_5/net21_15_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_0/MP1 XI11_5/net20_15_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_0/MP0 XI11_5/net21_15_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI0/MN0_15 gnd gnd XI11_5/net21_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_14 gnd gnd XI11_5/net21_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_13 gnd gnd XI11_5/net21_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_12 gnd gnd XI11_5/net21_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_11 gnd gnd XI11_5/net21_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_10 gnd gnd XI11_5/net21_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_9 gnd gnd XI11_5/net21_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_8 gnd gnd XI11_5/net21_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_7 gnd gnd XI11_5/net21_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_6 gnd gnd XI11_5/net21_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_5 gnd gnd XI11_5/net21_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_4 gnd gnd XI11_5/net21_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_3 gnd gnd XI11_5/net21_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_2 gnd gnd XI11_5/net21_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_1 gnd gnd XI11_5/net21_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_0 gnd gnd XI11_5/net21_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_15 gnd gnd XI11_5/net20_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_14 gnd gnd XI11_5/net20_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_13 gnd gnd XI11_5/net20_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_12 gnd gnd XI11_5/net20_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_11 gnd gnd XI11_5/net20_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_10 gnd gnd XI11_5/net20_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_9 gnd gnd XI11_5/net20_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_8 gnd gnd XI11_5/net20_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_7 gnd gnd XI11_5/net20_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_6 gnd gnd XI11_5/net20_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_5 gnd gnd XI11_5/net20_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_4 gnd gnd XI11_5/net20_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_3 gnd gnd XI11_5/net20_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_2 gnd gnd XI11_5/net20_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_1 gnd gnd XI11_5/net20_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_0 gnd gnd XI11_5/net20_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_15 XI11_5/net21_0_ xsel_63_ XI11_5/XI0/XI0_63/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_14 XI11_5/net21_1_ xsel_63_ XI11_5/XI0/XI0_63/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_13 XI11_5/net21_2_ xsel_63_ XI11_5/XI0/XI0_63/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_12 XI11_5/net21_3_ xsel_63_ XI11_5/XI0/XI0_63/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_11 XI11_5/net21_4_ xsel_63_ XI11_5/XI0/XI0_63/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_10 XI11_5/net21_5_ xsel_63_ XI11_5/XI0/XI0_63/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_9 XI11_5/net21_6_ xsel_63_ XI11_5/XI0/XI0_63/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_8 XI11_5/net21_7_ xsel_63_ XI11_5/XI0/XI0_63/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_7 XI11_5/net21_8_ xsel_63_ XI11_5/XI0/XI0_63/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_6 XI11_5/net21_9_ xsel_63_ XI11_5/XI0/XI0_63/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_5 XI11_5/net21_10_ xsel_63_ XI11_5/XI0/XI0_63/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_4 XI11_5/net21_11_ xsel_63_ XI11_5/XI0/XI0_63/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_3 XI11_5/net21_12_ xsel_63_ XI11_5/XI0/XI0_63/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_2 XI11_5/net21_13_ xsel_63_ XI11_5/XI0/XI0_63/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_1 XI11_5/net21_14_ xsel_63_ XI11_5/XI0/XI0_63/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_0 XI11_5/net21_15_ xsel_63_ XI11_5/XI0/XI0_63/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_15 XI11_5/XI0/XI0_63/d__15_ xsel_63_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_14 XI11_5/XI0/XI0_63/d__14_ xsel_63_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_13 XI11_5/XI0/XI0_63/d__13_ xsel_63_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_12 XI11_5/XI0/XI0_63/d__12_ xsel_63_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_11 XI11_5/XI0/XI0_63/d__11_ xsel_63_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_10 XI11_5/XI0/XI0_63/d__10_ xsel_63_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_9 XI11_5/XI0/XI0_63/d__9_ xsel_63_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_8 XI11_5/XI0/XI0_63/d__8_ xsel_63_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_7 XI11_5/XI0/XI0_63/d__7_ xsel_63_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_6 XI11_5/XI0/XI0_63/d__6_ xsel_63_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_5 XI11_5/XI0/XI0_63/d__5_ xsel_63_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_4 XI11_5/XI0/XI0_63/d__4_ xsel_63_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_3 XI11_5/XI0/XI0_63/d__3_ xsel_63_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_2 XI11_5/XI0/XI0_63/d__2_ xsel_63_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_1 XI11_5/XI0/XI0_63/d__1_ xsel_63_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_0 XI11_5/XI0/XI0_63/d__0_ xsel_63_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_15 XI11_5/net21_0_ xsel_62_ XI11_5/XI0/XI0_62/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_14 XI11_5/net21_1_ xsel_62_ XI11_5/XI0/XI0_62/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_13 XI11_5/net21_2_ xsel_62_ XI11_5/XI0/XI0_62/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_12 XI11_5/net21_3_ xsel_62_ XI11_5/XI0/XI0_62/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_11 XI11_5/net21_4_ xsel_62_ XI11_5/XI0/XI0_62/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_10 XI11_5/net21_5_ xsel_62_ XI11_5/XI0/XI0_62/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_9 XI11_5/net21_6_ xsel_62_ XI11_5/XI0/XI0_62/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_8 XI11_5/net21_7_ xsel_62_ XI11_5/XI0/XI0_62/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_7 XI11_5/net21_8_ xsel_62_ XI11_5/XI0/XI0_62/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_6 XI11_5/net21_9_ xsel_62_ XI11_5/XI0/XI0_62/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_5 XI11_5/net21_10_ xsel_62_ XI11_5/XI0/XI0_62/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_4 XI11_5/net21_11_ xsel_62_ XI11_5/XI0/XI0_62/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_3 XI11_5/net21_12_ xsel_62_ XI11_5/XI0/XI0_62/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_2 XI11_5/net21_13_ xsel_62_ XI11_5/XI0/XI0_62/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_1 XI11_5/net21_14_ xsel_62_ XI11_5/XI0/XI0_62/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_0 XI11_5/net21_15_ xsel_62_ XI11_5/XI0/XI0_62/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_15 XI11_5/XI0/XI0_62/d__15_ xsel_62_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_14 XI11_5/XI0/XI0_62/d__14_ xsel_62_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_13 XI11_5/XI0/XI0_62/d__13_ xsel_62_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_12 XI11_5/XI0/XI0_62/d__12_ xsel_62_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_11 XI11_5/XI0/XI0_62/d__11_ xsel_62_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_10 XI11_5/XI0/XI0_62/d__10_ xsel_62_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_9 XI11_5/XI0/XI0_62/d__9_ xsel_62_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_8 XI11_5/XI0/XI0_62/d__8_ xsel_62_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_7 XI11_5/XI0/XI0_62/d__7_ xsel_62_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_6 XI11_5/XI0/XI0_62/d__6_ xsel_62_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_5 XI11_5/XI0/XI0_62/d__5_ xsel_62_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_4 XI11_5/XI0/XI0_62/d__4_ xsel_62_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_3 XI11_5/XI0/XI0_62/d__3_ xsel_62_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_2 XI11_5/XI0/XI0_62/d__2_ xsel_62_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_1 XI11_5/XI0/XI0_62/d__1_ xsel_62_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_0 XI11_5/XI0/XI0_62/d__0_ xsel_62_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_15 XI11_5/net21_0_ xsel_61_ XI11_5/XI0/XI0_61/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_14 XI11_5/net21_1_ xsel_61_ XI11_5/XI0/XI0_61/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_13 XI11_5/net21_2_ xsel_61_ XI11_5/XI0/XI0_61/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_12 XI11_5/net21_3_ xsel_61_ XI11_5/XI0/XI0_61/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_11 XI11_5/net21_4_ xsel_61_ XI11_5/XI0/XI0_61/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_10 XI11_5/net21_5_ xsel_61_ XI11_5/XI0/XI0_61/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_9 XI11_5/net21_6_ xsel_61_ XI11_5/XI0/XI0_61/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_8 XI11_5/net21_7_ xsel_61_ XI11_5/XI0/XI0_61/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_7 XI11_5/net21_8_ xsel_61_ XI11_5/XI0/XI0_61/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_6 XI11_5/net21_9_ xsel_61_ XI11_5/XI0/XI0_61/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_5 XI11_5/net21_10_ xsel_61_ XI11_5/XI0/XI0_61/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_4 XI11_5/net21_11_ xsel_61_ XI11_5/XI0/XI0_61/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_3 XI11_5/net21_12_ xsel_61_ XI11_5/XI0/XI0_61/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_2 XI11_5/net21_13_ xsel_61_ XI11_5/XI0/XI0_61/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_1 XI11_5/net21_14_ xsel_61_ XI11_5/XI0/XI0_61/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_0 XI11_5/net21_15_ xsel_61_ XI11_5/XI0/XI0_61/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_15 XI11_5/XI0/XI0_61/d__15_ xsel_61_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_14 XI11_5/XI0/XI0_61/d__14_ xsel_61_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_13 XI11_5/XI0/XI0_61/d__13_ xsel_61_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_12 XI11_5/XI0/XI0_61/d__12_ xsel_61_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_11 XI11_5/XI0/XI0_61/d__11_ xsel_61_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_10 XI11_5/XI0/XI0_61/d__10_ xsel_61_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_9 XI11_5/XI0/XI0_61/d__9_ xsel_61_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_8 XI11_5/XI0/XI0_61/d__8_ xsel_61_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_7 XI11_5/XI0/XI0_61/d__7_ xsel_61_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_6 XI11_5/XI0/XI0_61/d__6_ xsel_61_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_5 XI11_5/XI0/XI0_61/d__5_ xsel_61_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_4 XI11_5/XI0/XI0_61/d__4_ xsel_61_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_3 XI11_5/XI0/XI0_61/d__3_ xsel_61_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_2 XI11_5/XI0/XI0_61/d__2_ xsel_61_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_1 XI11_5/XI0/XI0_61/d__1_ xsel_61_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_0 XI11_5/XI0/XI0_61/d__0_ xsel_61_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_15 XI11_5/net21_0_ xsel_60_ XI11_5/XI0/XI0_60/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_14 XI11_5/net21_1_ xsel_60_ XI11_5/XI0/XI0_60/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_13 XI11_5/net21_2_ xsel_60_ XI11_5/XI0/XI0_60/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_12 XI11_5/net21_3_ xsel_60_ XI11_5/XI0/XI0_60/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_11 XI11_5/net21_4_ xsel_60_ XI11_5/XI0/XI0_60/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_10 XI11_5/net21_5_ xsel_60_ XI11_5/XI0/XI0_60/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_9 XI11_5/net21_6_ xsel_60_ XI11_5/XI0/XI0_60/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_8 XI11_5/net21_7_ xsel_60_ XI11_5/XI0/XI0_60/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_7 XI11_5/net21_8_ xsel_60_ XI11_5/XI0/XI0_60/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_6 XI11_5/net21_9_ xsel_60_ XI11_5/XI0/XI0_60/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_5 XI11_5/net21_10_ xsel_60_ XI11_5/XI0/XI0_60/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_4 XI11_5/net21_11_ xsel_60_ XI11_5/XI0/XI0_60/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_3 XI11_5/net21_12_ xsel_60_ XI11_5/XI0/XI0_60/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_2 XI11_5/net21_13_ xsel_60_ XI11_5/XI0/XI0_60/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_1 XI11_5/net21_14_ xsel_60_ XI11_5/XI0/XI0_60/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_0 XI11_5/net21_15_ xsel_60_ XI11_5/XI0/XI0_60/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_15 XI11_5/XI0/XI0_60/d__15_ xsel_60_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_14 XI11_5/XI0/XI0_60/d__14_ xsel_60_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_13 XI11_5/XI0/XI0_60/d__13_ xsel_60_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_12 XI11_5/XI0/XI0_60/d__12_ xsel_60_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_11 XI11_5/XI0/XI0_60/d__11_ xsel_60_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_10 XI11_5/XI0/XI0_60/d__10_ xsel_60_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_9 XI11_5/XI0/XI0_60/d__9_ xsel_60_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_8 XI11_5/XI0/XI0_60/d__8_ xsel_60_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_7 XI11_5/XI0/XI0_60/d__7_ xsel_60_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_6 XI11_5/XI0/XI0_60/d__6_ xsel_60_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_5 XI11_5/XI0/XI0_60/d__5_ xsel_60_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_4 XI11_5/XI0/XI0_60/d__4_ xsel_60_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_3 XI11_5/XI0/XI0_60/d__3_ xsel_60_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_2 XI11_5/XI0/XI0_60/d__2_ xsel_60_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_1 XI11_5/XI0/XI0_60/d__1_ xsel_60_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_0 XI11_5/XI0/XI0_60/d__0_ xsel_60_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_15 XI11_5/net21_0_ xsel_59_ XI11_5/XI0/XI0_59/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_14 XI11_5/net21_1_ xsel_59_ XI11_5/XI0/XI0_59/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_13 XI11_5/net21_2_ xsel_59_ XI11_5/XI0/XI0_59/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_12 XI11_5/net21_3_ xsel_59_ XI11_5/XI0/XI0_59/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_11 XI11_5/net21_4_ xsel_59_ XI11_5/XI0/XI0_59/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_10 XI11_5/net21_5_ xsel_59_ XI11_5/XI0/XI0_59/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_9 XI11_5/net21_6_ xsel_59_ XI11_5/XI0/XI0_59/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_8 XI11_5/net21_7_ xsel_59_ XI11_5/XI0/XI0_59/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_7 XI11_5/net21_8_ xsel_59_ XI11_5/XI0/XI0_59/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_6 XI11_5/net21_9_ xsel_59_ XI11_5/XI0/XI0_59/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_5 XI11_5/net21_10_ xsel_59_ XI11_5/XI0/XI0_59/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_4 XI11_5/net21_11_ xsel_59_ XI11_5/XI0/XI0_59/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_3 XI11_5/net21_12_ xsel_59_ XI11_5/XI0/XI0_59/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_2 XI11_5/net21_13_ xsel_59_ XI11_5/XI0/XI0_59/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_1 XI11_5/net21_14_ xsel_59_ XI11_5/XI0/XI0_59/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_0 XI11_5/net21_15_ xsel_59_ XI11_5/XI0/XI0_59/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_15 XI11_5/XI0/XI0_59/d__15_ xsel_59_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_14 XI11_5/XI0/XI0_59/d__14_ xsel_59_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_13 XI11_5/XI0/XI0_59/d__13_ xsel_59_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_12 XI11_5/XI0/XI0_59/d__12_ xsel_59_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_11 XI11_5/XI0/XI0_59/d__11_ xsel_59_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_10 XI11_5/XI0/XI0_59/d__10_ xsel_59_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_9 XI11_5/XI0/XI0_59/d__9_ xsel_59_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_8 XI11_5/XI0/XI0_59/d__8_ xsel_59_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_7 XI11_5/XI0/XI0_59/d__7_ xsel_59_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_6 XI11_5/XI0/XI0_59/d__6_ xsel_59_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_5 XI11_5/XI0/XI0_59/d__5_ xsel_59_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_4 XI11_5/XI0/XI0_59/d__4_ xsel_59_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_3 XI11_5/XI0/XI0_59/d__3_ xsel_59_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_2 XI11_5/XI0/XI0_59/d__2_ xsel_59_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_1 XI11_5/XI0/XI0_59/d__1_ xsel_59_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_0 XI11_5/XI0/XI0_59/d__0_ xsel_59_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_15 XI11_5/net21_0_ xsel_58_ XI11_5/XI0/XI0_58/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_14 XI11_5/net21_1_ xsel_58_ XI11_5/XI0/XI0_58/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_13 XI11_5/net21_2_ xsel_58_ XI11_5/XI0/XI0_58/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_12 XI11_5/net21_3_ xsel_58_ XI11_5/XI0/XI0_58/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_11 XI11_5/net21_4_ xsel_58_ XI11_5/XI0/XI0_58/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_10 XI11_5/net21_5_ xsel_58_ XI11_5/XI0/XI0_58/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_9 XI11_5/net21_6_ xsel_58_ XI11_5/XI0/XI0_58/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_8 XI11_5/net21_7_ xsel_58_ XI11_5/XI0/XI0_58/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_7 XI11_5/net21_8_ xsel_58_ XI11_5/XI0/XI0_58/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_6 XI11_5/net21_9_ xsel_58_ XI11_5/XI0/XI0_58/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_5 XI11_5/net21_10_ xsel_58_ XI11_5/XI0/XI0_58/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_4 XI11_5/net21_11_ xsel_58_ XI11_5/XI0/XI0_58/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_3 XI11_5/net21_12_ xsel_58_ XI11_5/XI0/XI0_58/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_2 XI11_5/net21_13_ xsel_58_ XI11_5/XI0/XI0_58/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_1 XI11_5/net21_14_ xsel_58_ XI11_5/XI0/XI0_58/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_0 XI11_5/net21_15_ xsel_58_ XI11_5/XI0/XI0_58/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_15 XI11_5/XI0/XI0_58/d__15_ xsel_58_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_14 XI11_5/XI0/XI0_58/d__14_ xsel_58_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_13 XI11_5/XI0/XI0_58/d__13_ xsel_58_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_12 XI11_5/XI0/XI0_58/d__12_ xsel_58_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_11 XI11_5/XI0/XI0_58/d__11_ xsel_58_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_10 XI11_5/XI0/XI0_58/d__10_ xsel_58_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_9 XI11_5/XI0/XI0_58/d__9_ xsel_58_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_8 XI11_5/XI0/XI0_58/d__8_ xsel_58_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_7 XI11_5/XI0/XI0_58/d__7_ xsel_58_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_6 XI11_5/XI0/XI0_58/d__6_ xsel_58_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_5 XI11_5/XI0/XI0_58/d__5_ xsel_58_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_4 XI11_5/XI0/XI0_58/d__4_ xsel_58_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_3 XI11_5/XI0/XI0_58/d__3_ xsel_58_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_2 XI11_5/XI0/XI0_58/d__2_ xsel_58_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_1 XI11_5/XI0/XI0_58/d__1_ xsel_58_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_0 XI11_5/XI0/XI0_58/d__0_ xsel_58_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_15 XI11_5/net21_0_ xsel_57_ XI11_5/XI0/XI0_57/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_14 XI11_5/net21_1_ xsel_57_ XI11_5/XI0/XI0_57/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_13 XI11_5/net21_2_ xsel_57_ XI11_5/XI0/XI0_57/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_12 XI11_5/net21_3_ xsel_57_ XI11_5/XI0/XI0_57/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_11 XI11_5/net21_4_ xsel_57_ XI11_5/XI0/XI0_57/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_10 XI11_5/net21_5_ xsel_57_ XI11_5/XI0/XI0_57/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_9 XI11_5/net21_6_ xsel_57_ XI11_5/XI0/XI0_57/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_8 XI11_5/net21_7_ xsel_57_ XI11_5/XI0/XI0_57/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_7 XI11_5/net21_8_ xsel_57_ XI11_5/XI0/XI0_57/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_6 XI11_5/net21_9_ xsel_57_ XI11_5/XI0/XI0_57/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_5 XI11_5/net21_10_ xsel_57_ XI11_5/XI0/XI0_57/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_4 XI11_5/net21_11_ xsel_57_ XI11_5/XI0/XI0_57/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_3 XI11_5/net21_12_ xsel_57_ XI11_5/XI0/XI0_57/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_2 XI11_5/net21_13_ xsel_57_ XI11_5/XI0/XI0_57/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_1 XI11_5/net21_14_ xsel_57_ XI11_5/XI0/XI0_57/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_0 XI11_5/net21_15_ xsel_57_ XI11_5/XI0/XI0_57/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_15 XI11_5/XI0/XI0_57/d__15_ xsel_57_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_14 XI11_5/XI0/XI0_57/d__14_ xsel_57_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_13 XI11_5/XI0/XI0_57/d__13_ xsel_57_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_12 XI11_5/XI0/XI0_57/d__12_ xsel_57_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_11 XI11_5/XI0/XI0_57/d__11_ xsel_57_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_10 XI11_5/XI0/XI0_57/d__10_ xsel_57_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_9 XI11_5/XI0/XI0_57/d__9_ xsel_57_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_8 XI11_5/XI0/XI0_57/d__8_ xsel_57_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_7 XI11_5/XI0/XI0_57/d__7_ xsel_57_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_6 XI11_5/XI0/XI0_57/d__6_ xsel_57_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_5 XI11_5/XI0/XI0_57/d__5_ xsel_57_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_4 XI11_5/XI0/XI0_57/d__4_ xsel_57_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_3 XI11_5/XI0/XI0_57/d__3_ xsel_57_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_2 XI11_5/XI0/XI0_57/d__2_ xsel_57_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_1 XI11_5/XI0/XI0_57/d__1_ xsel_57_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_0 XI11_5/XI0/XI0_57/d__0_ xsel_57_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_15 XI11_5/net21_0_ xsel_56_ XI11_5/XI0/XI0_56/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_14 XI11_5/net21_1_ xsel_56_ XI11_5/XI0/XI0_56/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_13 XI11_5/net21_2_ xsel_56_ XI11_5/XI0/XI0_56/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_12 XI11_5/net21_3_ xsel_56_ XI11_5/XI0/XI0_56/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_11 XI11_5/net21_4_ xsel_56_ XI11_5/XI0/XI0_56/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_10 XI11_5/net21_5_ xsel_56_ XI11_5/XI0/XI0_56/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_9 XI11_5/net21_6_ xsel_56_ XI11_5/XI0/XI0_56/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_8 XI11_5/net21_7_ xsel_56_ XI11_5/XI0/XI0_56/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_7 XI11_5/net21_8_ xsel_56_ XI11_5/XI0/XI0_56/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_6 XI11_5/net21_9_ xsel_56_ XI11_5/XI0/XI0_56/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_5 XI11_5/net21_10_ xsel_56_ XI11_5/XI0/XI0_56/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_4 XI11_5/net21_11_ xsel_56_ XI11_5/XI0/XI0_56/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_3 XI11_5/net21_12_ xsel_56_ XI11_5/XI0/XI0_56/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_2 XI11_5/net21_13_ xsel_56_ XI11_5/XI0/XI0_56/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_1 XI11_5/net21_14_ xsel_56_ XI11_5/XI0/XI0_56/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_0 XI11_5/net21_15_ xsel_56_ XI11_5/XI0/XI0_56/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_15 XI11_5/XI0/XI0_56/d__15_ xsel_56_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_14 XI11_5/XI0/XI0_56/d__14_ xsel_56_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_13 XI11_5/XI0/XI0_56/d__13_ xsel_56_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_12 XI11_5/XI0/XI0_56/d__12_ xsel_56_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_11 XI11_5/XI0/XI0_56/d__11_ xsel_56_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_10 XI11_5/XI0/XI0_56/d__10_ xsel_56_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_9 XI11_5/XI0/XI0_56/d__9_ xsel_56_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_8 XI11_5/XI0/XI0_56/d__8_ xsel_56_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_7 XI11_5/XI0/XI0_56/d__7_ xsel_56_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_6 XI11_5/XI0/XI0_56/d__6_ xsel_56_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_5 XI11_5/XI0/XI0_56/d__5_ xsel_56_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_4 XI11_5/XI0/XI0_56/d__4_ xsel_56_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_3 XI11_5/XI0/XI0_56/d__3_ xsel_56_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_2 XI11_5/XI0/XI0_56/d__2_ xsel_56_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_1 XI11_5/XI0/XI0_56/d__1_ xsel_56_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_0 XI11_5/XI0/XI0_56/d__0_ xsel_56_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_15 XI11_5/net21_0_ xsel_55_ XI11_5/XI0/XI0_55/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_14 XI11_5/net21_1_ xsel_55_ XI11_5/XI0/XI0_55/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_13 XI11_5/net21_2_ xsel_55_ XI11_5/XI0/XI0_55/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_12 XI11_5/net21_3_ xsel_55_ XI11_5/XI0/XI0_55/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_11 XI11_5/net21_4_ xsel_55_ XI11_5/XI0/XI0_55/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_10 XI11_5/net21_5_ xsel_55_ XI11_5/XI0/XI0_55/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_9 XI11_5/net21_6_ xsel_55_ XI11_5/XI0/XI0_55/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_8 XI11_5/net21_7_ xsel_55_ XI11_5/XI0/XI0_55/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_7 XI11_5/net21_8_ xsel_55_ XI11_5/XI0/XI0_55/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_6 XI11_5/net21_9_ xsel_55_ XI11_5/XI0/XI0_55/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_5 XI11_5/net21_10_ xsel_55_ XI11_5/XI0/XI0_55/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_4 XI11_5/net21_11_ xsel_55_ XI11_5/XI0/XI0_55/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_3 XI11_5/net21_12_ xsel_55_ XI11_5/XI0/XI0_55/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_2 XI11_5/net21_13_ xsel_55_ XI11_5/XI0/XI0_55/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_1 XI11_5/net21_14_ xsel_55_ XI11_5/XI0/XI0_55/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_0 XI11_5/net21_15_ xsel_55_ XI11_5/XI0/XI0_55/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_15 XI11_5/XI0/XI0_55/d__15_ xsel_55_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_14 XI11_5/XI0/XI0_55/d__14_ xsel_55_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_13 XI11_5/XI0/XI0_55/d__13_ xsel_55_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_12 XI11_5/XI0/XI0_55/d__12_ xsel_55_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_11 XI11_5/XI0/XI0_55/d__11_ xsel_55_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_10 XI11_5/XI0/XI0_55/d__10_ xsel_55_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_9 XI11_5/XI0/XI0_55/d__9_ xsel_55_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_8 XI11_5/XI0/XI0_55/d__8_ xsel_55_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_7 XI11_5/XI0/XI0_55/d__7_ xsel_55_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_6 XI11_5/XI0/XI0_55/d__6_ xsel_55_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_5 XI11_5/XI0/XI0_55/d__5_ xsel_55_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_4 XI11_5/XI0/XI0_55/d__4_ xsel_55_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_3 XI11_5/XI0/XI0_55/d__3_ xsel_55_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_2 XI11_5/XI0/XI0_55/d__2_ xsel_55_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_1 XI11_5/XI0/XI0_55/d__1_ xsel_55_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_0 XI11_5/XI0/XI0_55/d__0_ xsel_55_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_15 XI11_5/net21_0_ xsel_54_ XI11_5/XI0/XI0_54/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_14 XI11_5/net21_1_ xsel_54_ XI11_5/XI0/XI0_54/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_13 XI11_5/net21_2_ xsel_54_ XI11_5/XI0/XI0_54/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_12 XI11_5/net21_3_ xsel_54_ XI11_5/XI0/XI0_54/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_11 XI11_5/net21_4_ xsel_54_ XI11_5/XI0/XI0_54/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_10 XI11_5/net21_5_ xsel_54_ XI11_5/XI0/XI0_54/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_9 XI11_5/net21_6_ xsel_54_ XI11_5/XI0/XI0_54/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_8 XI11_5/net21_7_ xsel_54_ XI11_5/XI0/XI0_54/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_7 XI11_5/net21_8_ xsel_54_ XI11_5/XI0/XI0_54/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_6 XI11_5/net21_9_ xsel_54_ XI11_5/XI0/XI0_54/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_5 XI11_5/net21_10_ xsel_54_ XI11_5/XI0/XI0_54/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_4 XI11_5/net21_11_ xsel_54_ XI11_5/XI0/XI0_54/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_3 XI11_5/net21_12_ xsel_54_ XI11_5/XI0/XI0_54/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_2 XI11_5/net21_13_ xsel_54_ XI11_5/XI0/XI0_54/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_1 XI11_5/net21_14_ xsel_54_ XI11_5/XI0/XI0_54/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_0 XI11_5/net21_15_ xsel_54_ XI11_5/XI0/XI0_54/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_15 XI11_5/XI0/XI0_54/d__15_ xsel_54_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_14 XI11_5/XI0/XI0_54/d__14_ xsel_54_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_13 XI11_5/XI0/XI0_54/d__13_ xsel_54_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_12 XI11_5/XI0/XI0_54/d__12_ xsel_54_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_11 XI11_5/XI0/XI0_54/d__11_ xsel_54_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_10 XI11_5/XI0/XI0_54/d__10_ xsel_54_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_9 XI11_5/XI0/XI0_54/d__9_ xsel_54_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_8 XI11_5/XI0/XI0_54/d__8_ xsel_54_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_7 XI11_5/XI0/XI0_54/d__7_ xsel_54_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_6 XI11_5/XI0/XI0_54/d__6_ xsel_54_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_5 XI11_5/XI0/XI0_54/d__5_ xsel_54_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_4 XI11_5/XI0/XI0_54/d__4_ xsel_54_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_3 XI11_5/XI0/XI0_54/d__3_ xsel_54_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_2 XI11_5/XI0/XI0_54/d__2_ xsel_54_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_1 XI11_5/XI0/XI0_54/d__1_ xsel_54_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_0 XI11_5/XI0/XI0_54/d__0_ xsel_54_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_15 XI11_5/net21_0_ xsel_53_ XI11_5/XI0/XI0_53/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_14 XI11_5/net21_1_ xsel_53_ XI11_5/XI0/XI0_53/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_13 XI11_5/net21_2_ xsel_53_ XI11_5/XI0/XI0_53/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_12 XI11_5/net21_3_ xsel_53_ XI11_5/XI0/XI0_53/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_11 XI11_5/net21_4_ xsel_53_ XI11_5/XI0/XI0_53/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_10 XI11_5/net21_5_ xsel_53_ XI11_5/XI0/XI0_53/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_9 XI11_5/net21_6_ xsel_53_ XI11_5/XI0/XI0_53/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_8 XI11_5/net21_7_ xsel_53_ XI11_5/XI0/XI0_53/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_7 XI11_5/net21_8_ xsel_53_ XI11_5/XI0/XI0_53/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_6 XI11_5/net21_9_ xsel_53_ XI11_5/XI0/XI0_53/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_5 XI11_5/net21_10_ xsel_53_ XI11_5/XI0/XI0_53/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_4 XI11_5/net21_11_ xsel_53_ XI11_5/XI0/XI0_53/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_3 XI11_5/net21_12_ xsel_53_ XI11_5/XI0/XI0_53/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_2 XI11_5/net21_13_ xsel_53_ XI11_5/XI0/XI0_53/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_1 XI11_5/net21_14_ xsel_53_ XI11_5/XI0/XI0_53/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_0 XI11_5/net21_15_ xsel_53_ XI11_5/XI0/XI0_53/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_15 XI11_5/XI0/XI0_53/d__15_ xsel_53_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_14 XI11_5/XI0/XI0_53/d__14_ xsel_53_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_13 XI11_5/XI0/XI0_53/d__13_ xsel_53_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_12 XI11_5/XI0/XI0_53/d__12_ xsel_53_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_11 XI11_5/XI0/XI0_53/d__11_ xsel_53_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_10 XI11_5/XI0/XI0_53/d__10_ xsel_53_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_9 XI11_5/XI0/XI0_53/d__9_ xsel_53_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_8 XI11_5/XI0/XI0_53/d__8_ xsel_53_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_7 XI11_5/XI0/XI0_53/d__7_ xsel_53_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_6 XI11_5/XI0/XI0_53/d__6_ xsel_53_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_5 XI11_5/XI0/XI0_53/d__5_ xsel_53_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_4 XI11_5/XI0/XI0_53/d__4_ xsel_53_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_3 XI11_5/XI0/XI0_53/d__3_ xsel_53_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_2 XI11_5/XI0/XI0_53/d__2_ xsel_53_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_1 XI11_5/XI0/XI0_53/d__1_ xsel_53_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_0 XI11_5/XI0/XI0_53/d__0_ xsel_53_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_15 XI11_5/net21_0_ xsel_52_ XI11_5/XI0/XI0_52/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_14 XI11_5/net21_1_ xsel_52_ XI11_5/XI0/XI0_52/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_13 XI11_5/net21_2_ xsel_52_ XI11_5/XI0/XI0_52/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_12 XI11_5/net21_3_ xsel_52_ XI11_5/XI0/XI0_52/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_11 XI11_5/net21_4_ xsel_52_ XI11_5/XI0/XI0_52/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_10 XI11_5/net21_5_ xsel_52_ XI11_5/XI0/XI0_52/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_9 XI11_5/net21_6_ xsel_52_ XI11_5/XI0/XI0_52/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_8 XI11_5/net21_7_ xsel_52_ XI11_5/XI0/XI0_52/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_7 XI11_5/net21_8_ xsel_52_ XI11_5/XI0/XI0_52/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_6 XI11_5/net21_9_ xsel_52_ XI11_5/XI0/XI0_52/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_5 XI11_5/net21_10_ xsel_52_ XI11_5/XI0/XI0_52/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_4 XI11_5/net21_11_ xsel_52_ XI11_5/XI0/XI0_52/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_3 XI11_5/net21_12_ xsel_52_ XI11_5/XI0/XI0_52/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_2 XI11_5/net21_13_ xsel_52_ XI11_5/XI0/XI0_52/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_1 XI11_5/net21_14_ xsel_52_ XI11_5/XI0/XI0_52/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_0 XI11_5/net21_15_ xsel_52_ XI11_5/XI0/XI0_52/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_15 XI11_5/XI0/XI0_52/d__15_ xsel_52_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_14 XI11_5/XI0/XI0_52/d__14_ xsel_52_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_13 XI11_5/XI0/XI0_52/d__13_ xsel_52_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_12 XI11_5/XI0/XI0_52/d__12_ xsel_52_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_11 XI11_5/XI0/XI0_52/d__11_ xsel_52_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_10 XI11_5/XI0/XI0_52/d__10_ xsel_52_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_9 XI11_5/XI0/XI0_52/d__9_ xsel_52_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_8 XI11_5/XI0/XI0_52/d__8_ xsel_52_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_7 XI11_5/XI0/XI0_52/d__7_ xsel_52_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_6 XI11_5/XI0/XI0_52/d__6_ xsel_52_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_5 XI11_5/XI0/XI0_52/d__5_ xsel_52_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_4 XI11_5/XI0/XI0_52/d__4_ xsel_52_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_3 XI11_5/XI0/XI0_52/d__3_ xsel_52_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_2 XI11_5/XI0/XI0_52/d__2_ xsel_52_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_1 XI11_5/XI0/XI0_52/d__1_ xsel_52_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_0 XI11_5/XI0/XI0_52/d__0_ xsel_52_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_15 XI11_5/net21_0_ xsel_51_ XI11_5/XI0/XI0_51/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_14 XI11_5/net21_1_ xsel_51_ XI11_5/XI0/XI0_51/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_13 XI11_5/net21_2_ xsel_51_ XI11_5/XI0/XI0_51/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_12 XI11_5/net21_3_ xsel_51_ XI11_5/XI0/XI0_51/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_11 XI11_5/net21_4_ xsel_51_ XI11_5/XI0/XI0_51/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_10 XI11_5/net21_5_ xsel_51_ XI11_5/XI0/XI0_51/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_9 XI11_5/net21_6_ xsel_51_ XI11_5/XI0/XI0_51/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_8 XI11_5/net21_7_ xsel_51_ XI11_5/XI0/XI0_51/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_7 XI11_5/net21_8_ xsel_51_ XI11_5/XI0/XI0_51/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_6 XI11_5/net21_9_ xsel_51_ XI11_5/XI0/XI0_51/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_5 XI11_5/net21_10_ xsel_51_ XI11_5/XI0/XI0_51/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_4 XI11_5/net21_11_ xsel_51_ XI11_5/XI0/XI0_51/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_3 XI11_5/net21_12_ xsel_51_ XI11_5/XI0/XI0_51/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_2 XI11_5/net21_13_ xsel_51_ XI11_5/XI0/XI0_51/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_1 XI11_5/net21_14_ xsel_51_ XI11_5/XI0/XI0_51/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_0 XI11_5/net21_15_ xsel_51_ XI11_5/XI0/XI0_51/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_15 XI11_5/XI0/XI0_51/d__15_ xsel_51_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_14 XI11_5/XI0/XI0_51/d__14_ xsel_51_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_13 XI11_5/XI0/XI0_51/d__13_ xsel_51_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_12 XI11_5/XI0/XI0_51/d__12_ xsel_51_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_11 XI11_5/XI0/XI0_51/d__11_ xsel_51_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_10 XI11_5/XI0/XI0_51/d__10_ xsel_51_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_9 XI11_5/XI0/XI0_51/d__9_ xsel_51_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_8 XI11_5/XI0/XI0_51/d__8_ xsel_51_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_7 XI11_5/XI0/XI0_51/d__7_ xsel_51_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_6 XI11_5/XI0/XI0_51/d__6_ xsel_51_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_5 XI11_5/XI0/XI0_51/d__5_ xsel_51_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_4 XI11_5/XI0/XI0_51/d__4_ xsel_51_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_3 XI11_5/XI0/XI0_51/d__3_ xsel_51_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_2 XI11_5/XI0/XI0_51/d__2_ xsel_51_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_1 XI11_5/XI0/XI0_51/d__1_ xsel_51_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_0 XI11_5/XI0/XI0_51/d__0_ xsel_51_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_15 XI11_5/net21_0_ xsel_50_ XI11_5/XI0/XI0_50/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_14 XI11_5/net21_1_ xsel_50_ XI11_5/XI0/XI0_50/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_13 XI11_5/net21_2_ xsel_50_ XI11_5/XI0/XI0_50/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_12 XI11_5/net21_3_ xsel_50_ XI11_5/XI0/XI0_50/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_11 XI11_5/net21_4_ xsel_50_ XI11_5/XI0/XI0_50/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_10 XI11_5/net21_5_ xsel_50_ XI11_5/XI0/XI0_50/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_9 XI11_5/net21_6_ xsel_50_ XI11_5/XI0/XI0_50/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_8 XI11_5/net21_7_ xsel_50_ XI11_5/XI0/XI0_50/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_7 XI11_5/net21_8_ xsel_50_ XI11_5/XI0/XI0_50/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_6 XI11_5/net21_9_ xsel_50_ XI11_5/XI0/XI0_50/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_5 XI11_5/net21_10_ xsel_50_ XI11_5/XI0/XI0_50/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_4 XI11_5/net21_11_ xsel_50_ XI11_5/XI0/XI0_50/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_3 XI11_5/net21_12_ xsel_50_ XI11_5/XI0/XI0_50/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_2 XI11_5/net21_13_ xsel_50_ XI11_5/XI0/XI0_50/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_1 XI11_5/net21_14_ xsel_50_ XI11_5/XI0/XI0_50/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_0 XI11_5/net21_15_ xsel_50_ XI11_5/XI0/XI0_50/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_15 XI11_5/XI0/XI0_50/d__15_ xsel_50_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_14 XI11_5/XI0/XI0_50/d__14_ xsel_50_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_13 XI11_5/XI0/XI0_50/d__13_ xsel_50_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_12 XI11_5/XI0/XI0_50/d__12_ xsel_50_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_11 XI11_5/XI0/XI0_50/d__11_ xsel_50_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_10 XI11_5/XI0/XI0_50/d__10_ xsel_50_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_9 XI11_5/XI0/XI0_50/d__9_ xsel_50_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_8 XI11_5/XI0/XI0_50/d__8_ xsel_50_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_7 XI11_5/XI0/XI0_50/d__7_ xsel_50_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_6 XI11_5/XI0/XI0_50/d__6_ xsel_50_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_5 XI11_5/XI0/XI0_50/d__5_ xsel_50_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_4 XI11_5/XI0/XI0_50/d__4_ xsel_50_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_3 XI11_5/XI0/XI0_50/d__3_ xsel_50_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_2 XI11_5/XI0/XI0_50/d__2_ xsel_50_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_1 XI11_5/XI0/XI0_50/d__1_ xsel_50_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_0 XI11_5/XI0/XI0_50/d__0_ xsel_50_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_15 XI11_5/net21_0_ xsel_49_ XI11_5/XI0/XI0_49/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_14 XI11_5/net21_1_ xsel_49_ XI11_5/XI0/XI0_49/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_13 XI11_5/net21_2_ xsel_49_ XI11_5/XI0/XI0_49/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_12 XI11_5/net21_3_ xsel_49_ XI11_5/XI0/XI0_49/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_11 XI11_5/net21_4_ xsel_49_ XI11_5/XI0/XI0_49/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_10 XI11_5/net21_5_ xsel_49_ XI11_5/XI0/XI0_49/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_9 XI11_5/net21_6_ xsel_49_ XI11_5/XI0/XI0_49/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_8 XI11_5/net21_7_ xsel_49_ XI11_5/XI0/XI0_49/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_7 XI11_5/net21_8_ xsel_49_ XI11_5/XI0/XI0_49/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_6 XI11_5/net21_9_ xsel_49_ XI11_5/XI0/XI0_49/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_5 XI11_5/net21_10_ xsel_49_ XI11_5/XI0/XI0_49/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_4 XI11_5/net21_11_ xsel_49_ XI11_5/XI0/XI0_49/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_3 XI11_5/net21_12_ xsel_49_ XI11_5/XI0/XI0_49/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_2 XI11_5/net21_13_ xsel_49_ XI11_5/XI0/XI0_49/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_1 XI11_5/net21_14_ xsel_49_ XI11_5/XI0/XI0_49/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_0 XI11_5/net21_15_ xsel_49_ XI11_5/XI0/XI0_49/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_15 XI11_5/XI0/XI0_49/d__15_ xsel_49_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_14 XI11_5/XI0/XI0_49/d__14_ xsel_49_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_13 XI11_5/XI0/XI0_49/d__13_ xsel_49_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_12 XI11_5/XI0/XI0_49/d__12_ xsel_49_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_11 XI11_5/XI0/XI0_49/d__11_ xsel_49_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_10 XI11_5/XI0/XI0_49/d__10_ xsel_49_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_9 XI11_5/XI0/XI0_49/d__9_ xsel_49_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_8 XI11_5/XI0/XI0_49/d__8_ xsel_49_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_7 XI11_5/XI0/XI0_49/d__7_ xsel_49_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_6 XI11_5/XI0/XI0_49/d__6_ xsel_49_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_5 XI11_5/XI0/XI0_49/d__5_ xsel_49_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_4 XI11_5/XI0/XI0_49/d__4_ xsel_49_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_3 XI11_5/XI0/XI0_49/d__3_ xsel_49_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_2 XI11_5/XI0/XI0_49/d__2_ xsel_49_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_1 XI11_5/XI0/XI0_49/d__1_ xsel_49_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_0 XI11_5/XI0/XI0_49/d__0_ xsel_49_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_15 XI11_5/net21_0_ xsel_48_ XI11_5/XI0/XI0_48/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_14 XI11_5/net21_1_ xsel_48_ XI11_5/XI0/XI0_48/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_13 XI11_5/net21_2_ xsel_48_ XI11_5/XI0/XI0_48/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_12 XI11_5/net21_3_ xsel_48_ XI11_5/XI0/XI0_48/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_11 XI11_5/net21_4_ xsel_48_ XI11_5/XI0/XI0_48/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_10 XI11_5/net21_5_ xsel_48_ XI11_5/XI0/XI0_48/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_9 XI11_5/net21_6_ xsel_48_ XI11_5/XI0/XI0_48/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_8 XI11_5/net21_7_ xsel_48_ XI11_5/XI0/XI0_48/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_7 XI11_5/net21_8_ xsel_48_ XI11_5/XI0/XI0_48/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_6 XI11_5/net21_9_ xsel_48_ XI11_5/XI0/XI0_48/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_5 XI11_5/net21_10_ xsel_48_ XI11_5/XI0/XI0_48/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_4 XI11_5/net21_11_ xsel_48_ XI11_5/XI0/XI0_48/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_3 XI11_5/net21_12_ xsel_48_ XI11_5/XI0/XI0_48/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_2 XI11_5/net21_13_ xsel_48_ XI11_5/XI0/XI0_48/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_1 XI11_5/net21_14_ xsel_48_ XI11_5/XI0/XI0_48/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_0 XI11_5/net21_15_ xsel_48_ XI11_5/XI0/XI0_48/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_15 XI11_5/XI0/XI0_48/d__15_ xsel_48_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_14 XI11_5/XI0/XI0_48/d__14_ xsel_48_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_13 XI11_5/XI0/XI0_48/d__13_ xsel_48_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_12 XI11_5/XI0/XI0_48/d__12_ xsel_48_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_11 XI11_5/XI0/XI0_48/d__11_ xsel_48_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_10 XI11_5/XI0/XI0_48/d__10_ xsel_48_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_9 XI11_5/XI0/XI0_48/d__9_ xsel_48_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_8 XI11_5/XI0/XI0_48/d__8_ xsel_48_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_7 XI11_5/XI0/XI0_48/d__7_ xsel_48_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_6 XI11_5/XI0/XI0_48/d__6_ xsel_48_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_5 XI11_5/XI0/XI0_48/d__5_ xsel_48_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_4 XI11_5/XI0/XI0_48/d__4_ xsel_48_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_3 XI11_5/XI0/XI0_48/d__3_ xsel_48_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_2 XI11_5/XI0/XI0_48/d__2_ xsel_48_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_1 XI11_5/XI0/XI0_48/d__1_ xsel_48_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_0 XI11_5/XI0/XI0_48/d__0_ xsel_48_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_15 XI11_5/net21_0_ xsel_47_ XI11_5/XI0/XI0_47/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_14 XI11_5/net21_1_ xsel_47_ XI11_5/XI0/XI0_47/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_13 XI11_5/net21_2_ xsel_47_ XI11_5/XI0/XI0_47/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_12 XI11_5/net21_3_ xsel_47_ XI11_5/XI0/XI0_47/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_11 XI11_5/net21_4_ xsel_47_ XI11_5/XI0/XI0_47/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_10 XI11_5/net21_5_ xsel_47_ XI11_5/XI0/XI0_47/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_9 XI11_5/net21_6_ xsel_47_ XI11_5/XI0/XI0_47/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_8 XI11_5/net21_7_ xsel_47_ XI11_5/XI0/XI0_47/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_7 XI11_5/net21_8_ xsel_47_ XI11_5/XI0/XI0_47/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_6 XI11_5/net21_9_ xsel_47_ XI11_5/XI0/XI0_47/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_5 XI11_5/net21_10_ xsel_47_ XI11_5/XI0/XI0_47/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_4 XI11_5/net21_11_ xsel_47_ XI11_5/XI0/XI0_47/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_3 XI11_5/net21_12_ xsel_47_ XI11_5/XI0/XI0_47/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_2 XI11_5/net21_13_ xsel_47_ XI11_5/XI0/XI0_47/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_1 XI11_5/net21_14_ xsel_47_ XI11_5/XI0/XI0_47/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_0 XI11_5/net21_15_ xsel_47_ XI11_5/XI0/XI0_47/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_15 XI11_5/XI0/XI0_47/d__15_ xsel_47_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_14 XI11_5/XI0/XI0_47/d__14_ xsel_47_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_13 XI11_5/XI0/XI0_47/d__13_ xsel_47_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_12 XI11_5/XI0/XI0_47/d__12_ xsel_47_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_11 XI11_5/XI0/XI0_47/d__11_ xsel_47_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_10 XI11_5/XI0/XI0_47/d__10_ xsel_47_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_9 XI11_5/XI0/XI0_47/d__9_ xsel_47_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_8 XI11_5/XI0/XI0_47/d__8_ xsel_47_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_7 XI11_5/XI0/XI0_47/d__7_ xsel_47_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_6 XI11_5/XI0/XI0_47/d__6_ xsel_47_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_5 XI11_5/XI0/XI0_47/d__5_ xsel_47_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_4 XI11_5/XI0/XI0_47/d__4_ xsel_47_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_3 XI11_5/XI0/XI0_47/d__3_ xsel_47_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_2 XI11_5/XI0/XI0_47/d__2_ xsel_47_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_1 XI11_5/XI0/XI0_47/d__1_ xsel_47_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_0 XI11_5/XI0/XI0_47/d__0_ xsel_47_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_15 XI11_5/net21_0_ xsel_46_ XI11_5/XI0/XI0_46/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_14 XI11_5/net21_1_ xsel_46_ XI11_5/XI0/XI0_46/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_13 XI11_5/net21_2_ xsel_46_ XI11_5/XI0/XI0_46/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_12 XI11_5/net21_3_ xsel_46_ XI11_5/XI0/XI0_46/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_11 XI11_5/net21_4_ xsel_46_ XI11_5/XI0/XI0_46/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_10 XI11_5/net21_5_ xsel_46_ XI11_5/XI0/XI0_46/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_9 XI11_5/net21_6_ xsel_46_ XI11_5/XI0/XI0_46/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_8 XI11_5/net21_7_ xsel_46_ XI11_5/XI0/XI0_46/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_7 XI11_5/net21_8_ xsel_46_ XI11_5/XI0/XI0_46/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_6 XI11_5/net21_9_ xsel_46_ XI11_5/XI0/XI0_46/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_5 XI11_5/net21_10_ xsel_46_ XI11_5/XI0/XI0_46/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_4 XI11_5/net21_11_ xsel_46_ XI11_5/XI0/XI0_46/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_3 XI11_5/net21_12_ xsel_46_ XI11_5/XI0/XI0_46/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_2 XI11_5/net21_13_ xsel_46_ XI11_5/XI0/XI0_46/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_1 XI11_5/net21_14_ xsel_46_ XI11_5/XI0/XI0_46/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_0 XI11_5/net21_15_ xsel_46_ XI11_5/XI0/XI0_46/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_15 XI11_5/XI0/XI0_46/d__15_ xsel_46_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_14 XI11_5/XI0/XI0_46/d__14_ xsel_46_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_13 XI11_5/XI0/XI0_46/d__13_ xsel_46_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_12 XI11_5/XI0/XI0_46/d__12_ xsel_46_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_11 XI11_5/XI0/XI0_46/d__11_ xsel_46_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_10 XI11_5/XI0/XI0_46/d__10_ xsel_46_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_9 XI11_5/XI0/XI0_46/d__9_ xsel_46_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_8 XI11_5/XI0/XI0_46/d__8_ xsel_46_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_7 XI11_5/XI0/XI0_46/d__7_ xsel_46_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_6 XI11_5/XI0/XI0_46/d__6_ xsel_46_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_5 XI11_5/XI0/XI0_46/d__5_ xsel_46_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_4 XI11_5/XI0/XI0_46/d__4_ xsel_46_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_3 XI11_5/XI0/XI0_46/d__3_ xsel_46_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_2 XI11_5/XI0/XI0_46/d__2_ xsel_46_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_1 XI11_5/XI0/XI0_46/d__1_ xsel_46_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_0 XI11_5/XI0/XI0_46/d__0_ xsel_46_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_15 XI11_5/net21_0_ xsel_45_ XI11_5/XI0/XI0_45/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_14 XI11_5/net21_1_ xsel_45_ XI11_5/XI0/XI0_45/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_13 XI11_5/net21_2_ xsel_45_ XI11_5/XI0/XI0_45/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_12 XI11_5/net21_3_ xsel_45_ XI11_5/XI0/XI0_45/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_11 XI11_5/net21_4_ xsel_45_ XI11_5/XI0/XI0_45/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_10 XI11_5/net21_5_ xsel_45_ XI11_5/XI0/XI0_45/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_9 XI11_5/net21_6_ xsel_45_ XI11_5/XI0/XI0_45/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_8 XI11_5/net21_7_ xsel_45_ XI11_5/XI0/XI0_45/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_7 XI11_5/net21_8_ xsel_45_ XI11_5/XI0/XI0_45/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_6 XI11_5/net21_9_ xsel_45_ XI11_5/XI0/XI0_45/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_5 XI11_5/net21_10_ xsel_45_ XI11_5/XI0/XI0_45/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_4 XI11_5/net21_11_ xsel_45_ XI11_5/XI0/XI0_45/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_3 XI11_5/net21_12_ xsel_45_ XI11_5/XI0/XI0_45/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_2 XI11_5/net21_13_ xsel_45_ XI11_5/XI0/XI0_45/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_1 XI11_5/net21_14_ xsel_45_ XI11_5/XI0/XI0_45/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_0 XI11_5/net21_15_ xsel_45_ XI11_5/XI0/XI0_45/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_15 XI11_5/XI0/XI0_45/d__15_ xsel_45_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_14 XI11_5/XI0/XI0_45/d__14_ xsel_45_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_13 XI11_5/XI0/XI0_45/d__13_ xsel_45_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_12 XI11_5/XI0/XI0_45/d__12_ xsel_45_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_11 XI11_5/XI0/XI0_45/d__11_ xsel_45_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_10 XI11_5/XI0/XI0_45/d__10_ xsel_45_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_9 XI11_5/XI0/XI0_45/d__9_ xsel_45_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_8 XI11_5/XI0/XI0_45/d__8_ xsel_45_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_7 XI11_5/XI0/XI0_45/d__7_ xsel_45_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_6 XI11_5/XI0/XI0_45/d__6_ xsel_45_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_5 XI11_5/XI0/XI0_45/d__5_ xsel_45_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_4 XI11_5/XI0/XI0_45/d__4_ xsel_45_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_3 XI11_5/XI0/XI0_45/d__3_ xsel_45_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_2 XI11_5/XI0/XI0_45/d__2_ xsel_45_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_1 XI11_5/XI0/XI0_45/d__1_ xsel_45_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_0 XI11_5/XI0/XI0_45/d__0_ xsel_45_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_15 XI11_5/net21_0_ xsel_44_ XI11_5/XI0/XI0_44/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_14 XI11_5/net21_1_ xsel_44_ XI11_5/XI0/XI0_44/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_13 XI11_5/net21_2_ xsel_44_ XI11_5/XI0/XI0_44/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_12 XI11_5/net21_3_ xsel_44_ XI11_5/XI0/XI0_44/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_11 XI11_5/net21_4_ xsel_44_ XI11_5/XI0/XI0_44/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_10 XI11_5/net21_5_ xsel_44_ XI11_5/XI0/XI0_44/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_9 XI11_5/net21_6_ xsel_44_ XI11_5/XI0/XI0_44/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_8 XI11_5/net21_7_ xsel_44_ XI11_5/XI0/XI0_44/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_7 XI11_5/net21_8_ xsel_44_ XI11_5/XI0/XI0_44/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_6 XI11_5/net21_9_ xsel_44_ XI11_5/XI0/XI0_44/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_5 XI11_5/net21_10_ xsel_44_ XI11_5/XI0/XI0_44/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_4 XI11_5/net21_11_ xsel_44_ XI11_5/XI0/XI0_44/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_3 XI11_5/net21_12_ xsel_44_ XI11_5/XI0/XI0_44/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_2 XI11_5/net21_13_ xsel_44_ XI11_5/XI0/XI0_44/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_1 XI11_5/net21_14_ xsel_44_ XI11_5/XI0/XI0_44/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_0 XI11_5/net21_15_ xsel_44_ XI11_5/XI0/XI0_44/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_15 XI11_5/XI0/XI0_44/d__15_ xsel_44_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_14 XI11_5/XI0/XI0_44/d__14_ xsel_44_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_13 XI11_5/XI0/XI0_44/d__13_ xsel_44_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_12 XI11_5/XI0/XI0_44/d__12_ xsel_44_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_11 XI11_5/XI0/XI0_44/d__11_ xsel_44_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_10 XI11_5/XI0/XI0_44/d__10_ xsel_44_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_9 XI11_5/XI0/XI0_44/d__9_ xsel_44_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_8 XI11_5/XI0/XI0_44/d__8_ xsel_44_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_7 XI11_5/XI0/XI0_44/d__7_ xsel_44_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_6 XI11_5/XI0/XI0_44/d__6_ xsel_44_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_5 XI11_5/XI0/XI0_44/d__5_ xsel_44_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_4 XI11_5/XI0/XI0_44/d__4_ xsel_44_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_3 XI11_5/XI0/XI0_44/d__3_ xsel_44_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_2 XI11_5/XI0/XI0_44/d__2_ xsel_44_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_1 XI11_5/XI0/XI0_44/d__1_ xsel_44_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_0 XI11_5/XI0/XI0_44/d__0_ xsel_44_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_15 XI11_5/net21_0_ xsel_43_ XI11_5/XI0/XI0_43/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_14 XI11_5/net21_1_ xsel_43_ XI11_5/XI0/XI0_43/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_13 XI11_5/net21_2_ xsel_43_ XI11_5/XI0/XI0_43/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_12 XI11_5/net21_3_ xsel_43_ XI11_5/XI0/XI0_43/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_11 XI11_5/net21_4_ xsel_43_ XI11_5/XI0/XI0_43/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_10 XI11_5/net21_5_ xsel_43_ XI11_5/XI0/XI0_43/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_9 XI11_5/net21_6_ xsel_43_ XI11_5/XI0/XI0_43/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_8 XI11_5/net21_7_ xsel_43_ XI11_5/XI0/XI0_43/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_7 XI11_5/net21_8_ xsel_43_ XI11_5/XI0/XI0_43/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_6 XI11_5/net21_9_ xsel_43_ XI11_5/XI0/XI0_43/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_5 XI11_5/net21_10_ xsel_43_ XI11_5/XI0/XI0_43/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_4 XI11_5/net21_11_ xsel_43_ XI11_5/XI0/XI0_43/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_3 XI11_5/net21_12_ xsel_43_ XI11_5/XI0/XI0_43/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_2 XI11_5/net21_13_ xsel_43_ XI11_5/XI0/XI0_43/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_1 XI11_5/net21_14_ xsel_43_ XI11_5/XI0/XI0_43/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_0 XI11_5/net21_15_ xsel_43_ XI11_5/XI0/XI0_43/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_15 XI11_5/XI0/XI0_43/d__15_ xsel_43_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_14 XI11_5/XI0/XI0_43/d__14_ xsel_43_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_13 XI11_5/XI0/XI0_43/d__13_ xsel_43_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_12 XI11_5/XI0/XI0_43/d__12_ xsel_43_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_11 XI11_5/XI0/XI0_43/d__11_ xsel_43_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_10 XI11_5/XI0/XI0_43/d__10_ xsel_43_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_9 XI11_5/XI0/XI0_43/d__9_ xsel_43_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_8 XI11_5/XI0/XI0_43/d__8_ xsel_43_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_7 XI11_5/XI0/XI0_43/d__7_ xsel_43_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_6 XI11_5/XI0/XI0_43/d__6_ xsel_43_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_5 XI11_5/XI0/XI0_43/d__5_ xsel_43_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_4 XI11_5/XI0/XI0_43/d__4_ xsel_43_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_3 XI11_5/XI0/XI0_43/d__3_ xsel_43_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_2 XI11_5/XI0/XI0_43/d__2_ xsel_43_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_1 XI11_5/XI0/XI0_43/d__1_ xsel_43_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_0 XI11_5/XI0/XI0_43/d__0_ xsel_43_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_15 XI11_5/net21_0_ xsel_42_ XI11_5/XI0/XI0_42/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_14 XI11_5/net21_1_ xsel_42_ XI11_5/XI0/XI0_42/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_13 XI11_5/net21_2_ xsel_42_ XI11_5/XI0/XI0_42/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_12 XI11_5/net21_3_ xsel_42_ XI11_5/XI0/XI0_42/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_11 XI11_5/net21_4_ xsel_42_ XI11_5/XI0/XI0_42/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_10 XI11_5/net21_5_ xsel_42_ XI11_5/XI0/XI0_42/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_9 XI11_5/net21_6_ xsel_42_ XI11_5/XI0/XI0_42/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_8 XI11_5/net21_7_ xsel_42_ XI11_5/XI0/XI0_42/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_7 XI11_5/net21_8_ xsel_42_ XI11_5/XI0/XI0_42/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_6 XI11_5/net21_9_ xsel_42_ XI11_5/XI0/XI0_42/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_5 XI11_5/net21_10_ xsel_42_ XI11_5/XI0/XI0_42/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_4 XI11_5/net21_11_ xsel_42_ XI11_5/XI0/XI0_42/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_3 XI11_5/net21_12_ xsel_42_ XI11_5/XI0/XI0_42/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_2 XI11_5/net21_13_ xsel_42_ XI11_5/XI0/XI0_42/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_1 XI11_5/net21_14_ xsel_42_ XI11_5/XI0/XI0_42/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_0 XI11_5/net21_15_ xsel_42_ XI11_5/XI0/XI0_42/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_15 XI11_5/XI0/XI0_42/d__15_ xsel_42_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_14 XI11_5/XI0/XI0_42/d__14_ xsel_42_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_13 XI11_5/XI0/XI0_42/d__13_ xsel_42_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_12 XI11_5/XI0/XI0_42/d__12_ xsel_42_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_11 XI11_5/XI0/XI0_42/d__11_ xsel_42_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_10 XI11_5/XI0/XI0_42/d__10_ xsel_42_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_9 XI11_5/XI0/XI0_42/d__9_ xsel_42_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_8 XI11_5/XI0/XI0_42/d__8_ xsel_42_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_7 XI11_5/XI0/XI0_42/d__7_ xsel_42_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_6 XI11_5/XI0/XI0_42/d__6_ xsel_42_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_5 XI11_5/XI0/XI0_42/d__5_ xsel_42_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_4 XI11_5/XI0/XI0_42/d__4_ xsel_42_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_3 XI11_5/XI0/XI0_42/d__3_ xsel_42_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_2 XI11_5/XI0/XI0_42/d__2_ xsel_42_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_1 XI11_5/XI0/XI0_42/d__1_ xsel_42_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_0 XI11_5/XI0/XI0_42/d__0_ xsel_42_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_15 XI11_5/net21_0_ xsel_41_ XI11_5/XI0/XI0_41/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_14 XI11_5/net21_1_ xsel_41_ XI11_5/XI0/XI0_41/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_13 XI11_5/net21_2_ xsel_41_ XI11_5/XI0/XI0_41/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_12 XI11_5/net21_3_ xsel_41_ XI11_5/XI0/XI0_41/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_11 XI11_5/net21_4_ xsel_41_ XI11_5/XI0/XI0_41/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_10 XI11_5/net21_5_ xsel_41_ XI11_5/XI0/XI0_41/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_9 XI11_5/net21_6_ xsel_41_ XI11_5/XI0/XI0_41/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_8 XI11_5/net21_7_ xsel_41_ XI11_5/XI0/XI0_41/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_7 XI11_5/net21_8_ xsel_41_ XI11_5/XI0/XI0_41/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_6 XI11_5/net21_9_ xsel_41_ XI11_5/XI0/XI0_41/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_5 XI11_5/net21_10_ xsel_41_ XI11_5/XI0/XI0_41/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_4 XI11_5/net21_11_ xsel_41_ XI11_5/XI0/XI0_41/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_3 XI11_5/net21_12_ xsel_41_ XI11_5/XI0/XI0_41/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_2 XI11_5/net21_13_ xsel_41_ XI11_5/XI0/XI0_41/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_1 XI11_5/net21_14_ xsel_41_ XI11_5/XI0/XI0_41/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_0 XI11_5/net21_15_ xsel_41_ XI11_5/XI0/XI0_41/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_15 XI11_5/XI0/XI0_41/d__15_ xsel_41_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_14 XI11_5/XI0/XI0_41/d__14_ xsel_41_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_13 XI11_5/XI0/XI0_41/d__13_ xsel_41_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_12 XI11_5/XI0/XI0_41/d__12_ xsel_41_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_11 XI11_5/XI0/XI0_41/d__11_ xsel_41_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_10 XI11_5/XI0/XI0_41/d__10_ xsel_41_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_9 XI11_5/XI0/XI0_41/d__9_ xsel_41_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_8 XI11_5/XI0/XI0_41/d__8_ xsel_41_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_7 XI11_5/XI0/XI0_41/d__7_ xsel_41_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_6 XI11_5/XI0/XI0_41/d__6_ xsel_41_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_5 XI11_5/XI0/XI0_41/d__5_ xsel_41_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_4 XI11_5/XI0/XI0_41/d__4_ xsel_41_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_3 XI11_5/XI0/XI0_41/d__3_ xsel_41_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_2 XI11_5/XI0/XI0_41/d__2_ xsel_41_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_1 XI11_5/XI0/XI0_41/d__1_ xsel_41_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_0 XI11_5/XI0/XI0_41/d__0_ xsel_41_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_15 XI11_5/net21_0_ xsel_40_ XI11_5/XI0/XI0_40/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_14 XI11_5/net21_1_ xsel_40_ XI11_5/XI0/XI0_40/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_13 XI11_5/net21_2_ xsel_40_ XI11_5/XI0/XI0_40/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_12 XI11_5/net21_3_ xsel_40_ XI11_5/XI0/XI0_40/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_11 XI11_5/net21_4_ xsel_40_ XI11_5/XI0/XI0_40/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_10 XI11_5/net21_5_ xsel_40_ XI11_5/XI0/XI0_40/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_9 XI11_5/net21_6_ xsel_40_ XI11_5/XI0/XI0_40/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_8 XI11_5/net21_7_ xsel_40_ XI11_5/XI0/XI0_40/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_7 XI11_5/net21_8_ xsel_40_ XI11_5/XI0/XI0_40/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_6 XI11_5/net21_9_ xsel_40_ XI11_5/XI0/XI0_40/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_5 XI11_5/net21_10_ xsel_40_ XI11_5/XI0/XI0_40/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_4 XI11_5/net21_11_ xsel_40_ XI11_5/XI0/XI0_40/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_3 XI11_5/net21_12_ xsel_40_ XI11_5/XI0/XI0_40/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_2 XI11_5/net21_13_ xsel_40_ XI11_5/XI0/XI0_40/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_1 XI11_5/net21_14_ xsel_40_ XI11_5/XI0/XI0_40/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_0 XI11_5/net21_15_ xsel_40_ XI11_5/XI0/XI0_40/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_15 XI11_5/XI0/XI0_40/d__15_ xsel_40_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_14 XI11_5/XI0/XI0_40/d__14_ xsel_40_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_13 XI11_5/XI0/XI0_40/d__13_ xsel_40_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_12 XI11_5/XI0/XI0_40/d__12_ xsel_40_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_11 XI11_5/XI0/XI0_40/d__11_ xsel_40_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_10 XI11_5/XI0/XI0_40/d__10_ xsel_40_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_9 XI11_5/XI0/XI0_40/d__9_ xsel_40_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_8 XI11_5/XI0/XI0_40/d__8_ xsel_40_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_7 XI11_5/XI0/XI0_40/d__7_ xsel_40_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_6 XI11_5/XI0/XI0_40/d__6_ xsel_40_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_5 XI11_5/XI0/XI0_40/d__5_ xsel_40_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_4 XI11_5/XI0/XI0_40/d__4_ xsel_40_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_3 XI11_5/XI0/XI0_40/d__3_ xsel_40_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_2 XI11_5/XI0/XI0_40/d__2_ xsel_40_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_1 XI11_5/XI0/XI0_40/d__1_ xsel_40_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_0 XI11_5/XI0/XI0_40/d__0_ xsel_40_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_15 XI11_5/net21_0_ xsel_39_ XI11_5/XI0/XI0_39/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_14 XI11_5/net21_1_ xsel_39_ XI11_5/XI0/XI0_39/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_13 XI11_5/net21_2_ xsel_39_ XI11_5/XI0/XI0_39/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_12 XI11_5/net21_3_ xsel_39_ XI11_5/XI0/XI0_39/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_11 XI11_5/net21_4_ xsel_39_ XI11_5/XI0/XI0_39/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_10 XI11_5/net21_5_ xsel_39_ XI11_5/XI0/XI0_39/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_9 XI11_5/net21_6_ xsel_39_ XI11_5/XI0/XI0_39/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_8 XI11_5/net21_7_ xsel_39_ XI11_5/XI0/XI0_39/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_7 XI11_5/net21_8_ xsel_39_ XI11_5/XI0/XI0_39/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_6 XI11_5/net21_9_ xsel_39_ XI11_5/XI0/XI0_39/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_5 XI11_5/net21_10_ xsel_39_ XI11_5/XI0/XI0_39/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_4 XI11_5/net21_11_ xsel_39_ XI11_5/XI0/XI0_39/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_3 XI11_5/net21_12_ xsel_39_ XI11_5/XI0/XI0_39/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_2 XI11_5/net21_13_ xsel_39_ XI11_5/XI0/XI0_39/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_1 XI11_5/net21_14_ xsel_39_ XI11_5/XI0/XI0_39/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_0 XI11_5/net21_15_ xsel_39_ XI11_5/XI0/XI0_39/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_15 XI11_5/XI0/XI0_39/d__15_ xsel_39_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_14 XI11_5/XI0/XI0_39/d__14_ xsel_39_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_13 XI11_5/XI0/XI0_39/d__13_ xsel_39_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_12 XI11_5/XI0/XI0_39/d__12_ xsel_39_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_11 XI11_5/XI0/XI0_39/d__11_ xsel_39_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_10 XI11_5/XI0/XI0_39/d__10_ xsel_39_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_9 XI11_5/XI0/XI0_39/d__9_ xsel_39_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_8 XI11_5/XI0/XI0_39/d__8_ xsel_39_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_7 XI11_5/XI0/XI0_39/d__7_ xsel_39_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_6 XI11_5/XI0/XI0_39/d__6_ xsel_39_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_5 XI11_5/XI0/XI0_39/d__5_ xsel_39_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_4 XI11_5/XI0/XI0_39/d__4_ xsel_39_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_3 XI11_5/XI0/XI0_39/d__3_ xsel_39_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_2 XI11_5/XI0/XI0_39/d__2_ xsel_39_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_1 XI11_5/XI0/XI0_39/d__1_ xsel_39_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_0 XI11_5/XI0/XI0_39/d__0_ xsel_39_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_15 XI11_5/net21_0_ xsel_38_ XI11_5/XI0/XI0_38/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_14 XI11_5/net21_1_ xsel_38_ XI11_5/XI0/XI0_38/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_13 XI11_5/net21_2_ xsel_38_ XI11_5/XI0/XI0_38/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_12 XI11_5/net21_3_ xsel_38_ XI11_5/XI0/XI0_38/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_11 XI11_5/net21_4_ xsel_38_ XI11_5/XI0/XI0_38/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_10 XI11_5/net21_5_ xsel_38_ XI11_5/XI0/XI0_38/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_9 XI11_5/net21_6_ xsel_38_ XI11_5/XI0/XI0_38/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_8 XI11_5/net21_7_ xsel_38_ XI11_5/XI0/XI0_38/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_7 XI11_5/net21_8_ xsel_38_ XI11_5/XI0/XI0_38/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_6 XI11_5/net21_9_ xsel_38_ XI11_5/XI0/XI0_38/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_5 XI11_5/net21_10_ xsel_38_ XI11_5/XI0/XI0_38/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_4 XI11_5/net21_11_ xsel_38_ XI11_5/XI0/XI0_38/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_3 XI11_5/net21_12_ xsel_38_ XI11_5/XI0/XI0_38/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_2 XI11_5/net21_13_ xsel_38_ XI11_5/XI0/XI0_38/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_1 XI11_5/net21_14_ xsel_38_ XI11_5/XI0/XI0_38/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_0 XI11_5/net21_15_ xsel_38_ XI11_5/XI0/XI0_38/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_15 XI11_5/XI0/XI0_38/d__15_ xsel_38_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_14 XI11_5/XI0/XI0_38/d__14_ xsel_38_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_13 XI11_5/XI0/XI0_38/d__13_ xsel_38_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_12 XI11_5/XI0/XI0_38/d__12_ xsel_38_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_11 XI11_5/XI0/XI0_38/d__11_ xsel_38_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_10 XI11_5/XI0/XI0_38/d__10_ xsel_38_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_9 XI11_5/XI0/XI0_38/d__9_ xsel_38_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_8 XI11_5/XI0/XI0_38/d__8_ xsel_38_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_7 XI11_5/XI0/XI0_38/d__7_ xsel_38_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_6 XI11_5/XI0/XI0_38/d__6_ xsel_38_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_5 XI11_5/XI0/XI0_38/d__5_ xsel_38_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_4 XI11_5/XI0/XI0_38/d__4_ xsel_38_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_3 XI11_5/XI0/XI0_38/d__3_ xsel_38_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_2 XI11_5/XI0/XI0_38/d__2_ xsel_38_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_1 XI11_5/XI0/XI0_38/d__1_ xsel_38_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_0 XI11_5/XI0/XI0_38/d__0_ xsel_38_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_15 XI11_5/net21_0_ xsel_37_ XI11_5/XI0/XI0_37/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_14 XI11_5/net21_1_ xsel_37_ XI11_5/XI0/XI0_37/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_13 XI11_5/net21_2_ xsel_37_ XI11_5/XI0/XI0_37/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_12 XI11_5/net21_3_ xsel_37_ XI11_5/XI0/XI0_37/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_11 XI11_5/net21_4_ xsel_37_ XI11_5/XI0/XI0_37/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_10 XI11_5/net21_5_ xsel_37_ XI11_5/XI0/XI0_37/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_9 XI11_5/net21_6_ xsel_37_ XI11_5/XI0/XI0_37/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_8 XI11_5/net21_7_ xsel_37_ XI11_5/XI0/XI0_37/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_7 XI11_5/net21_8_ xsel_37_ XI11_5/XI0/XI0_37/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_6 XI11_5/net21_9_ xsel_37_ XI11_5/XI0/XI0_37/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_5 XI11_5/net21_10_ xsel_37_ XI11_5/XI0/XI0_37/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_4 XI11_5/net21_11_ xsel_37_ XI11_5/XI0/XI0_37/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_3 XI11_5/net21_12_ xsel_37_ XI11_5/XI0/XI0_37/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_2 XI11_5/net21_13_ xsel_37_ XI11_5/XI0/XI0_37/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_1 XI11_5/net21_14_ xsel_37_ XI11_5/XI0/XI0_37/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_0 XI11_5/net21_15_ xsel_37_ XI11_5/XI0/XI0_37/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_15 XI11_5/XI0/XI0_37/d__15_ xsel_37_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_14 XI11_5/XI0/XI0_37/d__14_ xsel_37_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_13 XI11_5/XI0/XI0_37/d__13_ xsel_37_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_12 XI11_5/XI0/XI0_37/d__12_ xsel_37_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_11 XI11_5/XI0/XI0_37/d__11_ xsel_37_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_10 XI11_5/XI0/XI0_37/d__10_ xsel_37_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_9 XI11_5/XI0/XI0_37/d__9_ xsel_37_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_8 XI11_5/XI0/XI0_37/d__8_ xsel_37_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_7 XI11_5/XI0/XI0_37/d__7_ xsel_37_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_6 XI11_5/XI0/XI0_37/d__6_ xsel_37_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_5 XI11_5/XI0/XI0_37/d__5_ xsel_37_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_4 XI11_5/XI0/XI0_37/d__4_ xsel_37_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_3 XI11_5/XI0/XI0_37/d__3_ xsel_37_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_2 XI11_5/XI0/XI0_37/d__2_ xsel_37_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_1 XI11_5/XI0/XI0_37/d__1_ xsel_37_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_0 XI11_5/XI0/XI0_37/d__0_ xsel_37_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_15 XI11_5/net21_0_ xsel_36_ XI11_5/XI0/XI0_36/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_14 XI11_5/net21_1_ xsel_36_ XI11_5/XI0/XI0_36/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_13 XI11_5/net21_2_ xsel_36_ XI11_5/XI0/XI0_36/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_12 XI11_5/net21_3_ xsel_36_ XI11_5/XI0/XI0_36/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_11 XI11_5/net21_4_ xsel_36_ XI11_5/XI0/XI0_36/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_10 XI11_5/net21_5_ xsel_36_ XI11_5/XI0/XI0_36/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_9 XI11_5/net21_6_ xsel_36_ XI11_5/XI0/XI0_36/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_8 XI11_5/net21_7_ xsel_36_ XI11_5/XI0/XI0_36/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_7 XI11_5/net21_8_ xsel_36_ XI11_5/XI0/XI0_36/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_6 XI11_5/net21_9_ xsel_36_ XI11_5/XI0/XI0_36/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_5 XI11_5/net21_10_ xsel_36_ XI11_5/XI0/XI0_36/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_4 XI11_5/net21_11_ xsel_36_ XI11_5/XI0/XI0_36/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_3 XI11_5/net21_12_ xsel_36_ XI11_5/XI0/XI0_36/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_2 XI11_5/net21_13_ xsel_36_ XI11_5/XI0/XI0_36/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_1 XI11_5/net21_14_ xsel_36_ XI11_5/XI0/XI0_36/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_0 XI11_5/net21_15_ xsel_36_ XI11_5/XI0/XI0_36/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_15 XI11_5/XI0/XI0_36/d__15_ xsel_36_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_14 XI11_5/XI0/XI0_36/d__14_ xsel_36_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_13 XI11_5/XI0/XI0_36/d__13_ xsel_36_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_12 XI11_5/XI0/XI0_36/d__12_ xsel_36_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_11 XI11_5/XI0/XI0_36/d__11_ xsel_36_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_10 XI11_5/XI0/XI0_36/d__10_ xsel_36_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_9 XI11_5/XI0/XI0_36/d__9_ xsel_36_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_8 XI11_5/XI0/XI0_36/d__8_ xsel_36_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_7 XI11_5/XI0/XI0_36/d__7_ xsel_36_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_6 XI11_5/XI0/XI0_36/d__6_ xsel_36_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_5 XI11_5/XI0/XI0_36/d__5_ xsel_36_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_4 XI11_5/XI0/XI0_36/d__4_ xsel_36_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_3 XI11_5/XI0/XI0_36/d__3_ xsel_36_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_2 XI11_5/XI0/XI0_36/d__2_ xsel_36_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_1 XI11_5/XI0/XI0_36/d__1_ xsel_36_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_0 XI11_5/XI0/XI0_36/d__0_ xsel_36_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_15 XI11_5/net21_0_ xsel_35_ XI11_5/XI0/XI0_35/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_14 XI11_5/net21_1_ xsel_35_ XI11_5/XI0/XI0_35/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_13 XI11_5/net21_2_ xsel_35_ XI11_5/XI0/XI0_35/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_12 XI11_5/net21_3_ xsel_35_ XI11_5/XI0/XI0_35/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_11 XI11_5/net21_4_ xsel_35_ XI11_5/XI0/XI0_35/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_10 XI11_5/net21_5_ xsel_35_ XI11_5/XI0/XI0_35/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_9 XI11_5/net21_6_ xsel_35_ XI11_5/XI0/XI0_35/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_8 XI11_5/net21_7_ xsel_35_ XI11_5/XI0/XI0_35/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_7 XI11_5/net21_8_ xsel_35_ XI11_5/XI0/XI0_35/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_6 XI11_5/net21_9_ xsel_35_ XI11_5/XI0/XI0_35/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_5 XI11_5/net21_10_ xsel_35_ XI11_5/XI0/XI0_35/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_4 XI11_5/net21_11_ xsel_35_ XI11_5/XI0/XI0_35/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_3 XI11_5/net21_12_ xsel_35_ XI11_5/XI0/XI0_35/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_2 XI11_5/net21_13_ xsel_35_ XI11_5/XI0/XI0_35/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_1 XI11_5/net21_14_ xsel_35_ XI11_5/XI0/XI0_35/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_0 XI11_5/net21_15_ xsel_35_ XI11_5/XI0/XI0_35/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_15 XI11_5/XI0/XI0_35/d__15_ xsel_35_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_14 XI11_5/XI0/XI0_35/d__14_ xsel_35_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_13 XI11_5/XI0/XI0_35/d__13_ xsel_35_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_12 XI11_5/XI0/XI0_35/d__12_ xsel_35_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_11 XI11_5/XI0/XI0_35/d__11_ xsel_35_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_10 XI11_5/XI0/XI0_35/d__10_ xsel_35_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_9 XI11_5/XI0/XI0_35/d__9_ xsel_35_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_8 XI11_5/XI0/XI0_35/d__8_ xsel_35_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_7 XI11_5/XI0/XI0_35/d__7_ xsel_35_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_6 XI11_5/XI0/XI0_35/d__6_ xsel_35_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_5 XI11_5/XI0/XI0_35/d__5_ xsel_35_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_4 XI11_5/XI0/XI0_35/d__4_ xsel_35_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_3 XI11_5/XI0/XI0_35/d__3_ xsel_35_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_2 XI11_5/XI0/XI0_35/d__2_ xsel_35_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_1 XI11_5/XI0/XI0_35/d__1_ xsel_35_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_0 XI11_5/XI0/XI0_35/d__0_ xsel_35_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_15 XI11_5/net21_0_ xsel_34_ XI11_5/XI0/XI0_34/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_14 XI11_5/net21_1_ xsel_34_ XI11_5/XI0/XI0_34/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_13 XI11_5/net21_2_ xsel_34_ XI11_5/XI0/XI0_34/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_12 XI11_5/net21_3_ xsel_34_ XI11_5/XI0/XI0_34/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_11 XI11_5/net21_4_ xsel_34_ XI11_5/XI0/XI0_34/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_10 XI11_5/net21_5_ xsel_34_ XI11_5/XI0/XI0_34/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_9 XI11_5/net21_6_ xsel_34_ XI11_5/XI0/XI0_34/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_8 XI11_5/net21_7_ xsel_34_ XI11_5/XI0/XI0_34/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_7 XI11_5/net21_8_ xsel_34_ XI11_5/XI0/XI0_34/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_6 XI11_5/net21_9_ xsel_34_ XI11_5/XI0/XI0_34/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_5 XI11_5/net21_10_ xsel_34_ XI11_5/XI0/XI0_34/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_4 XI11_5/net21_11_ xsel_34_ XI11_5/XI0/XI0_34/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_3 XI11_5/net21_12_ xsel_34_ XI11_5/XI0/XI0_34/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_2 XI11_5/net21_13_ xsel_34_ XI11_5/XI0/XI0_34/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_1 XI11_5/net21_14_ xsel_34_ XI11_5/XI0/XI0_34/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_0 XI11_5/net21_15_ xsel_34_ XI11_5/XI0/XI0_34/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_15 XI11_5/XI0/XI0_34/d__15_ xsel_34_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_14 XI11_5/XI0/XI0_34/d__14_ xsel_34_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_13 XI11_5/XI0/XI0_34/d__13_ xsel_34_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_12 XI11_5/XI0/XI0_34/d__12_ xsel_34_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_11 XI11_5/XI0/XI0_34/d__11_ xsel_34_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_10 XI11_5/XI0/XI0_34/d__10_ xsel_34_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_9 XI11_5/XI0/XI0_34/d__9_ xsel_34_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_8 XI11_5/XI0/XI0_34/d__8_ xsel_34_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_7 XI11_5/XI0/XI0_34/d__7_ xsel_34_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_6 XI11_5/XI0/XI0_34/d__6_ xsel_34_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_5 XI11_5/XI0/XI0_34/d__5_ xsel_34_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_4 XI11_5/XI0/XI0_34/d__4_ xsel_34_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_3 XI11_5/XI0/XI0_34/d__3_ xsel_34_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_2 XI11_5/XI0/XI0_34/d__2_ xsel_34_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_1 XI11_5/XI0/XI0_34/d__1_ xsel_34_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_0 XI11_5/XI0/XI0_34/d__0_ xsel_34_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_15 XI11_5/net21_0_ xsel_33_ XI11_5/XI0/XI0_33/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_14 XI11_5/net21_1_ xsel_33_ XI11_5/XI0/XI0_33/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_13 XI11_5/net21_2_ xsel_33_ XI11_5/XI0/XI0_33/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_12 XI11_5/net21_3_ xsel_33_ XI11_5/XI0/XI0_33/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_11 XI11_5/net21_4_ xsel_33_ XI11_5/XI0/XI0_33/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_10 XI11_5/net21_5_ xsel_33_ XI11_5/XI0/XI0_33/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_9 XI11_5/net21_6_ xsel_33_ XI11_5/XI0/XI0_33/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_8 XI11_5/net21_7_ xsel_33_ XI11_5/XI0/XI0_33/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_7 XI11_5/net21_8_ xsel_33_ XI11_5/XI0/XI0_33/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_6 XI11_5/net21_9_ xsel_33_ XI11_5/XI0/XI0_33/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_5 XI11_5/net21_10_ xsel_33_ XI11_5/XI0/XI0_33/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_4 XI11_5/net21_11_ xsel_33_ XI11_5/XI0/XI0_33/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_3 XI11_5/net21_12_ xsel_33_ XI11_5/XI0/XI0_33/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_2 XI11_5/net21_13_ xsel_33_ XI11_5/XI0/XI0_33/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_1 XI11_5/net21_14_ xsel_33_ XI11_5/XI0/XI0_33/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_0 XI11_5/net21_15_ xsel_33_ XI11_5/XI0/XI0_33/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_15 XI11_5/XI0/XI0_33/d__15_ xsel_33_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_14 XI11_5/XI0/XI0_33/d__14_ xsel_33_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_13 XI11_5/XI0/XI0_33/d__13_ xsel_33_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_12 XI11_5/XI0/XI0_33/d__12_ xsel_33_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_11 XI11_5/XI0/XI0_33/d__11_ xsel_33_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_10 XI11_5/XI0/XI0_33/d__10_ xsel_33_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_9 XI11_5/XI0/XI0_33/d__9_ xsel_33_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_8 XI11_5/XI0/XI0_33/d__8_ xsel_33_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_7 XI11_5/XI0/XI0_33/d__7_ xsel_33_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_6 XI11_5/XI0/XI0_33/d__6_ xsel_33_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_5 XI11_5/XI0/XI0_33/d__5_ xsel_33_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_4 XI11_5/XI0/XI0_33/d__4_ xsel_33_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_3 XI11_5/XI0/XI0_33/d__3_ xsel_33_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_2 XI11_5/XI0/XI0_33/d__2_ xsel_33_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_1 XI11_5/XI0/XI0_33/d__1_ xsel_33_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_0 XI11_5/XI0/XI0_33/d__0_ xsel_33_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_15 XI11_5/net21_0_ xsel_32_ XI11_5/XI0/XI0_32/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_14 XI11_5/net21_1_ xsel_32_ XI11_5/XI0/XI0_32/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_13 XI11_5/net21_2_ xsel_32_ XI11_5/XI0/XI0_32/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_12 XI11_5/net21_3_ xsel_32_ XI11_5/XI0/XI0_32/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_11 XI11_5/net21_4_ xsel_32_ XI11_5/XI0/XI0_32/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_10 XI11_5/net21_5_ xsel_32_ XI11_5/XI0/XI0_32/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_9 XI11_5/net21_6_ xsel_32_ XI11_5/XI0/XI0_32/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_8 XI11_5/net21_7_ xsel_32_ XI11_5/XI0/XI0_32/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_7 XI11_5/net21_8_ xsel_32_ XI11_5/XI0/XI0_32/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_6 XI11_5/net21_9_ xsel_32_ XI11_5/XI0/XI0_32/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_5 XI11_5/net21_10_ xsel_32_ XI11_5/XI0/XI0_32/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_4 XI11_5/net21_11_ xsel_32_ XI11_5/XI0/XI0_32/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_3 XI11_5/net21_12_ xsel_32_ XI11_5/XI0/XI0_32/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_2 XI11_5/net21_13_ xsel_32_ XI11_5/XI0/XI0_32/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_1 XI11_5/net21_14_ xsel_32_ XI11_5/XI0/XI0_32/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_0 XI11_5/net21_15_ xsel_32_ XI11_5/XI0/XI0_32/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_15 XI11_5/XI0/XI0_32/d__15_ xsel_32_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_14 XI11_5/XI0/XI0_32/d__14_ xsel_32_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_13 XI11_5/XI0/XI0_32/d__13_ xsel_32_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_12 XI11_5/XI0/XI0_32/d__12_ xsel_32_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_11 XI11_5/XI0/XI0_32/d__11_ xsel_32_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_10 XI11_5/XI0/XI0_32/d__10_ xsel_32_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_9 XI11_5/XI0/XI0_32/d__9_ xsel_32_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_8 XI11_5/XI0/XI0_32/d__8_ xsel_32_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_7 XI11_5/XI0/XI0_32/d__7_ xsel_32_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_6 XI11_5/XI0/XI0_32/d__6_ xsel_32_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_5 XI11_5/XI0/XI0_32/d__5_ xsel_32_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_4 XI11_5/XI0/XI0_32/d__4_ xsel_32_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_3 XI11_5/XI0/XI0_32/d__3_ xsel_32_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_2 XI11_5/XI0/XI0_32/d__2_ xsel_32_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_1 XI11_5/XI0/XI0_32/d__1_ xsel_32_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_0 XI11_5/XI0/XI0_32/d__0_ xsel_32_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_15 XI11_5/net21_0_ xsel_31_ XI11_5/XI0/XI0_31/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_14 XI11_5/net21_1_ xsel_31_ XI11_5/XI0/XI0_31/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_13 XI11_5/net21_2_ xsel_31_ XI11_5/XI0/XI0_31/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_12 XI11_5/net21_3_ xsel_31_ XI11_5/XI0/XI0_31/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_11 XI11_5/net21_4_ xsel_31_ XI11_5/XI0/XI0_31/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_10 XI11_5/net21_5_ xsel_31_ XI11_5/XI0/XI0_31/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_9 XI11_5/net21_6_ xsel_31_ XI11_5/XI0/XI0_31/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_8 XI11_5/net21_7_ xsel_31_ XI11_5/XI0/XI0_31/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_7 XI11_5/net21_8_ xsel_31_ XI11_5/XI0/XI0_31/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_6 XI11_5/net21_9_ xsel_31_ XI11_5/XI0/XI0_31/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_5 XI11_5/net21_10_ xsel_31_ XI11_5/XI0/XI0_31/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_4 XI11_5/net21_11_ xsel_31_ XI11_5/XI0/XI0_31/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_3 XI11_5/net21_12_ xsel_31_ XI11_5/XI0/XI0_31/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_2 XI11_5/net21_13_ xsel_31_ XI11_5/XI0/XI0_31/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_1 XI11_5/net21_14_ xsel_31_ XI11_5/XI0/XI0_31/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_0 XI11_5/net21_15_ xsel_31_ XI11_5/XI0/XI0_31/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_15 XI11_5/XI0/XI0_31/d__15_ xsel_31_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_14 XI11_5/XI0/XI0_31/d__14_ xsel_31_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_13 XI11_5/XI0/XI0_31/d__13_ xsel_31_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_12 XI11_5/XI0/XI0_31/d__12_ xsel_31_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_11 XI11_5/XI0/XI0_31/d__11_ xsel_31_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_10 XI11_5/XI0/XI0_31/d__10_ xsel_31_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_9 XI11_5/XI0/XI0_31/d__9_ xsel_31_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_8 XI11_5/XI0/XI0_31/d__8_ xsel_31_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_7 XI11_5/XI0/XI0_31/d__7_ xsel_31_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_6 XI11_5/XI0/XI0_31/d__6_ xsel_31_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_5 XI11_5/XI0/XI0_31/d__5_ xsel_31_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_4 XI11_5/XI0/XI0_31/d__4_ xsel_31_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_3 XI11_5/XI0/XI0_31/d__3_ xsel_31_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_2 XI11_5/XI0/XI0_31/d__2_ xsel_31_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_1 XI11_5/XI0/XI0_31/d__1_ xsel_31_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_0 XI11_5/XI0/XI0_31/d__0_ xsel_31_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_15 XI11_5/net21_0_ xsel_30_ XI11_5/XI0/XI0_30/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_14 XI11_5/net21_1_ xsel_30_ XI11_5/XI0/XI0_30/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_13 XI11_5/net21_2_ xsel_30_ XI11_5/XI0/XI0_30/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_12 XI11_5/net21_3_ xsel_30_ XI11_5/XI0/XI0_30/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_11 XI11_5/net21_4_ xsel_30_ XI11_5/XI0/XI0_30/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_10 XI11_5/net21_5_ xsel_30_ XI11_5/XI0/XI0_30/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_9 XI11_5/net21_6_ xsel_30_ XI11_5/XI0/XI0_30/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_8 XI11_5/net21_7_ xsel_30_ XI11_5/XI0/XI0_30/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_7 XI11_5/net21_8_ xsel_30_ XI11_5/XI0/XI0_30/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_6 XI11_5/net21_9_ xsel_30_ XI11_5/XI0/XI0_30/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_5 XI11_5/net21_10_ xsel_30_ XI11_5/XI0/XI0_30/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_4 XI11_5/net21_11_ xsel_30_ XI11_5/XI0/XI0_30/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_3 XI11_5/net21_12_ xsel_30_ XI11_5/XI0/XI0_30/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_2 XI11_5/net21_13_ xsel_30_ XI11_5/XI0/XI0_30/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_1 XI11_5/net21_14_ xsel_30_ XI11_5/XI0/XI0_30/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_0 XI11_5/net21_15_ xsel_30_ XI11_5/XI0/XI0_30/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_15 XI11_5/XI0/XI0_30/d__15_ xsel_30_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_14 XI11_5/XI0/XI0_30/d__14_ xsel_30_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_13 XI11_5/XI0/XI0_30/d__13_ xsel_30_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_12 XI11_5/XI0/XI0_30/d__12_ xsel_30_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_11 XI11_5/XI0/XI0_30/d__11_ xsel_30_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_10 XI11_5/XI0/XI0_30/d__10_ xsel_30_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_9 XI11_5/XI0/XI0_30/d__9_ xsel_30_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_8 XI11_5/XI0/XI0_30/d__8_ xsel_30_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_7 XI11_5/XI0/XI0_30/d__7_ xsel_30_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_6 XI11_5/XI0/XI0_30/d__6_ xsel_30_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_5 XI11_5/XI0/XI0_30/d__5_ xsel_30_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_4 XI11_5/XI0/XI0_30/d__4_ xsel_30_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_3 XI11_5/XI0/XI0_30/d__3_ xsel_30_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_2 XI11_5/XI0/XI0_30/d__2_ xsel_30_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_1 XI11_5/XI0/XI0_30/d__1_ xsel_30_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_0 XI11_5/XI0/XI0_30/d__0_ xsel_30_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_15 XI11_5/net21_0_ xsel_29_ XI11_5/XI0/XI0_29/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_14 XI11_5/net21_1_ xsel_29_ XI11_5/XI0/XI0_29/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_13 XI11_5/net21_2_ xsel_29_ XI11_5/XI0/XI0_29/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_12 XI11_5/net21_3_ xsel_29_ XI11_5/XI0/XI0_29/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_11 XI11_5/net21_4_ xsel_29_ XI11_5/XI0/XI0_29/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_10 XI11_5/net21_5_ xsel_29_ XI11_5/XI0/XI0_29/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_9 XI11_5/net21_6_ xsel_29_ XI11_5/XI0/XI0_29/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_8 XI11_5/net21_7_ xsel_29_ XI11_5/XI0/XI0_29/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_7 XI11_5/net21_8_ xsel_29_ XI11_5/XI0/XI0_29/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_6 XI11_5/net21_9_ xsel_29_ XI11_5/XI0/XI0_29/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_5 XI11_5/net21_10_ xsel_29_ XI11_5/XI0/XI0_29/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_4 XI11_5/net21_11_ xsel_29_ XI11_5/XI0/XI0_29/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_3 XI11_5/net21_12_ xsel_29_ XI11_5/XI0/XI0_29/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_2 XI11_5/net21_13_ xsel_29_ XI11_5/XI0/XI0_29/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_1 XI11_5/net21_14_ xsel_29_ XI11_5/XI0/XI0_29/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_0 XI11_5/net21_15_ xsel_29_ XI11_5/XI0/XI0_29/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_15 XI11_5/XI0/XI0_29/d__15_ xsel_29_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_14 XI11_5/XI0/XI0_29/d__14_ xsel_29_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_13 XI11_5/XI0/XI0_29/d__13_ xsel_29_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_12 XI11_5/XI0/XI0_29/d__12_ xsel_29_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_11 XI11_5/XI0/XI0_29/d__11_ xsel_29_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_10 XI11_5/XI0/XI0_29/d__10_ xsel_29_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_9 XI11_5/XI0/XI0_29/d__9_ xsel_29_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_8 XI11_5/XI0/XI0_29/d__8_ xsel_29_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_7 XI11_5/XI0/XI0_29/d__7_ xsel_29_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_6 XI11_5/XI0/XI0_29/d__6_ xsel_29_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_5 XI11_5/XI0/XI0_29/d__5_ xsel_29_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_4 XI11_5/XI0/XI0_29/d__4_ xsel_29_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_3 XI11_5/XI0/XI0_29/d__3_ xsel_29_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_2 XI11_5/XI0/XI0_29/d__2_ xsel_29_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_1 XI11_5/XI0/XI0_29/d__1_ xsel_29_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_0 XI11_5/XI0/XI0_29/d__0_ xsel_29_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_15 XI11_5/net21_0_ xsel_28_ XI11_5/XI0/XI0_28/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_14 XI11_5/net21_1_ xsel_28_ XI11_5/XI0/XI0_28/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_13 XI11_5/net21_2_ xsel_28_ XI11_5/XI0/XI0_28/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_12 XI11_5/net21_3_ xsel_28_ XI11_5/XI0/XI0_28/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_11 XI11_5/net21_4_ xsel_28_ XI11_5/XI0/XI0_28/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_10 XI11_5/net21_5_ xsel_28_ XI11_5/XI0/XI0_28/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_9 XI11_5/net21_6_ xsel_28_ XI11_5/XI0/XI0_28/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_8 XI11_5/net21_7_ xsel_28_ XI11_5/XI0/XI0_28/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_7 XI11_5/net21_8_ xsel_28_ XI11_5/XI0/XI0_28/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_6 XI11_5/net21_9_ xsel_28_ XI11_5/XI0/XI0_28/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_5 XI11_5/net21_10_ xsel_28_ XI11_5/XI0/XI0_28/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_4 XI11_5/net21_11_ xsel_28_ XI11_5/XI0/XI0_28/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_3 XI11_5/net21_12_ xsel_28_ XI11_5/XI0/XI0_28/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_2 XI11_5/net21_13_ xsel_28_ XI11_5/XI0/XI0_28/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_1 XI11_5/net21_14_ xsel_28_ XI11_5/XI0/XI0_28/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_0 XI11_5/net21_15_ xsel_28_ XI11_5/XI0/XI0_28/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_15 XI11_5/XI0/XI0_28/d__15_ xsel_28_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_14 XI11_5/XI0/XI0_28/d__14_ xsel_28_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_13 XI11_5/XI0/XI0_28/d__13_ xsel_28_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_12 XI11_5/XI0/XI0_28/d__12_ xsel_28_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_11 XI11_5/XI0/XI0_28/d__11_ xsel_28_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_10 XI11_5/XI0/XI0_28/d__10_ xsel_28_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_9 XI11_5/XI0/XI0_28/d__9_ xsel_28_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_8 XI11_5/XI0/XI0_28/d__8_ xsel_28_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_7 XI11_5/XI0/XI0_28/d__7_ xsel_28_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_6 XI11_5/XI0/XI0_28/d__6_ xsel_28_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_5 XI11_5/XI0/XI0_28/d__5_ xsel_28_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_4 XI11_5/XI0/XI0_28/d__4_ xsel_28_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_3 XI11_5/XI0/XI0_28/d__3_ xsel_28_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_2 XI11_5/XI0/XI0_28/d__2_ xsel_28_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_1 XI11_5/XI0/XI0_28/d__1_ xsel_28_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_0 XI11_5/XI0/XI0_28/d__0_ xsel_28_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_15 XI11_5/net21_0_ xsel_27_ XI11_5/XI0/XI0_27/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_14 XI11_5/net21_1_ xsel_27_ XI11_5/XI0/XI0_27/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_13 XI11_5/net21_2_ xsel_27_ XI11_5/XI0/XI0_27/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_12 XI11_5/net21_3_ xsel_27_ XI11_5/XI0/XI0_27/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_11 XI11_5/net21_4_ xsel_27_ XI11_5/XI0/XI0_27/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_10 XI11_5/net21_5_ xsel_27_ XI11_5/XI0/XI0_27/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_9 XI11_5/net21_6_ xsel_27_ XI11_5/XI0/XI0_27/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_8 XI11_5/net21_7_ xsel_27_ XI11_5/XI0/XI0_27/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_7 XI11_5/net21_8_ xsel_27_ XI11_5/XI0/XI0_27/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_6 XI11_5/net21_9_ xsel_27_ XI11_5/XI0/XI0_27/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_5 XI11_5/net21_10_ xsel_27_ XI11_5/XI0/XI0_27/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_4 XI11_5/net21_11_ xsel_27_ XI11_5/XI0/XI0_27/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_3 XI11_5/net21_12_ xsel_27_ XI11_5/XI0/XI0_27/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_2 XI11_5/net21_13_ xsel_27_ XI11_5/XI0/XI0_27/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_1 XI11_5/net21_14_ xsel_27_ XI11_5/XI0/XI0_27/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_0 XI11_5/net21_15_ xsel_27_ XI11_5/XI0/XI0_27/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_15 XI11_5/XI0/XI0_27/d__15_ xsel_27_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_14 XI11_5/XI0/XI0_27/d__14_ xsel_27_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_13 XI11_5/XI0/XI0_27/d__13_ xsel_27_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_12 XI11_5/XI0/XI0_27/d__12_ xsel_27_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_11 XI11_5/XI0/XI0_27/d__11_ xsel_27_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_10 XI11_5/XI0/XI0_27/d__10_ xsel_27_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_9 XI11_5/XI0/XI0_27/d__9_ xsel_27_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_8 XI11_5/XI0/XI0_27/d__8_ xsel_27_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_7 XI11_5/XI0/XI0_27/d__7_ xsel_27_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_6 XI11_5/XI0/XI0_27/d__6_ xsel_27_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_5 XI11_5/XI0/XI0_27/d__5_ xsel_27_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_4 XI11_5/XI0/XI0_27/d__4_ xsel_27_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_3 XI11_5/XI0/XI0_27/d__3_ xsel_27_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_2 XI11_5/XI0/XI0_27/d__2_ xsel_27_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_1 XI11_5/XI0/XI0_27/d__1_ xsel_27_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_0 XI11_5/XI0/XI0_27/d__0_ xsel_27_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_15 XI11_5/net21_0_ xsel_26_ XI11_5/XI0/XI0_26/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_14 XI11_5/net21_1_ xsel_26_ XI11_5/XI0/XI0_26/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_13 XI11_5/net21_2_ xsel_26_ XI11_5/XI0/XI0_26/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_12 XI11_5/net21_3_ xsel_26_ XI11_5/XI0/XI0_26/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_11 XI11_5/net21_4_ xsel_26_ XI11_5/XI0/XI0_26/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_10 XI11_5/net21_5_ xsel_26_ XI11_5/XI0/XI0_26/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_9 XI11_5/net21_6_ xsel_26_ XI11_5/XI0/XI0_26/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_8 XI11_5/net21_7_ xsel_26_ XI11_5/XI0/XI0_26/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_7 XI11_5/net21_8_ xsel_26_ XI11_5/XI0/XI0_26/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_6 XI11_5/net21_9_ xsel_26_ XI11_5/XI0/XI0_26/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_5 XI11_5/net21_10_ xsel_26_ XI11_5/XI0/XI0_26/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_4 XI11_5/net21_11_ xsel_26_ XI11_5/XI0/XI0_26/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_3 XI11_5/net21_12_ xsel_26_ XI11_5/XI0/XI0_26/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_2 XI11_5/net21_13_ xsel_26_ XI11_5/XI0/XI0_26/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_1 XI11_5/net21_14_ xsel_26_ XI11_5/XI0/XI0_26/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_0 XI11_5/net21_15_ xsel_26_ XI11_5/XI0/XI0_26/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_15 XI11_5/XI0/XI0_26/d__15_ xsel_26_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_14 XI11_5/XI0/XI0_26/d__14_ xsel_26_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_13 XI11_5/XI0/XI0_26/d__13_ xsel_26_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_12 XI11_5/XI0/XI0_26/d__12_ xsel_26_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_11 XI11_5/XI0/XI0_26/d__11_ xsel_26_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_10 XI11_5/XI0/XI0_26/d__10_ xsel_26_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_9 XI11_5/XI0/XI0_26/d__9_ xsel_26_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_8 XI11_5/XI0/XI0_26/d__8_ xsel_26_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_7 XI11_5/XI0/XI0_26/d__7_ xsel_26_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_6 XI11_5/XI0/XI0_26/d__6_ xsel_26_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_5 XI11_5/XI0/XI0_26/d__5_ xsel_26_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_4 XI11_5/XI0/XI0_26/d__4_ xsel_26_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_3 XI11_5/XI0/XI0_26/d__3_ xsel_26_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_2 XI11_5/XI0/XI0_26/d__2_ xsel_26_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_1 XI11_5/XI0/XI0_26/d__1_ xsel_26_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_0 XI11_5/XI0/XI0_26/d__0_ xsel_26_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_15 XI11_5/net21_0_ xsel_25_ XI11_5/XI0/XI0_25/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_14 XI11_5/net21_1_ xsel_25_ XI11_5/XI0/XI0_25/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_13 XI11_5/net21_2_ xsel_25_ XI11_5/XI0/XI0_25/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_12 XI11_5/net21_3_ xsel_25_ XI11_5/XI0/XI0_25/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_11 XI11_5/net21_4_ xsel_25_ XI11_5/XI0/XI0_25/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_10 XI11_5/net21_5_ xsel_25_ XI11_5/XI0/XI0_25/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_9 XI11_5/net21_6_ xsel_25_ XI11_5/XI0/XI0_25/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_8 XI11_5/net21_7_ xsel_25_ XI11_5/XI0/XI0_25/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_7 XI11_5/net21_8_ xsel_25_ XI11_5/XI0/XI0_25/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_6 XI11_5/net21_9_ xsel_25_ XI11_5/XI0/XI0_25/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_5 XI11_5/net21_10_ xsel_25_ XI11_5/XI0/XI0_25/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_4 XI11_5/net21_11_ xsel_25_ XI11_5/XI0/XI0_25/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_3 XI11_5/net21_12_ xsel_25_ XI11_5/XI0/XI0_25/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_2 XI11_5/net21_13_ xsel_25_ XI11_5/XI0/XI0_25/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_1 XI11_5/net21_14_ xsel_25_ XI11_5/XI0/XI0_25/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_0 XI11_5/net21_15_ xsel_25_ XI11_5/XI0/XI0_25/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_15 XI11_5/XI0/XI0_25/d__15_ xsel_25_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_14 XI11_5/XI0/XI0_25/d__14_ xsel_25_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_13 XI11_5/XI0/XI0_25/d__13_ xsel_25_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_12 XI11_5/XI0/XI0_25/d__12_ xsel_25_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_11 XI11_5/XI0/XI0_25/d__11_ xsel_25_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_10 XI11_5/XI0/XI0_25/d__10_ xsel_25_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_9 XI11_5/XI0/XI0_25/d__9_ xsel_25_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_8 XI11_5/XI0/XI0_25/d__8_ xsel_25_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_7 XI11_5/XI0/XI0_25/d__7_ xsel_25_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_6 XI11_5/XI0/XI0_25/d__6_ xsel_25_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_5 XI11_5/XI0/XI0_25/d__5_ xsel_25_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_4 XI11_5/XI0/XI0_25/d__4_ xsel_25_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_3 XI11_5/XI0/XI0_25/d__3_ xsel_25_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_2 XI11_5/XI0/XI0_25/d__2_ xsel_25_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_1 XI11_5/XI0/XI0_25/d__1_ xsel_25_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_0 XI11_5/XI0/XI0_25/d__0_ xsel_25_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_15 XI11_5/net21_0_ xsel_24_ XI11_5/XI0/XI0_24/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_14 XI11_5/net21_1_ xsel_24_ XI11_5/XI0/XI0_24/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_13 XI11_5/net21_2_ xsel_24_ XI11_5/XI0/XI0_24/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_12 XI11_5/net21_3_ xsel_24_ XI11_5/XI0/XI0_24/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_11 XI11_5/net21_4_ xsel_24_ XI11_5/XI0/XI0_24/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_10 XI11_5/net21_5_ xsel_24_ XI11_5/XI0/XI0_24/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_9 XI11_5/net21_6_ xsel_24_ XI11_5/XI0/XI0_24/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_8 XI11_5/net21_7_ xsel_24_ XI11_5/XI0/XI0_24/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_7 XI11_5/net21_8_ xsel_24_ XI11_5/XI0/XI0_24/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_6 XI11_5/net21_9_ xsel_24_ XI11_5/XI0/XI0_24/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_5 XI11_5/net21_10_ xsel_24_ XI11_5/XI0/XI0_24/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_4 XI11_5/net21_11_ xsel_24_ XI11_5/XI0/XI0_24/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_3 XI11_5/net21_12_ xsel_24_ XI11_5/XI0/XI0_24/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_2 XI11_5/net21_13_ xsel_24_ XI11_5/XI0/XI0_24/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_1 XI11_5/net21_14_ xsel_24_ XI11_5/XI0/XI0_24/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_0 XI11_5/net21_15_ xsel_24_ XI11_5/XI0/XI0_24/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_15 XI11_5/XI0/XI0_24/d__15_ xsel_24_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_14 XI11_5/XI0/XI0_24/d__14_ xsel_24_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_13 XI11_5/XI0/XI0_24/d__13_ xsel_24_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_12 XI11_5/XI0/XI0_24/d__12_ xsel_24_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_11 XI11_5/XI0/XI0_24/d__11_ xsel_24_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_10 XI11_5/XI0/XI0_24/d__10_ xsel_24_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_9 XI11_5/XI0/XI0_24/d__9_ xsel_24_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_8 XI11_5/XI0/XI0_24/d__8_ xsel_24_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_7 XI11_5/XI0/XI0_24/d__7_ xsel_24_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_6 XI11_5/XI0/XI0_24/d__6_ xsel_24_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_5 XI11_5/XI0/XI0_24/d__5_ xsel_24_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_4 XI11_5/XI0/XI0_24/d__4_ xsel_24_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_3 XI11_5/XI0/XI0_24/d__3_ xsel_24_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_2 XI11_5/XI0/XI0_24/d__2_ xsel_24_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_1 XI11_5/XI0/XI0_24/d__1_ xsel_24_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_0 XI11_5/XI0/XI0_24/d__0_ xsel_24_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_15 XI11_5/net21_0_ xsel_23_ XI11_5/XI0/XI0_23/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_14 XI11_5/net21_1_ xsel_23_ XI11_5/XI0/XI0_23/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_13 XI11_5/net21_2_ xsel_23_ XI11_5/XI0/XI0_23/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_12 XI11_5/net21_3_ xsel_23_ XI11_5/XI0/XI0_23/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_11 XI11_5/net21_4_ xsel_23_ XI11_5/XI0/XI0_23/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_10 XI11_5/net21_5_ xsel_23_ XI11_5/XI0/XI0_23/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_9 XI11_5/net21_6_ xsel_23_ XI11_5/XI0/XI0_23/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_8 XI11_5/net21_7_ xsel_23_ XI11_5/XI0/XI0_23/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_7 XI11_5/net21_8_ xsel_23_ XI11_5/XI0/XI0_23/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_6 XI11_5/net21_9_ xsel_23_ XI11_5/XI0/XI0_23/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_5 XI11_5/net21_10_ xsel_23_ XI11_5/XI0/XI0_23/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_4 XI11_5/net21_11_ xsel_23_ XI11_5/XI0/XI0_23/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_3 XI11_5/net21_12_ xsel_23_ XI11_5/XI0/XI0_23/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_2 XI11_5/net21_13_ xsel_23_ XI11_5/XI0/XI0_23/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_1 XI11_5/net21_14_ xsel_23_ XI11_5/XI0/XI0_23/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_0 XI11_5/net21_15_ xsel_23_ XI11_5/XI0/XI0_23/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_15 XI11_5/XI0/XI0_23/d__15_ xsel_23_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_14 XI11_5/XI0/XI0_23/d__14_ xsel_23_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_13 XI11_5/XI0/XI0_23/d__13_ xsel_23_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_12 XI11_5/XI0/XI0_23/d__12_ xsel_23_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_11 XI11_5/XI0/XI0_23/d__11_ xsel_23_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_10 XI11_5/XI0/XI0_23/d__10_ xsel_23_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_9 XI11_5/XI0/XI0_23/d__9_ xsel_23_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_8 XI11_5/XI0/XI0_23/d__8_ xsel_23_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_7 XI11_5/XI0/XI0_23/d__7_ xsel_23_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_6 XI11_5/XI0/XI0_23/d__6_ xsel_23_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_5 XI11_5/XI0/XI0_23/d__5_ xsel_23_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_4 XI11_5/XI0/XI0_23/d__4_ xsel_23_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_3 XI11_5/XI0/XI0_23/d__3_ xsel_23_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_2 XI11_5/XI0/XI0_23/d__2_ xsel_23_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_1 XI11_5/XI0/XI0_23/d__1_ xsel_23_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_0 XI11_5/XI0/XI0_23/d__0_ xsel_23_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_15 XI11_5/net21_0_ xsel_22_ XI11_5/XI0/XI0_22/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_14 XI11_5/net21_1_ xsel_22_ XI11_5/XI0/XI0_22/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_13 XI11_5/net21_2_ xsel_22_ XI11_5/XI0/XI0_22/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_12 XI11_5/net21_3_ xsel_22_ XI11_5/XI0/XI0_22/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_11 XI11_5/net21_4_ xsel_22_ XI11_5/XI0/XI0_22/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_10 XI11_5/net21_5_ xsel_22_ XI11_5/XI0/XI0_22/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_9 XI11_5/net21_6_ xsel_22_ XI11_5/XI0/XI0_22/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_8 XI11_5/net21_7_ xsel_22_ XI11_5/XI0/XI0_22/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_7 XI11_5/net21_8_ xsel_22_ XI11_5/XI0/XI0_22/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_6 XI11_5/net21_9_ xsel_22_ XI11_5/XI0/XI0_22/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_5 XI11_5/net21_10_ xsel_22_ XI11_5/XI0/XI0_22/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_4 XI11_5/net21_11_ xsel_22_ XI11_5/XI0/XI0_22/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_3 XI11_5/net21_12_ xsel_22_ XI11_5/XI0/XI0_22/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_2 XI11_5/net21_13_ xsel_22_ XI11_5/XI0/XI0_22/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_1 XI11_5/net21_14_ xsel_22_ XI11_5/XI0/XI0_22/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_0 XI11_5/net21_15_ xsel_22_ XI11_5/XI0/XI0_22/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_15 XI11_5/XI0/XI0_22/d__15_ xsel_22_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_14 XI11_5/XI0/XI0_22/d__14_ xsel_22_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_13 XI11_5/XI0/XI0_22/d__13_ xsel_22_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_12 XI11_5/XI0/XI0_22/d__12_ xsel_22_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_11 XI11_5/XI0/XI0_22/d__11_ xsel_22_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_10 XI11_5/XI0/XI0_22/d__10_ xsel_22_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_9 XI11_5/XI0/XI0_22/d__9_ xsel_22_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_8 XI11_5/XI0/XI0_22/d__8_ xsel_22_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_7 XI11_5/XI0/XI0_22/d__7_ xsel_22_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_6 XI11_5/XI0/XI0_22/d__6_ xsel_22_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_5 XI11_5/XI0/XI0_22/d__5_ xsel_22_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_4 XI11_5/XI0/XI0_22/d__4_ xsel_22_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_3 XI11_5/XI0/XI0_22/d__3_ xsel_22_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_2 XI11_5/XI0/XI0_22/d__2_ xsel_22_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_1 XI11_5/XI0/XI0_22/d__1_ xsel_22_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_0 XI11_5/XI0/XI0_22/d__0_ xsel_22_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_15 XI11_5/net21_0_ xsel_21_ XI11_5/XI0/XI0_21/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_14 XI11_5/net21_1_ xsel_21_ XI11_5/XI0/XI0_21/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_13 XI11_5/net21_2_ xsel_21_ XI11_5/XI0/XI0_21/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_12 XI11_5/net21_3_ xsel_21_ XI11_5/XI0/XI0_21/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_11 XI11_5/net21_4_ xsel_21_ XI11_5/XI0/XI0_21/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_10 XI11_5/net21_5_ xsel_21_ XI11_5/XI0/XI0_21/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_9 XI11_5/net21_6_ xsel_21_ XI11_5/XI0/XI0_21/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_8 XI11_5/net21_7_ xsel_21_ XI11_5/XI0/XI0_21/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_7 XI11_5/net21_8_ xsel_21_ XI11_5/XI0/XI0_21/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_6 XI11_5/net21_9_ xsel_21_ XI11_5/XI0/XI0_21/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_5 XI11_5/net21_10_ xsel_21_ XI11_5/XI0/XI0_21/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_4 XI11_5/net21_11_ xsel_21_ XI11_5/XI0/XI0_21/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_3 XI11_5/net21_12_ xsel_21_ XI11_5/XI0/XI0_21/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_2 XI11_5/net21_13_ xsel_21_ XI11_5/XI0/XI0_21/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_1 XI11_5/net21_14_ xsel_21_ XI11_5/XI0/XI0_21/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_0 XI11_5/net21_15_ xsel_21_ XI11_5/XI0/XI0_21/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_15 XI11_5/XI0/XI0_21/d__15_ xsel_21_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_14 XI11_5/XI0/XI0_21/d__14_ xsel_21_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_13 XI11_5/XI0/XI0_21/d__13_ xsel_21_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_12 XI11_5/XI0/XI0_21/d__12_ xsel_21_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_11 XI11_5/XI0/XI0_21/d__11_ xsel_21_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_10 XI11_5/XI0/XI0_21/d__10_ xsel_21_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_9 XI11_5/XI0/XI0_21/d__9_ xsel_21_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_8 XI11_5/XI0/XI0_21/d__8_ xsel_21_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_7 XI11_5/XI0/XI0_21/d__7_ xsel_21_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_6 XI11_5/XI0/XI0_21/d__6_ xsel_21_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_5 XI11_5/XI0/XI0_21/d__5_ xsel_21_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_4 XI11_5/XI0/XI0_21/d__4_ xsel_21_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_3 XI11_5/XI0/XI0_21/d__3_ xsel_21_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_2 XI11_5/XI0/XI0_21/d__2_ xsel_21_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_1 XI11_5/XI0/XI0_21/d__1_ xsel_21_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_0 XI11_5/XI0/XI0_21/d__0_ xsel_21_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_15 XI11_5/net21_0_ xsel_20_ XI11_5/XI0/XI0_20/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_14 XI11_5/net21_1_ xsel_20_ XI11_5/XI0/XI0_20/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_13 XI11_5/net21_2_ xsel_20_ XI11_5/XI0/XI0_20/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_12 XI11_5/net21_3_ xsel_20_ XI11_5/XI0/XI0_20/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_11 XI11_5/net21_4_ xsel_20_ XI11_5/XI0/XI0_20/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_10 XI11_5/net21_5_ xsel_20_ XI11_5/XI0/XI0_20/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_9 XI11_5/net21_6_ xsel_20_ XI11_5/XI0/XI0_20/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_8 XI11_5/net21_7_ xsel_20_ XI11_5/XI0/XI0_20/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_7 XI11_5/net21_8_ xsel_20_ XI11_5/XI0/XI0_20/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_6 XI11_5/net21_9_ xsel_20_ XI11_5/XI0/XI0_20/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_5 XI11_5/net21_10_ xsel_20_ XI11_5/XI0/XI0_20/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_4 XI11_5/net21_11_ xsel_20_ XI11_5/XI0/XI0_20/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_3 XI11_5/net21_12_ xsel_20_ XI11_5/XI0/XI0_20/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_2 XI11_5/net21_13_ xsel_20_ XI11_5/XI0/XI0_20/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_1 XI11_5/net21_14_ xsel_20_ XI11_5/XI0/XI0_20/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_0 XI11_5/net21_15_ xsel_20_ XI11_5/XI0/XI0_20/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_15 XI11_5/XI0/XI0_20/d__15_ xsel_20_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_14 XI11_5/XI0/XI0_20/d__14_ xsel_20_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_13 XI11_5/XI0/XI0_20/d__13_ xsel_20_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_12 XI11_5/XI0/XI0_20/d__12_ xsel_20_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_11 XI11_5/XI0/XI0_20/d__11_ xsel_20_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_10 XI11_5/XI0/XI0_20/d__10_ xsel_20_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_9 XI11_5/XI0/XI0_20/d__9_ xsel_20_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_8 XI11_5/XI0/XI0_20/d__8_ xsel_20_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_7 XI11_5/XI0/XI0_20/d__7_ xsel_20_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_6 XI11_5/XI0/XI0_20/d__6_ xsel_20_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_5 XI11_5/XI0/XI0_20/d__5_ xsel_20_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_4 XI11_5/XI0/XI0_20/d__4_ xsel_20_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_3 XI11_5/XI0/XI0_20/d__3_ xsel_20_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_2 XI11_5/XI0/XI0_20/d__2_ xsel_20_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_1 XI11_5/XI0/XI0_20/d__1_ xsel_20_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_0 XI11_5/XI0/XI0_20/d__0_ xsel_20_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_15 XI11_5/net21_0_ xsel_19_ XI11_5/XI0/XI0_19/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_14 XI11_5/net21_1_ xsel_19_ XI11_5/XI0/XI0_19/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_13 XI11_5/net21_2_ xsel_19_ XI11_5/XI0/XI0_19/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_12 XI11_5/net21_3_ xsel_19_ XI11_5/XI0/XI0_19/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_11 XI11_5/net21_4_ xsel_19_ XI11_5/XI0/XI0_19/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_10 XI11_5/net21_5_ xsel_19_ XI11_5/XI0/XI0_19/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_9 XI11_5/net21_6_ xsel_19_ XI11_5/XI0/XI0_19/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_8 XI11_5/net21_7_ xsel_19_ XI11_5/XI0/XI0_19/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_7 XI11_5/net21_8_ xsel_19_ XI11_5/XI0/XI0_19/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_6 XI11_5/net21_9_ xsel_19_ XI11_5/XI0/XI0_19/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_5 XI11_5/net21_10_ xsel_19_ XI11_5/XI0/XI0_19/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_4 XI11_5/net21_11_ xsel_19_ XI11_5/XI0/XI0_19/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_3 XI11_5/net21_12_ xsel_19_ XI11_5/XI0/XI0_19/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_2 XI11_5/net21_13_ xsel_19_ XI11_5/XI0/XI0_19/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_1 XI11_5/net21_14_ xsel_19_ XI11_5/XI0/XI0_19/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_0 XI11_5/net21_15_ xsel_19_ XI11_5/XI0/XI0_19/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_15 XI11_5/XI0/XI0_19/d__15_ xsel_19_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_14 XI11_5/XI0/XI0_19/d__14_ xsel_19_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_13 XI11_5/XI0/XI0_19/d__13_ xsel_19_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_12 XI11_5/XI0/XI0_19/d__12_ xsel_19_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_11 XI11_5/XI0/XI0_19/d__11_ xsel_19_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_10 XI11_5/XI0/XI0_19/d__10_ xsel_19_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_9 XI11_5/XI0/XI0_19/d__9_ xsel_19_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_8 XI11_5/XI0/XI0_19/d__8_ xsel_19_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_7 XI11_5/XI0/XI0_19/d__7_ xsel_19_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_6 XI11_5/XI0/XI0_19/d__6_ xsel_19_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_5 XI11_5/XI0/XI0_19/d__5_ xsel_19_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_4 XI11_5/XI0/XI0_19/d__4_ xsel_19_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_3 XI11_5/XI0/XI0_19/d__3_ xsel_19_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_2 XI11_5/XI0/XI0_19/d__2_ xsel_19_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_1 XI11_5/XI0/XI0_19/d__1_ xsel_19_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_0 XI11_5/XI0/XI0_19/d__0_ xsel_19_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_15 XI11_5/net21_0_ xsel_18_ XI11_5/XI0/XI0_18/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_14 XI11_5/net21_1_ xsel_18_ XI11_5/XI0/XI0_18/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_13 XI11_5/net21_2_ xsel_18_ XI11_5/XI0/XI0_18/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_12 XI11_5/net21_3_ xsel_18_ XI11_5/XI0/XI0_18/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_11 XI11_5/net21_4_ xsel_18_ XI11_5/XI0/XI0_18/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_10 XI11_5/net21_5_ xsel_18_ XI11_5/XI0/XI0_18/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_9 XI11_5/net21_6_ xsel_18_ XI11_5/XI0/XI0_18/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_8 XI11_5/net21_7_ xsel_18_ XI11_5/XI0/XI0_18/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_7 XI11_5/net21_8_ xsel_18_ XI11_5/XI0/XI0_18/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_6 XI11_5/net21_9_ xsel_18_ XI11_5/XI0/XI0_18/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_5 XI11_5/net21_10_ xsel_18_ XI11_5/XI0/XI0_18/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_4 XI11_5/net21_11_ xsel_18_ XI11_5/XI0/XI0_18/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_3 XI11_5/net21_12_ xsel_18_ XI11_5/XI0/XI0_18/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_2 XI11_5/net21_13_ xsel_18_ XI11_5/XI0/XI0_18/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_1 XI11_5/net21_14_ xsel_18_ XI11_5/XI0/XI0_18/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_0 XI11_5/net21_15_ xsel_18_ XI11_5/XI0/XI0_18/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_15 XI11_5/XI0/XI0_18/d__15_ xsel_18_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_14 XI11_5/XI0/XI0_18/d__14_ xsel_18_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_13 XI11_5/XI0/XI0_18/d__13_ xsel_18_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_12 XI11_5/XI0/XI0_18/d__12_ xsel_18_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_11 XI11_5/XI0/XI0_18/d__11_ xsel_18_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_10 XI11_5/XI0/XI0_18/d__10_ xsel_18_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_9 XI11_5/XI0/XI0_18/d__9_ xsel_18_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_8 XI11_5/XI0/XI0_18/d__8_ xsel_18_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_7 XI11_5/XI0/XI0_18/d__7_ xsel_18_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_6 XI11_5/XI0/XI0_18/d__6_ xsel_18_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_5 XI11_5/XI0/XI0_18/d__5_ xsel_18_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_4 XI11_5/XI0/XI0_18/d__4_ xsel_18_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_3 XI11_5/XI0/XI0_18/d__3_ xsel_18_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_2 XI11_5/XI0/XI0_18/d__2_ xsel_18_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_1 XI11_5/XI0/XI0_18/d__1_ xsel_18_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_0 XI11_5/XI0/XI0_18/d__0_ xsel_18_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_15 XI11_5/net21_0_ xsel_17_ XI11_5/XI0/XI0_17/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_14 XI11_5/net21_1_ xsel_17_ XI11_5/XI0/XI0_17/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_13 XI11_5/net21_2_ xsel_17_ XI11_5/XI0/XI0_17/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_12 XI11_5/net21_3_ xsel_17_ XI11_5/XI0/XI0_17/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_11 XI11_5/net21_4_ xsel_17_ XI11_5/XI0/XI0_17/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_10 XI11_5/net21_5_ xsel_17_ XI11_5/XI0/XI0_17/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_9 XI11_5/net21_6_ xsel_17_ XI11_5/XI0/XI0_17/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_8 XI11_5/net21_7_ xsel_17_ XI11_5/XI0/XI0_17/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_7 XI11_5/net21_8_ xsel_17_ XI11_5/XI0/XI0_17/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_6 XI11_5/net21_9_ xsel_17_ XI11_5/XI0/XI0_17/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_5 XI11_5/net21_10_ xsel_17_ XI11_5/XI0/XI0_17/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_4 XI11_5/net21_11_ xsel_17_ XI11_5/XI0/XI0_17/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_3 XI11_5/net21_12_ xsel_17_ XI11_5/XI0/XI0_17/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_2 XI11_5/net21_13_ xsel_17_ XI11_5/XI0/XI0_17/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_1 XI11_5/net21_14_ xsel_17_ XI11_5/XI0/XI0_17/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_0 XI11_5/net21_15_ xsel_17_ XI11_5/XI0/XI0_17/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_15 XI11_5/XI0/XI0_17/d__15_ xsel_17_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_14 XI11_5/XI0/XI0_17/d__14_ xsel_17_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_13 XI11_5/XI0/XI0_17/d__13_ xsel_17_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_12 XI11_5/XI0/XI0_17/d__12_ xsel_17_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_11 XI11_5/XI0/XI0_17/d__11_ xsel_17_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_10 XI11_5/XI0/XI0_17/d__10_ xsel_17_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_9 XI11_5/XI0/XI0_17/d__9_ xsel_17_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_8 XI11_5/XI0/XI0_17/d__8_ xsel_17_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_7 XI11_5/XI0/XI0_17/d__7_ xsel_17_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_6 XI11_5/XI0/XI0_17/d__6_ xsel_17_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_5 XI11_5/XI0/XI0_17/d__5_ xsel_17_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_4 XI11_5/XI0/XI0_17/d__4_ xsel_17_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_3 XI11_5/XI0/XI0_17/d__3_ xsel_17_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_2 XI11_5/XI0/XI0_17/d__2_ xsel_17_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_1 XI11_5/XI0/XI0_17/d__1_ xsel_17_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_0 XI11_5/XI0/XI0_17/d__0_ xsel_17_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_15 XI11_5/net21_0_ xsel_16_ XI11_5/XI0/XI0_16/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_14 XI11_5/net21_1_ xsel_16_ XI11_5/XI0/XI0_16/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_13 XI11_5/net21_2_ xsel_16_ XI11_5/XI0/XI0_16/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_12 XI11_5/net21_3_ xsel_16_ XI11_5/XI0/XI0_16/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_11 XI11_5/net21_4_ xsel_16_ XI11_5/XI0/XI0_16/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_10 XI11_5/net21_5_ xsel_16_ XI11_5/XI0/XI0_16/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_9 XI11_5/net21_6_ xsel_16_ XI11_5/XI0/XI0_16/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_8 XI11_5/net21_7_ xsel_16_ XI11_5/XI0/XI0_16/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_7 XI11_5/net21_8_ xsel_16_ XI11_5/XI0/XI0_16/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_6 XI11_5/net21_9_ xsel_16_ XI11_5/XI0/XI0_16/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_5 XI11_5/net21_10_ xsel_16_ XI11_5/XI0/XI0_16/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_4 XI11_5/net21_11_ xsel_16_ XI11_5/XI0/XI0_16/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_3 XI11_5/net21_12_ xsel_16_ XI11_5/XI0/XI0_16/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_2 XI11_5/net21_13_ xsel_16_ XI11_5/XI0/XI0_16/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_1 XI11_5/net21_14_ xsel_16_ XI11_5/XI0/XI0_16/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_0 XI11_5/net21_15_ xsel_16_ XI11_5/XI0/XI0_16/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_15 XI11_5/XI0/XI0_16/d__15_ xsel_16_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_14 XI11_5/XI0/XI0_16/d__14_ xsel_16_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_13 XI11_5/XI0/XI0_16/d__13_ xsel_16_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_12 XI11_5/XI0/XI0_16/d__12_ xsel_16_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_11 XI11_5/XI0/XI0_16/d__11_ xsel_16_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_10 XI11_5/XI0/XI0_16/d__10_ xsel_16_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_9 XI11_5/XI0/XI0_16/d__9_ xsel_16_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_8 XI11_5/XI0/XI0_16/d__8_ xsel_16_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_7 XI11_5/XI0/XI0_16/d__7_ xsel_16_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_6 XI11_5/XI0/XI0_16/d__6_ xsel_16_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_5 XI11_5/XI0/XI0_16/d__5_ xsel_16_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_4 XI11_5/XI0/XI0_16/d__4_ xsel_16_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_3 XI11_5/XI0/XI0_16/d__3_ xsel_16_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_2 XI11_5/XI0/XI0_16/d__2_ xsel_16_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_1 XI11_5/XI0/XI0_16/d__1_ xsel_16_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_0 XI11_5/XI0/XI0_16/d__0_ xsel_16_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_15 XI11_5/net21_0_ xsel_15_ XI11_5/XI0/XI0_15/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_14 XI11_5/net21_1_ xsel_15_ XI11_5/XI0/XI0_15/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_13 XI11_5/net21_2_ xsel_15_ XI11_5/XI0/XI0_15/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_12 XI11_5/net21_3_ xsel_15_ XI11_5/XI0/XI0_15/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_11 XI11_5/net21_4_ xsel_15_ XI11_5/XI0/XI0_15/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_10 XI11_5/net21_5_ xsel_15_ XI11_5/XI0/XI0_15/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_9 XI11_5/net21_6_ xsel_15_ XI11_5/XI0/XI0_15/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_8 XI11_5/net21_7_ xsel_15_ XI11_5/XI0/XI0_15/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_7 XI11_5/net21_8_ xsel_15_ XI11_5/XI0/XI0_15/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_6 XI11_5/net21_9_ xsel_15_ XI11_5/XI0/XI0_15/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_5 XI11_5/net21_10_ xsel_15_ XI11_5/XI0/XI0_15/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_4 XI11_5/net21_11_ xsel_15_ XI11_5/XI0/XI0_15/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_3 XI11_5/net21_12_ xsel_15_ XI11_5/XI0/XI0_15/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_2 XI11_5/net21_13_ xsel_15_ XI11_5/XI0/XI0_15/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_1 XI11_5/net21_14_ xsel_15_ XI11_5/XI0/XI0_15/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_0 XI11_5/net21_15_ xsel_15_ XI11_5/XI0/XI0_15/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_15 XI11_5/XI0/XI0_15/d__15_ xsel_15_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_14 XI11_5/XI0/XI0_15/d__14_ xsel_15_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_13 XI11_5/XI0/XI0_15/d__13_ xsel_15_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_12 XI11_5/XI0/XI0_15/d__12_ xsel_15_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_11 XI11_5/XI0/XI0_15/d__11_ xsel_15_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_10 XI11_5/XI0/XI0_15/d__10_ xsel_15_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_9 XI11_5/XI0/XI0_15/d__9_ xsel_15_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_8 XI11_5/XI0/XI0_15/d__8_ xsel_15_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_7 XI11_5/XI0/XI0_15/d__7_ xsel_15_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_6 XI11_5/XI0/XI0_15/d__6_ xsel_15_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_5 XI11_5/XI0/XI0_15/d__5_ xsel_15_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_4 XI11_5/XI0/XI0_15/d__4_ xsel_15_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_3 XI11_5/XI0/XI0_15/d__3_ xsel_15_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_2 XI11_5/XI0/XI0_15/d__2_ xsel_15_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_1 XI11_5/XI0/XI0_15/d__1_ xsel_15_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_0 XI11_5/XI0/XI0_15/d__0_ xsel_15_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_15 XI11_5/net21_0_ xsel_14_ XI11_5/XI0/XI0_14/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_14 XI11_5/net21_1_ xsel_14_ XI11_5/XI0/XI0_14/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_13 XI11_5/net21_2_ xsel_14_ XI11_5/XI0/XI0_14/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_12 XI11_5/net21_3_ xsel_14_ XI11_5/XI0/XI0_14/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_11 XI11_5/net21_4_ xsel_14_ XI11_5/XI0/XI0_14/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_10 XI11_5/net21_5_ xsel_14_ XI11_5/XI0/XI0_14/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_9 XI11_5/net21_6_ xsel_14_ XI11_5/XI0/XI0_14/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_8 XI11_5/net21_7_ xsel_14_ XI11_5/XI0/XI0_14/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_7 XI11_5/net21_8_ xsel_14_ XI11_5/XI0/XI0_14/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_6 XI11_5/net21_9_ xsel_14_ XI11_5/XI0/XI0_14/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_5 XI11_5/net21_10_ xsel_14_ XI11_5/XI0/XI0_14/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_4 XI11_5/net21_11_ xsel_14_ XI11_5/XI0/XI0_14/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_3 XI11_5/net21_12_ xsel_14_ XI11_5/XI0/XI0_14/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_2 XI11_5/net21_13_ xsel_14_ XI11_5/XI0/XI0_14/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_1 XI11_5/net21_14_ xsel_14_ XI11_5/XI0/XI0_14/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_0 XI11_5/net21_15_ xsel_14_ XI11_5/XI0/XI0_14/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_15 XI11_5/XI0/XI0_14/d__15_ xsel_14_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_14 XI11_5/XI0/XI0_14/d__14_ xsel_14_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_13 XI11_5/XI0/XI0_14/d__13_ xsel_14_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_12 XI11_5/XI0/XI0_14/d__12_ xsel_14_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_11 XI11_5/XI0/XI0_14/d__11_ xsel_14_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_10 XI11_5/XI0/XI0_14/d__10_ xsel_14_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_9 XI11_5/XI0/XI0_14/d__9_ xsel_14_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_8 XI11_5/XI0/XI0_14/d__8_ xsel_14_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_7 XI11_5/XI0/XI0_14/d__7_ xsel_14_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_6 XI11_5/XI0/XI0_14/d__6_ xsel_14_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_5 XI11_5/XI0/XI0_14/d__5_ xsel_14_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_4 XI11_5/XI0/XI0_14/d__4_ xsel_14_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_3 XI11_5/XI0/XI0_14/d__3_ xsel_14_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_2 XI11_5/XI0/XI0_14/d__2_ xsel_14_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_1 XI11_5/XI0/XI0_14/d__1_ xsel_14_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_0 XI11_5/XI0/XI0_14/d__0_ xsel_14_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_15 XI11_5/net21_0_ xsel_13_ XI11_5/XI0/XI0_13/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_14 XI11_5/net21_1_ xsel_13_ XI11_5/XI0/XI0_13/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_13 XI11_5/net21_2_ xsel_13_ XI11_5/XI0/XI0_13/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_12 XI11_5/net21_3_ xsel_13_ XI11_5/XI0/XI0_13/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_11 XI11_5/net21_4_ xsel_13_ XI11_5/XI0/XI0_13/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_10 XI11_5/net21_5_ xsel_13_ XI11_5/XI0/XI0_13/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_9 XI11_5/net21_6_ xsel_13_ XI11_5/XI0/XI0_13/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_8 XI11_5/net21_7_ xsel_13_ XI11_5/XI0/XI0_13/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_7 XI11_5/net21_8_ xsel_13_ XI11_5/XI0/XI0_13/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_6 XI11_5/net21_9_ xsel_13_ XI11_5/XI0/XI0_13/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_5 XI11_5/net21_10_ xsel_13_ XI11_5/XI0/XI0_13/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_4 XI11_5/net21_11_ xsel_13_ XI11_5/XI0/XI0_13/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_3 XI11_5/net21_12_ xsel_13_ XI11_5/XI0/XI0_13/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_2 XI11_5/net21_13_ xsel_13_ XI11_5/XI0/XI0_13/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_1 XI11_5/net21_14_ xsel_13_ XI11_5/XI0/XI0_13/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_0 XI11_5/net21_15_ xsel_13_ XI11_5/XI0/XI0_13/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_15 XI11_5/XI0/XI0_13/d__15_ xsel_13_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_14 XI11_5/XI0/XI0_13/d__14_ xsel_13_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_13 XI11_5/XI0/XI0_13/d__13_ xsel_13_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_12 XI11_5/XI0/XI0_13/d__12_ xsel_13_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_11 XI11_5/XI0/XI0_13/d__11_ xsel_13_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_10 XI11_5/XI0/XI0_13/d__10_ xsel_13_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_9 XI11_5/XI0/XI0_13/d__9_ xsel_13_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_8 XI11_5/XI0/XI0_13/d__8_ xsel_13_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_7 XI11_5/XI0/XI0_13/d__7_ xsel_13_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_6 XI11_5/XI0/XI0_13/d__6_ xsel_13_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_5 XI11_5/XI0/XI0_13/d__5_ xsel_13_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_4 XI11_5/XI0/XI0_13/d__4_ xsel_13_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_3 XI11_5/XI0/XI0_13/d__3_ xsel_13_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_2 XI11_5/XI0/XI0_13/d__2_ xsel_13_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_1 XI11_5/XI0/XI0_13/d__1_ xsel_13_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_0 XI11_5/XI0/XI0_13/d__0_ xsel_13_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_15 XI11_5/net21_0_ xsel_12_ XI11_5/XI0/XI0_12/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_14 XI11_5/net21_1_ xsel_12_ XI11_5/XI0/XI0_12/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_13 XI11_5/net21_2_ xsel_12_ XI11_5/XI0/XI0_12/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_12 XI11_5/net21_3_ xsel_12_ XI11_5/XI0/XI0_12/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_11 XI11_5/net21_4_ xsel_12_ XI11_5/XI0/XI0_12/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_10 XI11_5/net21_5_ xsel_12_ XI11_5/XI0/XI0_12/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_9 XI11_5/net21_6_ xsel_12_ XI11_5/XI0/XI0_12/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_8 XI11_5/net21_7_ xsel_12_ XI11_5/XI0/XI0_12/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_7 XI11_5/net21_8_ xsel_12_ XI11_5/XI0/XI0_12/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_6 XI11_5/net21_9_ xsel_12_ XI11_5/XI0/XI0_12/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_5 XI11_5/net21_10_ xsel_12_ XI11_5/XI0/XI0_12/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_4 XI11_5/net21_11_ xsel_12_ XI11_5/XI0/XI0_12/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_3 XI11_5/net21_12_ xsel_12_ XI11_5/XI0/XI0_12/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_2 XI11_5/net21_13_ xsel_12_ XI11_5/XI0/XI0_12/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_1 XI11_5/net21_14_ xsel_12_ XI11_5/XI0/XI0_12/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_0 XI11_5/net21_15_ xsel_12_ XI11_5/XI0/XI0_12/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_15 XI11_5/XI0/XI0_12/d__15_ xsel_12_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_14 XI11_5/XI0/XI0_12/d__14_ xsel_12_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_13 XI11_5/XI0/XI0_12/d__13_ xsel_12_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_12 XI11_5/XI0/XI0_12/d__12_ xsel_12_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_11 XI11_5/XI0/XI0_12/d__11_ xsel_12_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_10 XI11_5/XI0/XI0_12/d__10_ xsel_12_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_9 XI11_5/XI0/XI0_12/d__9_ xsel_12_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_8 XI11_5/XI0/XI0_12/d__8_ xsel_12_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_7 XI11_5/XI0/XI0_12/d__7_ xsel_12_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_6 XI11_5/XI0/XI0_12/d__6_ xsel_12_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_5 XI11_5/XI0/XI0_12/d__5_ xsel_12_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_4 XI11_5/XI0/XI0_12/d__4_ xsel_12_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_3 XI11_5/XI0/XI0_12/d__3_ xsel_12_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_2 XI11_5/XI0/XI0_12/d__2_ xsel_12_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_1 XI11_5/XI0/XI0_12/d__1_ xsel_12_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_0 XI11_5/XI0/XI0_12/d__0_ xsel_12_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_15 XI11_5/net21_0_ xsel_11_ XI11_5/XI0/XI0_11/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_14 XI11_5/net21_1_ xsel_11_ XI11_5/XI0/XI0_11/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_13 XI11_5/net21_2_ xsel_11_ XI11_5/XI0/XI0_11/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_12 XI11_5/net21_3_ xsel_11_ XI11_5/XI0/XI0_11/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_11 XI11_5/net21_4_ xsel_11_ XI11_5/XI0/XI0_11/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_10 XI11_5/net21_5_ xsel_11_ XI11_5/XI0/XI0_11/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_9 XI11_5/net21_6_ xsel_11_ XI11_5/XI0/XI0_11/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_8 XI11_5/net21_7_ xsel_11_ XI11_5/XI0/XI0_11/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_7 XI11_5/net21_8_ xsel_11_ XI11_5/XI0/XI0_11/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_6 XI11_5/net21_9_ xsel_11_ XI11_5/XI0/XI0_11/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_5 XI11_5/net21_10_ xsel_11_ XI11_5/XI0/XI0_11/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_4 XI11_5/net21_11_ xsel_11_ XI11_5/XI0/XI0_11/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_3 XI11_5/net21_12_ xsel_11_ XI11_5/XI0/XI0_11/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_2 XI11_5/net21_13_ xsel_11_ XI11_5/XI0/XI0_11/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_1 XI11_5/net21_14_ xsel_11_ XI11_5/XI0/XI0_11/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_0 XI11_5/net21_15_ xsel_11_ XI11_5/XI0/XI0_11/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_15 XI11_5/XI0/XI0_11/d__15_ xsel_11_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_14 XI11_5/XI0/XI0_11/d__14_ xsel_11_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_13 XI11_5/XI0/XI0_11/d__13_ xsel_11_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_12 XI11_5/XI0/XI0_11/d__12_ xsel_11_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_11 XI11_5/XI0/XI0_11/d__11_ xsel_11_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_10 XI11_5/XI0/XI0_11/d__10_ xsel_11_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_9 XI11_5/XI0/XI0_11/d__9_ xsel_11_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_8 XI11_5/XI0/XI0_11/d__8_ xsel_11_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_7 XI11_5/XI0/XI0_11/d__7_ xsel_11_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_6 XI11_5/XI0/XI0_11/d__6_ xsel_11_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_5 XI11_5/XI0/XI0_11/d__5_ xsel_11_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_4 XI11_5/XI0/XI0_11/d__4_ xsel_11_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_3 XI11_5/XI0/XI0_11/d__3_ xsel_11_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_2 XI11_5/XI0/XI0_11/d__2_ xsel_11_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_1 XI11_5/XI0/XI0_11/d__1_ xsel_11_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_0 XI11_5/XI0/XI0_11/d__0_ xsel_11_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_15 XI11_5/net21_0_ xsel_10_ XI11_5/XI0/XI0_10/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_14 XI11_5/net21_1_ xsel_10_ XI11_5/XI0/XI0_10/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_13 XI11_5/net21_2_ xsel_10_ XI11_5/XI0/XI0_10/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_12 XI11_5/net21_3_ xsel_10_ XI11_5/XI0/XI0_10/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_11 XI11_5/net21_4_ xsel_10_ XI11_5/XI0/XI0_10/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_10 XI11_5/net21_5_ xsel_10_ XI11_5/XI0/XI0_10/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_9 XI11_5/net21_6_ xsel_10_ XI11_5/XI0/XI0_10/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_8 XI11_5/net21_7_ xsel_10_ XI11_5/XI0/XI0_10/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_7 XI11_5/net21_8_ xsel_10_ XI11_5/XI0/XI0_10/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_6 XI11_5/net21_9_ xsel_10_ XI11_5/XI0/XI0_10/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_5 XI11_5/net21_10_ xsel_10_ XI11_5/XI0/XI0_10/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_4 XI11_5/net21_11_ xsel_10_ XI11_5/XI0/XI0_10/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_3 XI11_5/net21_12_ xsel_10_ XI11_5/XI0/XI0_10/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_2 XI11_5/net21_13_ xsel_10_ XI11_5/XI0/XI0_10/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_1 XI11_5/net21_14_ xsel_10_ XI11_5/XI0/XI0_10/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_0 XI11_5/net21_15_ xsel_10_ XI11_5/XI0/XI0_10/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_15 XI11_5/XI0/XI0_10/d__15_ xsel_10_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_14 XI11_5/XI0/XI0_10/d__14_ xsel_10_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_13 XI11_5/XI0/XI0_10/d__13_ xsel_10_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_12 XI11_5/XI0/XI0_10/d__12_ xsel_10_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_11 XI11_5/XI0/XI0_10/d__11_ xsel_10_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_10 XI11_5/XI0/XI0_10/d__10_ xsel_10_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_9 XI11_5/XI0/XI0_10/d__9_ xsel_10_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_8 XI11_5/XI0/XI0_10/d__8_ xsel_10_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_7 XI11_5/XI0/XI0_10/d__7_ xsel_10_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_6 XI11_5/XI0/XI0_10/d__6_ xsel_10_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_5 XI11_5/XI0/XI0_10/d__5_ xsel_10_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_4 XI11_5/XI0/XI0_10/d__4_ xsel_10_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_3 XI11_5/XI0/XI0_10/d__3_ xsel_10_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_2 XI11_5/XI0/XI0_10/d__2_ xsel_10_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_1 XI11_5/XI0/XI0_10/d__1_ xsel_10_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_0 XI11_5/XI0/XI0_10/d__0_ xsel_10_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_15 XI11_5/net21_0_ xsel_9_ XI11_5/XI0/XI0_9/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_14 XI11_5/net21_1_ xsel_9_ XI11_5/XI0/XI0_9/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_13 XI11_5/net21_2_ xsel_9_ XI11_5/XI0/XI0_9/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_12 XI11_5/net21_3_ xsel_9_ XI11_5/XI0/XI0_9/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_11 XI11_5/net21_4_ xsel_9_ XI11_5/XI0/XI0_9/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_10 XI11_5/net21_5_ xsel_9_ XI11_5/XI0/XI0_9/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_9 XI11_5/net21_6_ xsel_9_ XI11_5/XI0/XI0_9/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_8 XI11_5/net21_7_ xsel_9_ XI11_5/XI0/XI0_9/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_7 XI11_5/net21_8_ xsel_9_ XI11_5/XI0/XI0_9/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_6 XI11_5/net21_9_ xsel_9_ XI11_5/XI0/XI0_9/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_5 XI11_5/net21_10_ xsel_9_ XI11_5/XI0/XI0_9/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_4 XI11_5/net21_11_ xsel_9_ XI11_5/XI0/XI0_9/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_3 XI11_5/net21_12_ xsel_9_ XI11_5/XI0/XI0_9/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_2 XI11_5/net21_13_ xsel_9_ XI11_5/XI0/XI0_9/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_1 XI11_5/net21_14_ xsel_9_ XI11_5/XI0/XI0_9/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_0 XI11_5/net21_15_ xsel_9_ XI11_5/XI0/XI0_9/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_15 XI11_5/XI0/XI0_9/d__15_ xsel_9_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_14 XI11_5/XI0/XI0_9/d__14_ xsel_9_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_13 XI11_5/XI0/XI0_9/d__13_ xsel_9_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_12 XI11_5/XI0/XI0_9/d__12_ xsel_9_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_11 XI11_5/XI0/XI0_9/d__11_ xsel_9_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_10 XI11_5/XI0/XI0_9/d__10_ xsel_9_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_9 XI11_5/XI0/XI0_9/d__9_ xsel_9_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_8 XI11_5/XI0/XI0_9/d__8_ xsel_9_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_7 XI11_5/XI0/XI0_9/d__7_ xsel_9_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_6 XI11_5/XI0/XI0_9/d__6_ xsel_9_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_5 XI11_5/XI0/XI0_9/d__5_ xsel_9_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_4 XI11_5/XI0/XI0_9/d__4_ xsel_9_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_3 XI11_5/XI0/XI0_9/d__3_ xsel_9_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_2 XI11_5/XI0/XI0_9/d__2_ xsel_9_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_1 XI11_5/XI0/XI0_9/d__1_ xsel_9_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_0 XI11_5/XI0/XI0_9/d__0_ xsel_9_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_15 XI11_5/net21_0_ xsel_8_ XI11_5/XI0/XI0_8/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_14 XI11_5/net21_1_ xsel_8_ XI11_5/XI0/XI0_8/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_13 XI11_5/net21_2_ xsel_8_ XI11_5/XI0/XI0_8/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_12 XI11_5/net21_3_ xsel_8_ XI11_5/XI0/XI0_8/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_11 XI11_5/net21_4_ xsel_8_ XI11_5/XI0/XI0_8/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_10 XI11_5/net21_5_ xsel_8_ XI11_5/XI0/XI0_8/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_9 XI11_5/net21_6_ xsel_8_ XI11_5/XI0/XI0_8/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_8 XI11_5/net21_7_ xsel_8_ XI11_5/XI0/XI0_8/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_7 XI11_5/net21_8_ xsel_8_ XI11_5/XI0/XI0_8/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_6 XI11_5/net21_9_ xsel_8_ XI11_5/XI0/XI0_8/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_5 XI11_5/net21_10_ xsel_8_ XI11_5/XI0/XI0_8/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_4 XI11_5/net21_11_ xsel_8_ XI11_5/XI0/XI0_8/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_3 XI11_5/net21_12_ xsel_8_ XI11_5/XI0/XI0_8/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_2 XI11_5/net21_13_ xsel_8_ XI11_5/XI0/XI0_8/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_1 XI11_5/net21_14_ xsel_8_ XI11_5/XI0/XI0_8/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_0 XI11_5/net21_15_ xsel_8_ XI11_5/XI0/XI0_8/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_15 XI11_5/XI0/XI0_8/d__15_ xsel_8_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_14 XI11_5/XI0/XI0_8/d__14_ xsel_8_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_13 XI11_5/XI0/XI0_8/d__13_ xsel_8_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_12 XI11_5/XI0/XI0_8/d__12_ xsel_8_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_11 XI11_5/XI0/XI0_8/d__11_ xsel_8_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_10 XI11_5/XI0/XI0_8/d__10_ xsel_8_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_9 XI11_5/XI0/XI0_8/d__9_ xsel_8_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_8 XI11_5/XI0/XI0_8/d__8_ xsel_8_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_7 XI11_5/XI0/XI0_8/d__7_ xsel_8_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_6 XI11_5/XI0/XI0_8/d__6_ xsel_8_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_5 XI11_5/XI0/XI0_8/d__5_ xsel_8_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_4 XI11_5/XI0/XI0_8/d__4_ xsel_8_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_3 XI11_5/XI0/XI0_8/d__3_ xsel_8_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_2 XI11_5/XI0/XI0_8/d__2_ xsel_8_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_1 XI11_5/XI0/XI0_8/d__1_ xsel_8_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_0 XI11_5/XI0/XI0_8/d__0_ xsel_8_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_15 XI11_5/net21_0_ xsel_7_ XI11_5/XI0/XI0_7/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_14 XI11_5/net21_1_ xsel_7_ XI11_5/XI0/XI0_7/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_13 XI11_5/net21_2_ xsel_7_ XI11_5/XI0/XI0_7/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_12 XI11_5/net21_3_ xsel_7_ XI11_5/XI0/XI0_7/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_11 XI11_5/net21_4_ xsel_7_ XI11_5/XI0/XI0_7/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_10 XI11_5/net21_5_ xsel_7_ XI11_5/XI0/XI0_7/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_9 XI11_5/net21_6_ xsel_7_ XI11_5/XI0/XI0_7/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_8 XI11_5/net21_7_ xsel_7_ XI11_5/XI0/XI0_7/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_7 XI11_5/net21_8_ xsel_7_ XI11_5/XI0/XI0_7/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_6 XI11_5/net21_9_ xsel_7_ XI11_5/XI0/XI0_7/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_5 XI11_5/net21_10_ xsel_7_ XI11_5/XI0/XI0_7/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_4 XI11_5/net21_11_ xsel_7_ XI11_5/XI0/XI0_7/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_3 XI11_5/net21_12_ xsel_7_ XI11_5/XI0/XI0_7/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_2 XI11_5/net21_13_ xsel_7_ XI11_5/XI0/XI0_7/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_1 XI11_5/net21_14_ xsel_7_ XI11_5/XI0/XI0_7/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_0 XI11_5/net21_15_ xsel_7_ XI11_5/XI0/XI0_7/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_15 XI11_5/XI0/XI0_7/d__15_ xsel_7_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_14 XI11_5/XI0/XI0_7/d__14_ xsel_7_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_13 XI11_5/XI0/XI0_7/d__13_ xsel_7_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_12 XI11_5/XI0/XI0_7/d__12_ xsel_7_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_11 XI11_5/XI0/XI0_7/d__11_ xsel_7_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_10 XI11_5/XI0/XI0_7/d__10_ xsel_7_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_9 XI11_5/XI0/XI0_7/d__9_ xsel_7_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_8 XI11_5/XI0/XI0_7/d__8_ xsel_7_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_7 XI11_5/XI0/XI0_7/d__7_ xsel_7_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_6 XI11_5/XI0/XI0_7/d__6_ xsel_7_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_5 XI11_5/XI0/XI0_7/d__5_ xsel_7_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_4 XI11_5/XI0/XI0_7/d__4_ xsel_7_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_3 XI11_5/XI0/XI0_7/d__3_ xsel_7_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_2 XI11_5/XI0/XI0_7/d__2_ xsel_7_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_1 XI11_5/XI0/XI0_7/d__1_ xsel_7_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_0 XI11_5/XI0/XI0_7/d__0_ xsel_7_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_15 XI11_5/net21_0_ xsel_6_ XI11_5/XI0/XI0_6/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_14 XI11_5/net21_1_ xsel_6_ XI11_5/XI0/XI0_6/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_13 XI11_5/net21_2_ xsel_6_ XI11_5/XI0/XI0_6/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_12 XI11_5/net21_3_ xsel_6_ XI11_5/XI0/XI0_6/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_11 XI11_5/net21_4_ xsel_6_ XI11_5/XI0/XI0_6/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_10 XI11_5/net21_5_ xsel_6_ XI11_5/XI0/XI0_6/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_9 XI11_5/net21_6_ xsel_6_ XI11_5/XI0/XI0_6/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_8 XI11_5/net21_7_ xsel_6_ XI11_5/XI0/XI0_6/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_7 XI11_5/net21_8_ xsel_6_ XI11_5/XI0/XI0_6/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_6 XI11_5/net21_9_ xsel_6_ XI11_5/XI0/XI0_6/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_5 XI11_5/net21_10_ xsel_6_ XI11_5/XI0/XI0_6/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_4 XI11_5/net21_11_ xsel_6_ XI11_5/XI0/XI0_6/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_3 XI11_5/net21_12_ xsel_6_ XI11_5/XI0/XI0_6/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_2 XI11_5/net21_13_ xsel_6_ XI11_5/XI0/XI0_6/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_1 XI11_5/net21_14_ xsel_6_ XI11_5/XI0/XI0_6/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_0 XI11_5/net21_15_ xsel_6_ XI11_5/XI0/XI0_6/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_15 XI11_5/XI0/XI0_6/d__15_ xsel_6_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_14 XI11_5/XI0/XI0_6/d__14_ xsel_6_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_13 XI11_5/XI0/XI0_6/d__13_ xsel_6_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_12 XI11_5/XI0/XI0_6/d__12_ xsel_6_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_11 XI11_5/XI0/XI0_6/d__11_ xsel_6_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_10 XI11_5/XI0/XI0_6/d__10_ xsel_6_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_9 XI11_5/XI0/XI0_6/d__9_ xsel_6_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_8 XI11_5/XI0/XI0_6/d__8_ xsel_6_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_7 XI11_5/XI0/XI0_6/d__7_ xsel_6_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_6 XI11_5/XI0/XI0_6/d__6_ xsel_6_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_5 XI11_5/XI0/XI0_6/d__5_ xsel_6_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_4 XI11_5/XI0/XI0_6/d__4_ xsel_6_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_3 XI11_5/XI0/XI0_6/d__3_ xsel_6_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_2 XI11_5/XI0/XI0_6/d__2_ xsel_6_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_1 XI11_5/XI0/XI0_6/d__1_ xsel_6_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_0 XI11_5/XI0/XI0_6/d__0_ xsel_6_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_15 XI11_5/net21_0_ xsel_5_ XI11_5/XI0/XI0_5/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_14 XI11_5/net21_1_ xsel_5_ XI11_5/XI0/XI0_5/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_13 XI11_5/net21_2_ xsel_5_ XI11_5/XI0/XI0_5/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_12 XI11_5/net21_3_ xsel_5_ XI11_5/XI0/XI0_5/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_11 XI11_5/net21_4_ xsel_5_ XI11_5/XI0/XI0_5/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_10 XI11_5/net21_5_ xsel_5_ XI11_5/XI0/XI0_5/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_9 XI11_5/net21_6_ xsel_5_ XI11_5/XI0/XI0_5/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_8 XI11_5/net21_7_ xsel_5_ XI11_5/XI0/XI0_5/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_7 XI11_5/net21_8_ xsel_5_ XI11_5/XI0/XI0_5/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_6 XI11_5/net21_9_ xsel_5_ XI11_5/XI0/XI0_5/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_5 XI11_5/net21_10_ xsel_5_ XI11_5/XI0/XI0_5/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_4 XI11_5/net21_11_ xsel_5_ XI11_5/XI0/XI0_5/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_3 XI11_5/net21_12_ xsel_5_ XI11_5/XI0/XI0_5/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_2 XI11_5/net21_13_ xsel_5_ XI11_5/XI0/XI0_5/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_1 XI11_5/net21_14_ xsel_5_ XI11_5/XI0/XI0_5/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_0 XI11_5/net21_15_ xsel_5_ XI11_5/XI0/XI0_5/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_15 XI11_5/XI0/XI0_5/d__15_ xsel_5_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_14 XI11_5/XI0/XI0_5/d__14_ xsel_5_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_13 XI11_5/XI0/XI0_5/d__13_ xsel_5_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_12 XI11_5/XI0/XI0_5/d__12_ xsel_5_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_11 XI11_5/XI0/XI0_5/d__11_ xsel_5_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_10 XI11_5/XI0/XI0_5/d__10_ xsel_5_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_9 XI11_5/XI0/XI0_5/d__9_ xsel_5_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_8 XI11_5/XI0/XI0_5/d__8_ xsel_5_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_7 XI11_5/XI0/XI0_5/d__7_ xsel_5_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_6 XI11_5/XI0/XI0_5/d__6_ xsel_5_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_5 XI11_5/XI0/XI0_5/d__5_ xsel_5_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_4 XI11_5/XI0/XI0_5/d__4_ xsel_5_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_3 XI11_5/XI0/XI0_5/d__3_ xsel_5_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_2 XI11_5/XI0/XI0_5/d__2_ xsel_5_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_1 XI11_5/XI0/XI0_5/d__1_ xsel_5_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_0 XI11_5/XI0/XI0_5/d__0_ xsel_5_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_15 XI11_5/net21_0_ xsel_4_ XI11_5/XI0/XI0_4/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_14 XI11_5/net21_1_ xsel_4_ XI11_5/XI0/XI0_4/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_13 XI11_5/net21_2_ xsel_4_ XI11_5/XI0/XI0_4/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_12 XI11_5/net21_3_ xsel_4_ XI11_5/XI0/XI0_4/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_11 XI11_5/net21_4_ xsel_4_ XI11_5/XI0/XI0_4/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_10 XI11_5/net21_5_ xsel_4_ XI11_5/XI0/XI0_4/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_9 XI11_5/net21_6_ xsel_4_ XI11_5/XI0/XI0_4/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_8 XI11_5/net21_7_ xsel_4_ XI11_5/XI0/XI0_4/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_7 XI11_5/net21_8_ xsel_4_ XI11_5/XI0/XI0_4/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_6 XI11_5/net21_9_ xsel_4_ XI11_5/XI0/XI0_4/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_5 XI11_5/net21_10_ xsel_4_ XI11_5/XI0/XI0_4/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_4 XI11_5/net21_11_ xsel_4_ XI11_5/XI0/XI0_4/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_3 XI11_5/net21_12_ xsel_4_ XI11_5/XI0/XI0_4/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_2 XI11_5/net21_13_ xsel_4_ XI11_5/XI0/XI0_4/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_1 XI11_5/net21_14_ xsel_4_ XI11_5/XI0/XI0_4/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_0 XI11_5/net21_15_ xsel_4_ XI11_5/XI0/XI0_4/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_15 XI11_5/XI0/XI0_4/d__15_ xsel_4_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_14 XI11_5/XI0/XI0_4/d__14_ xsel_4_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_13 XI11_5/XI0/XI0_4/d__13_ xsel_4_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_12 XI11_5/XI0/XI0_4/d__12_ xsel_4_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_11 XI11_5/XI0/XI0_4/d__11_ xsel_4_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_10 XI11_5/XI0/XI0_4/d__10_ xsel_4_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_9 XI11_5/XI0/XI0_4/d__9_ xsel_4_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_8 XI11_5/XI0/XI0_4/d__8_ xsel_4_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_7 XI11_5/XI0/XI0_4/d__7_ xsel_4_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_6 XI11_5/XI0/XI0_4/d__6_ xsel_4_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_5 XI11_5/XI0/XI0_4/d__5_ xsel_4_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_4 XI11_5/XI0/XI0_4/d__4_ xsel_4_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_3 XI11_5/XI0/XI0_4/d__3_ xsel_4_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_2 XI11_5/XI0/XI0_4/d__2_ xsel_4_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_1 XI11_5/XI0/XI0_4/d__1_ xsel_4_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_0 XI11_5/XI0/XI0_4/d__0_ xsel_4_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_15 XI11_5/net21_0_ xsel_3_ XI11_5/XI0/XI0_3/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_14 XI11_5/net21_1_ xsel_3_ XI11_5/XI0/XI0_3/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_13 XI11_5/net21_2_ xsel_3_ XI11_5/XI0/XI0_3/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_12 XI11_5/net21_3_ xsel_3_ XI11_5/XI0/XI0_3/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_11 XI11_5/net21_4_ xsel_3_ XI11_5/XI0/XI0_3/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_10 XI11_5/net21_5_ xsel_3_ XI11_5/XI0/XI0_3/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_9 XI11_5/net21_6_ xsel_3_ XI11_5/XI0/XI0_3/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_8 XI11_5/net21_7_ xsel_3_ XI11_5/XI0/XI0_3/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_7 XI11_5/net21_8_ xsel_3_ XI11_5/XI0/XI0_3/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_6 XI11_5/net21_9_ xsel_3_ XI11_5/XI0/XI0_3/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_5 XI11_5/net21_10_ xsel_3_ XI11_5/XI0/XI0_3/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_4 XI11_5/net21_11_ xsel_3_ XI11_5/XI0/XI0_3/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_3 XI11_5/net21_12_ xsel_3_ XI11_5/XI0/XI0_3/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_2 XI11_5/net21_13_ xsel_3_ XI11_5/XI0/XI0_3/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_1 XI11_5/net21_14_ xsel_3_ XI11_5/XI0/XI0_3/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_0 XI11_5/net21_15_ xsel_3_ XI11_5/XI0/XI0_3/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_15 XI11_5/XI0/XI0_3/d__15_ xsel_3_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_14 XI11_5/XI0/XI0_3/d__14_ xsel_3_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_13 XI11_5/XI0/XI0_3/d__13_ xsel_3_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_12 XI11_5/XI0/XI0_3/d__12_ xsel_3_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_11 XI11_5/XI0/XI0_3/d__11_ xsel_3_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_10 XI11_5/XI0/XI0_3/d__10_ xsel_3_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_9 XI11_5/XI0/XI0_3/d__9_ xsel_3_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_8 XI11_5/XI0/XI0_3/d__8_ xsel_3_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_7 XI11_5/XI0/XI0_3/d__7_ xsel_3_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_6 XI11_5/XI0/XI0_3/d__6_ xsel_3_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_5 XI11_5/XI0/XI0_3/d__5_ xsel_3_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_4 XI11_5/XI0/XI0_3/d__4_ xsel_3_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_3 XI11_5/XI0/XI0_3/d__3_ xsel_3_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_2 XI11_5/XI0/XI0_3/d__2_ xsel_3_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_1 XI11_5/XI0/XI0_3/d__1_ xsel_3_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_0 XI11_5/XI0/XI0_3/d__0_ xsel_3_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_15 XI11_5/net21_0_ xsel_2_ XI11_5/XI0/XI0_2/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_14 XI11_5/net21_1_ xsel_2_ XI11_5/XI0/XI0_2/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_13 XI11_5/net21_2_ xsel_2_ XI11_5/XI0/XI0_2/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_12 XI11_5/net21_3_ xsel_2_ XI11_5/XI0/XI0_2/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_11 XI11_5/net21_4_ xsel_2_ XI11_5/XI0/XI0_2/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_10 XI11_5/net21_5_ xsel_2_ XI11_5/XI0/XI0_2/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_9 XI11_5/net21_6_ xsel_2_ XI11_5/XI0/XI0_2/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_8 XI11_5/net21_7_ xsel_2_ XI11_5/XI0/XI0_2/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_7 XI11_5/net21_8_ xsel_2_ XI11_5/XI0/XI0_2/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_6 XI11_5/net21_9_ xsel_2_ XI11_5/XI0/XI0_2/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_5 XI11_5/net21_10_ xsel_2_ XI11_5/XI0/XI0_2/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_4 XI11_5/net21_11_ xsel_2_ XI11_5/XI0/XI0_2/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_3 XI11_5/net21_12_ xsel_2_ XI11_5/XI0/XI0_2/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_2 XI11_5/net21_13_ xsel_2_ XI11_5/XI0/XI0_2/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_1 XI11_5/net21_14_ xsel_2_ XI11_5/XI0/XI0_2/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_0 XI11_5/net21_15_ xsel_2_ XI11_5/XI0/XI0_2/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_15 XI11_5/XI0/XI0_2/d__15_ xsel_2_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_14 XI11_5/XI0/XI0_2/d__14_ xsel_2_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_13 XI11_5/XI0/XI0_2/d__13_ xsel_2_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_12 XI11_5/XI0/XI0_2/d__12_ xsel_2_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_11 XI11_5/XI0/XI0_2/d__11_ xsel_2_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_10 XI11_5/XI0/XI0_2/d__10_ xsel_2_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_9 XI11_5/XI0/XI0_2/d__9_ xsel_2_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_8 XI11_5/XI0/XI0_2/d__8_ xsel_2_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_7 XI11_5/XI0/XI0_2/d__7_ xsel_2_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_6 XI11_5/XI0/XI0_2/d__6_ xsel_2_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_5 XI11_5/XI0/XI0_2/d__5_ xsel_2_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_4 XI11_5/XI0/XI0_2/d__4_ xsel_2_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_3 XI11_5/XI0/XI0_2/d__3_ xsel_2_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_2 XI11_5/XI0/XI0_2/d__2_ xsel_2_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_1 XI11_5/XI0/XI0_2/d__1_ xsel_2_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_0 XI11_5/XI0/XI0_2/d__0_ xsel_2_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_15 XI11_5/net21_0_ xsel_1_ XI11_5/XI0/XI0_1/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_14 XI11_5/net21_1_ xsel_1_ XI11_5/XI0/XI0_1/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_13 XI11_5/net21_2_ xsel_1_ XI11_5/XI0/XI0_1/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_12 XI11_5/net21_3_ xsel_1_ XI11_5/XI0/XI0_1/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_11 XI11_5/net21_4_ xsel_1_ XI11_5/XI0/XI0_1/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_10 XI11_5/net21_5_ xsel_1_ XI11_5/XI0/XI0_1/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_9 XI11_5/net21_6_ xsel_1_ XI11_5/XI0/XI0_1/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_8 XI11_5/net21_7_ xsel_1_ XI11_5/XI0/XI0_1/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_7 XI11_5/net21_8_ xsel_1_ XI11_5/XI0/XI0_1/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_6 XI11_5/net21_9_ xsel_1_ XI11_5/XI0/XI0_1/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_5 XI11_5/net21_10_ xsel_1_ XI11_5/XI0/XI0_1/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_4 XI11_5/net21_11_ xsel_1_ XI11_5/XI0/XI0_1/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_3 XI11_5/net21_12_ xsel_1_ XI11_5/XI0/XI0_1/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_2 XI11_5/net21_13_ xsel_1_ XI11_5/XI0/XI0_1/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_1 XI11_5/net21_14_ xsel_1_ XI11_5/XI0/XI0_1/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_0 XI11_5/net21_15_ xsel_1_ XI11_5/XI0/XI0_1/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_15 XI11_5/XI0/XI0_1/d__15_ xsel_1_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_14 XI11_5/XI0/XI0_1/d__14_ xsel_1_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_13 XI11_5/XI0/XI0_1/d__13_ xsel_1_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_12 XI11_5/XI0/XI0_1/d__12_ xsel_1_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_11 XI11_5/XI0/XI0_1/d__11_ xsel_1_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_10 XI11_5/XI0/XI0_1/d__10_ xsel_1_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_9 XI11_5/XI0/XI0_1/d__9_ xsel_1_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_8 XI11_5/XI0/XI0_1/d__8_ xsel_1_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_7 XI11_5/XI0/XI0_1/d__7_ xsel_1_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_6 XI11_5/XI0/XI0_1/d__6_ xsel_1_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_5 XI11_5/XI0/XI0_1/d__5_ xsel_1_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_4 XI11_5/XI0/XI0_1/d__4_ xsel_1_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_3 XI11_5/XI0/XI0_1/d__3_ xsel_1_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_2 XI11_5/XI0/XI0_1/d__2_ xsel_1_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_1 XI11_5/XI0/XI0_1/d__1_ xsel_1_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_0 XI11_5/XI0/XI0_1/d__0_ xsel_1_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_15 XI11_5/net21_0_ xsel_0_ XI11_5/XI0/XI0_0/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_14 XI11_5/net21_1_ xsel_0_ XI11_5/XI0/XI0_0/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_13 XI11_5/net21_2_ xsel_0_ XI11_5/XI0/XI0_0/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_12 XI11_5/net21_3_ xsel_0_ XI11_5/XI0/XI0_0/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_11 XI11_5/net21_4_ xsel_0_ XI11_5/XI0/XI0_0/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_10 XI11_5/net21_5_ xsel_0_ XI11_5/XI0/XI0_0/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_9 XI11_5/net21_6_ xsel_0_ XI11_5/XI0/XI0_0/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_8 XI11_5/net21_7_ xsel_0_ XI11_5/XI0/XI0_0/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_7 XI11_5/net21_8_ xsel_0_ XI11_5/XI0/XI0_0/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_6 XI11_5/net21_9_ xsel_0_ XI11_5/XI0/XI0_0/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_5 XI11_5/net21_10_ xsel_0_ XI11_5/XI0/XI0_0/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_4 XI11_5/net21_11_ xsel_0_ XI11_5/XI0/XI0_0/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_3 XI11_5/net21_12_ xsel_0_ XI11_5/XI0/XI0_0/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_2 XI11_5/net21_13_ xsel_0_ XI11_5/XI0/XI0_0/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_1 XI11_5/net21_14_ xsel_0_ XI11_5/XI0/XI0_0/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_0 XI11_5/net21_15_ xsel_0_ XI11_5/XI0/XI0_0/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_15 XI11_5/XI0/XI0_0/d__15_ xsel_0_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_14 XI11_5/XI0/XI0_0/d__14_ xsel_0_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_13 XI11_5/XI0/XI0_0/d__13_ xsel_0_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_12 XI11_5/XI0/XI0_0/d__12_ xsel_0_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_11 XI11_5/XI0/XI0_0/d__11_ xsel_0_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_10 XI11_5/XI0/XI0_0/d__10_ xsel_0_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_9 XI11_5/XI0/XI0_0/d__9_ xsel_0_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_8 XI11_5/XI0/XI0_0/d__8_ xsel_0_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_7 XI11_5/XI0/XI0_0/d__7_ xsel_0_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_6 XI11_5/XI0/XI0_0/d__6_ xsel_0_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_5 XI11_5/XI0/XI0_0/d__5_ xsel_0_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_4 XI11_5/XI0/XI0_0/d__4_ xsel_0_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_3 XI11_5/XI0/XI0_0/d__3_ xsel_0_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_2 XI11_5/XI0/XI0_0/d__2_ xsel_0_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_1 XI11_5/XI0/XI0_0/d__1_ xsel_0_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_0 XI11_5/XI0/XI0_0/d__0_ xsel_0_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI2/MN0_15 XI11_4/net21_0_ ysel_15_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_14 XI11_4/net21_1_ ysel_14_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_13 XI11_4/net21_2_ ysel_13_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_12 XI11_4/net21_3_ ysel_12_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_11 XI11_4/net21_4_ ysel_11_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_10 XI11_4/net21_5_ ysel_10_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_9 XI11_4/net21_6_ ysel_9_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_8 XI11_4/net21_7_ ysel_8_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_7 XI11_4/net21_8_ ysel_7_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_6 XI11_4/net21_9_ ysel_6_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_5 XI11_4/net21_10_ ysel_5_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_4 XI11_4/net21_11_ ysel_4_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_3 XI11_4/net21_12_ ysel_3_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_2 XI11_4/net21_13_ ysel_2_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_1 XI11_4/net21_14_ ysel_1_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_0 XI11_4/net21_15_ ysel_0_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_15 XI11_4/net20_0_ ysel_15_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_14 XI11_4/net20_1_ ysel_14_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_13 XI11_4/net20_2_ ysel_13_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_12 XI11_4/net20_3_ ysel_12_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_11 XI11_4/net20_4_ ysel_11_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_10 XI11_4/net20_5_ ysel_10_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_9 XI11_4/net20_6_ ysel_9_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_8 XI11_4/net20_7_ ysel_8_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_7 XI11_4/net20_8_ ysel_7_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_6 XI11_4/net20_9_ ysel_6_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_5 XI11_4/net20_10_ ysel_5_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_4 XI11_4/net20_11_ ysel_4_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_3 XI11_4/net20_12_ ysel_3_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_2 XI11_4/net20_13_ ysel_2_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_1 XI11_4/net20_14_ ysel_1_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_0 XI11_4/net20_15_ ysel_0_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI4/MN8 vdd XI11_4/XI4/net8 XI11_4/net12 vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_4/XI4/MP0 XI11_4/net9 XI11_4/XI4/net23 vdd vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_4/XI4/MP4 XI11_4/net12 XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI4/MP1 XI11_4/net9 XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI4/MP5 XI11_4/net12 XI11_4/preck XI11_4/net9 vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI4/MN7 vdd XI11_4/XI4/net090 DOUT_4_ vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_4/XI4/MP3 gnd XI11_4/XI4/net089 XI11_4/net12 gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_4/XI4/MN5 XI11_4/net9 XI11_4/XI4/net0103 gnd gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_4/XI4/MN4 XI11_4/XI4/data_out_ XI11_4/XI4/net32 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_4/XI4/MN0 XI11_4/XI4/data_out XI11_4/XI4/net52 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_4/XI4/MN9 gnd XI11_4/XI4/net0112 DOUT_4_ gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_4/XI1_15/MP2 XI11_4/net20_0_ XI11_4/preck XI11_4/net21_0_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_15/MP1 XI11_4/net20_0_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_15/MP0 XI11_4/net21_0_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_14/MP2 XI11_4/net20_1_ XI11_4/preck XI11_4/net21_1_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_14/MP1 XI11_4/net20_1_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_14/MP0 XI11_4/net21_1_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_13/MP2 XI11_4/net20_2_ XI11_4/preck XI11_4/net21_2_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_13/MP1 XI11_4/net20_2_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_13/MP0 XI11_4/net21_2_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_12/MP2 XI11_4/net20_3_ XI11_4/preck XI11_4/net21_3_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_12/MP1 XI11_4/net20_3_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_12/MP0 XI11_4/net21_3_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_11/MP2 XI11_4/net20_4_ XI11_4/preck XI11_4/net21_4_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_11/MP1 XI11_4/net20_4_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_11/MP0 XI11_4/net21_4_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_10/MP2 XI11_4/net20_5_ XI11_4/preck XI11_4/net21_5_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_10/MP1 XI11_4/net20_5_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_10/MP0 XI11_4/net21_5_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_9/MP2 XI11_4/net20_6_ XI11_4/preck XI11_4/net21_6_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_9/MP1 XI11_4/net20_6_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_9/MP0 XI11_4/net21_6_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_8/MP2 XI11_4/net20_7_ XI11_4/preck XI11_4/net21_7_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_8/MP1 XI11_4/net20_7_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_8/MP0 XI11_4/net21_7_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_7/MP2 XI11_4/net20_8_ XI11_4/preck XI11_4/net21_8_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_7/MP1 XI11_4/net20_8_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_7/MP0 XI11_4/net21_8_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_6/MP2 XI11_4/net20_9_ XI11_4/preck XI11_4/net21_9_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_6/MP1 XI11_4/net20_9_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_6/MP0 XI11_4/net21_9_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_5/MP2 XI11_4/net20_10_ XI11_4/preck XI11_4/net21_10_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_5/MP1 XI11_4/net20_10_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_5/MP0 XI11_4/net21_10_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_4/MP2 XI11_4/net20_11_ XI11_4/preck XI11_4/net21_11_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_4/MP1 XI11_4/net20_11_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_4/MP0 XI11_4/net21_11_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_3/MP2 XI11_4/net20_12_ XI11_4/preck XI11_4/net21_12_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_3/MP1 XI11_4/net20_12_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_3/MP0 XI11_4/net21_12_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_2/MP2 XI11_4/net20_13_ XI11_4/preck XI11_4/net21_13_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_2/MP1 XI11_4/net20_13_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_2/MP0 XI11_4/net21_13_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_1/MP2 XI11_4/net20_14_ XI11_4/preck XI11_4/net21_14_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_1/MP1 XI11_4/net20_14_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_1/MP0 XI11_4/net21_14_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_0/MP2 XI11_4/net20_15_ XI11_4/preck XI11_4/net21_15_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_0/MP1 XI11_4/net20_15_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_0/MP0 XI11_4/net21_15_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI0/MN0_15 gnd gnd XI11_4/net21_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_14 gnd gnd XI11_4/net21_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_13 gnd gnd XI11_4/net21_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_12 gnd gnd XI11_4/net21_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_11 gnd gnd XI11_4/net21_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_10 gnd gnd XI11_4/net21_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_9 gnd gnd XI11_4/net21_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_8 gnd gnd XI11_4/net21_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_7 gnd gnd XI11_4/net21_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_6 gnd gnd XI11_4/net21_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_5 gnd gnd XI11_4/net21_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_4 gnd gnd XI11_4/net21_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_3 gnd gnd XI11_4/net21_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_2 gnd gnd XI11_4/net21_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_1 gnd gnd XI11_4/net21_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_0 gnd gnd XI11_4/net21_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_15 gnd gnd XI11_4/net20_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_14 gnd gnd XI11_4/net20_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_13 gnd gnd XI11_4/net20_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_12 gnd gnd XI11_4/net20_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_11 gnd gnd XI11_4/net20_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_10 gnd gnd XI11_4/net20_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_9 gnd gnd XI11_4/net20_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_8 gnd gnd XI11_4/net20_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_7 gnd gnd XI11_4/net20_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_6 gnd gnd XI11_4/net20_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_5 gnd gnd XI11_4/net20_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_4 gnd gnd XI11_4/net20_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_3 gnd gnd XI11_4/net20_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_2 gnd gnd XI11_4/net20_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_1 gnd gnd XI11_4/net20_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_0 gnd gnd XI11_4/net20_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_15 XI11_4/net21_0_ xsel_63_ XI11_4/XI0/XI0_63/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_14 XI11_4/net21_1_ xsel_63_ XI11_4/XI0/XI0_63/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_13 XI11_4/net21_2_ xsel_63_ XI11_4/XI0/XI0_63/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_12 XI11_4/net21_3_ xsel_63_ XI11_4/XI0/XI0_63/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_11 XI11_4/net21_4_ xsel_63_ XI11_4/XI0/XI0_63/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_10 XI11_4/net21_5_ xsel_63_ XI11_4/XI0/XI0_63/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_9 XI11_4/net21_6_ xsel_63_ XI11_4/XI0/XI0_63/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_8 XI11_4/net21_7_ xsel_63_ XI11_4/XI0/XI0_63/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_7 XI11_4/net21_8_ xsel_63_ XI11_4/XI0/XI0_63/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_6 XI11_4/net21_9_ xsel_63_ XI11_4/XI0/XI0_63/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_5 XI11_4/net21_10_ xsel_63_ XI11_4/XI0/XI0_63/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_4 XI11_4/net21_11_ xsel_63_ XI11_4/XI0/XI0_63/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_3 XI11_4/net21_12_ xsel_63_ XI11_4/XI0/XI0_63/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_2 XI11_4/net21_13_ xsel_63_ XI11_4/XI0/XI0_63/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_1 XI11_4/net21_14_ xsel_63_ XI11_4/XI0/XI0_63/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_0 XI11_4/net21_15_ xsel_63_ XI11_4/XI0/XI0_63/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_15 XI11_4/XI0/XI0_63/d__15_ xsel_63_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_14 XI11_4/XI0/XI0_63/d__14_ xsel_63_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_13 XI11_4/XI0/XI0_63/d__13_ xsel_63_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_12 XI11_4/XI0/XI0_63/d__12_ xsel_63_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_11 XI11_4/XI0/XI0_63/d__11_ xsel_63_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_10 XI11_4/XI0/XI0_63/d__10_ xsel_63_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_9 XI11_4/XI0/XI0_63/d__9_ xsel_63_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_8 XI11_4/XI0/XI0_63/d__8_ xsel_63_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_7 XI11_4/XI0/XI0_63/d__7_ xsel_63_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_6 XI11_4/XI0/XI0_63/d__6_ xsel_63_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_5 XI11_4/XI0/XI0_63/d__5_ xsel_63_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_4 XI11_4/XI0/XI0_63/d__4_ xsel_63_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_3 XI11_4/XI0/XI0_63/d__3_ xsel_63_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_2 XI11_4/XI0/XI0_63/d__2_ xsel_63_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_1 XI11_4/XI0/XI0_63/d__1_ xsel_63_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_0 XI11_4/XI0/XI0_63/d__0_ xsel_63_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_15 XI11_4/net21_0_ xsel_62_ XI11_4/XI0/XI0_62/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_14 XI11_4/net21_1_ xsel_62_ XI11_4/XI0/XI0_62/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_13 XI11_4/net21_2_ xsel_62_ XI11_4/XI0/XI0_62/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_12 XI11_4/net21_3_ xsel_62_ XI11_4/XI0/XI0_62/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_11 XI11_4/net21_4_ xsel_62_ XI11_4/XI0/XI0_62/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_10 XI11_4/net21_5_ xsel_62_ XI11_4/XI0/XI0_62/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_9 XI11_4/net21_6_ xsel_62_ XI11_4/XI0/XI0_62/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_8 XI11_4/net21_7_ xsel_62_ XI11_4/XI0/XI0_62/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_7 XI11_4/net21_8_ xsel_62_ XI11_4/XI0/XI0_62/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_6 XI11_4/net21_9_ xsel_62_ XI11_4/XI0/XI0_62/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_5 XI11_4/net21_10_ xsel_62_ XI11_4/XI0/XI0_62/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_4 XI11_4/net21_11_ xsel_62_ XI11_4/XI0/XI0_62/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_3 XI11_4/net21_12_ xsel_62_ XI11_4/XI0/XI0_62/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_2 XI11_4/net21_13_ xsel_62_ XI11_4/XI0/XI0_62/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_1 XI11_4/net21_14_ xsel_62_ XI11_4/XI0/XI0_62/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_0 XI11_4/net21_15_ xsel_62_ XI11_4/XI0/XI0_62/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_15 XI11_4/XI0/XI0_62/d__15_ xsel_62_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_14 XI11_4/XI0/XI0_62/d__14_ xsel_62_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_13 XI11_4/XI0/XI0_62/d__13_ xsel_62_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_12 XI11_4/XI0/XI0_62/d__12_ xsel_62_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_11 XI11_4/XI0/XI0_62/d__11_ xsel_62_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_10 XI11_4/XI0/XI0_62/d__10_ xsel_62_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_9 XI11_4/XI0/XI0_62/d__9_ xsel_62_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_8 XI11_4/XI0/XI0_62/d__8_ xsel_62_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_7 XI11_4/XI0/XI0_62/d__7_ xsel_62_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_6 XI11_4/XI0/XI0_62/d__6_ xsel_62_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_5 XI11_4/XI0/XI0_62/d__5_ xsel_62_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_4 XI11_4/XI0/XI0_62/d__4_ xsel_62_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_3 XI11_4/XI0/XI0_62/d__3_ xsel_62_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_2 XI11_4/XI0/XI0_62/d__2_ xsel_62_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_1 XI11_4/XI0/XI0_62/d__1_ xsel_62_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_0 XI11_4/XI0/XI0_62/d__0_ xsel_62_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_15 XI11_4/net21_0_ xsel_61_ XI11_4/XI0/XI0_61/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_14 XI11_4/net21_1_ xsel_61_ XI11_4/XI0/XI0_61/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_13 XI11_4/net21_2_ xsel_61_ XI11_4/XI0/XI0_61/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_12 XI11_4/net21_3_ xsel_61_ XI11_4/XI0/XI0_61/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_11 XI11_4/net21_4_ xsel_61_ XI11_4/XI0/XI0_61/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_10 XI11_4/net21_5_ xsel_61_ XI11_4/XI0/XI0_61/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_9 XI11_4/net21_6_ xsel_61_ XI11_4/XI0/XI0_61/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_8 XI11_4/net21_7_ xsel_61_ XI11_4/XI0/XI0_61/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_7 XI11_4/net21_8_ xsel_61_ XI11_4/XI0/XI0_61/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_6 XI11_4/net21_9_ xsel_61_ XI11_4/XI0/XI0_61/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_5 XI11_4/net21_10_ xsel_61_ XI11_4/XI0/XI0_61/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_4 XI11_4/net21_11_ xsel_61_ XI11_4/XI0/XI0_61/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_3 XI11_4/net21_12_ xsel_61_ XI11_4/XI0/XI0_61/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_2 XI11_4/net21_13_ xsel_61_ XI11_4/XI0/XI0_61/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_1 XI11_4/net21_14_ xsel_61_ XI11_4/XI0/XI0_61/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_0 XI11_4/net21_15_ xsel_61_ XI11_4/XI0/XI0_61/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_15 XI11_4/XI0/XI0_61/d__15_ xsel_61_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_14 XI11_4/XI0/XI0_61/d__14_ xsel_61_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_13 XI11_4/XI0/XI0_61/d__13_ xsel_61_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_12 XI11_4/XI0/XI0_61/d__12_ xsel_61_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_11 XI11_4/XI0/XI0_61/d__11_ xsel_61_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_10 XI11_4/XI0/XI0_61/d__10_ xsel_61_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_9 XI11_4/XI0/XI0_61/d__9_ xsel_61_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_8 XI11_4/XI0/XI0_61/d__8_ xsel_61_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_7 XI11_4/XI0/XI0_61/d__7_ xsel_61_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_6 XI11_4/XI0/XI0_61/d__6_ xsel_61_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_5 XI11_4/XI0/XI0_61/d__5_ xsel_61_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_4 XI11_4/XI0/XI0_61/d__4_ xsel_61_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_3 XI11_4/XI0/XI0_61/d__3_ xsel_61_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_2 XI11_4/XI0/XI0_61/d__2_ xsel_61_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_1 XI11_4/XI0/XI0_61/d__1_ xsel_61_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_0 XI11_4/XI0/XI0_61/d__0_ xsel_61_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_15 XI11_4/net21_0_ xsel_60_ XI11_4/XI0/XI0_60/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_14 XI11_4/net21_1_ xsel_60_ XI11_4/XI0/XI0_60/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_13 XI11_4/net21_2_ xsel_60_ XI11_4/XI0/XI0_60/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_12 XI11_4/net21_3_ xsel_60_ XI11_4/XI0/XI0_60/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_11 XI11_4/net21_4_ xsel_60_ XI11_4/XI0/XI0_60/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_10 XI11_4/net21_5_ xsel_60_ XI11_4/XI0/XI0_60/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_9 XI11_4/net21_6_ xsel_60_ XI11_4/XI0/XI0_60/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_8 XI11_4/net21_7_ xsel_60_ XI11_4/XI0/XI0_60/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_7 XI11_4/net21_8_ xsel_60_ XI11_4/XI0/XI0_60/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_6 XI11_4/net21_9_ xsel_60_ XI11_4/XI0/XI0_60/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_5 XI11_4/net21_10_ xsel_60_ XI11_4/XI0/XI0_60/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_4 XI11_4/net21_11_ xsel_60_ XI11_4/XI0/XI0_60/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_3 XI11_4/net21_12_ xsel_60_ XI11_4/XI0/XI0_60/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_2 XI11_4/net21_13_ xsel_60_ XI11_4/XI0/XI0_60/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_1 XI11_4/net21_14_ xsel_60_ XI11_4/XI0/XI0_60/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_0 XI11_4/net21_15_ xsel_60_ XI11_4/XI0/XI0_60/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_15 XI11_4/XI0/XI0_60/d__15_ xsel_60_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_14 XI11_4/XI0/XI0_60/d__14_ xsel_60_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_13 XI11_4/XI0/XI0_60/d__13_ xsel_60_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_12 XI11_4/XI0/XI0_60/d__12_ xsel_60_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_11 XI11_4/XI0/XI0_60/d__11_ xsel_60_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_10 XI11_4/XI0/XI0_60/d__10_ xsel_60_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_9 XI11_4/XI0/XI0_60/d__9_ xsel_60_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_8 XI11_4/XI0/XI0_60/d__8_ xsel_60_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_7 XI11_4/XI0/XI0_60/d__7_ xsel_60_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_6 XI11_4/XI0/XI0_60/d__6_ xsel_60_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_5 XI11_4/XI0/XI0_60/d__5_ xsel_60_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_4 XI11_4/XI0/XI0_60/d__4_ xsel_60_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_3 XI11_4/XI0/XI0_60/d__3_ xsel_60_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_2 XI11_4/XI0/XI0_60/d__2_ xsel_60_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_1 XI11_4/XI0/XI0_60/d__1_ xsel_60_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_0 XI11_4/XI0/XI0_60/d__0_ xsel_60_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_15 XI11_4/net21_0_ xsel_59_ XI11_4/XI0/XI0_59/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_14 XI11_4/net21_1_ xsel_59_ XI11_4/XI0/XI0_59/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_13 XI11_4/net21_2_ xsel_59_ XI11_4/XI0/XI0_59/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_12 XI11_4/net21_3_ xsel_59_ XI11_4/XI0/XI0_59/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_11 XI11_4/net21_4_ xsel_59_ XI11_4/XI0/XI0_59/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_10 XI11_4/net21_5_ xsel_59_ XI11_4/XI0/XI0_59/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_9 XI11_4/net21_6_ xsel_59_ XI11_4/XI0/XI0_59/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_8 XI11_4/net21_7_ xsel_59_ XI11_4/XI0/XI0_59/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_7 XI11_4/net21_8_ xsel_59_ XI11_4/XI0/XI0_59/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_6 XI11_4/net21_9_ xsel_59_ XI11_4/XI0/XI0_59/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_5 XI11_4/net21_10_ xsel_59_ XI11_4/XI0/XI0_59/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_4 XI11_4/net21_11_ xsel_59_ XI11_4/XI0/XI0_59/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_3 XI11_4/net21_12_ xsel_59_ XI11_4/XI0/XI0_59/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_2 XI11_4/net21_13_ xsel_59_ XI11_4/XI0/XI0_59/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_1 XI11_4/net21_14_ xsel_59_ XI11_4/XI0/XI0_59/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_0 XI11_4/net21_15_ xsel_59_ XI11_4/XI0/XI0_59/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_15 XI11_4/XI0/XI0_59/d__15_ xsel_59_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_14 XI11_4/XI0/XI0_59/d__14_ xsel_59_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_13 XI11_4/XI0/XI0_59/d__13_ xsel_59_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_12 XI11_4/XI0/XI0_59/d__12_ xsel_59_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_11 XI11_4/XI0/XI0_59/d__11_ xsel_59_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_10 XI11_4/XI0/XI0_59/d__10_ xsel_59_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_9 XI11_4/XI0/XI0_59/d__9_ xsel_59_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_8 XI11_4/XI0/XI0_59/d__8_ xsel_59_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_7 XI11_4/XI0/XI0_59/d__7_ xsel_59_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_6 XI11_4/XI0/XI0_59/d__6_ xsel_59_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_5 XI11_4/XI0/XI0_59/d__5_ xsel_59_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_4 XI11_4/XI0/XI0_59/d__4_ xsel_59_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_3 XI11_4/XI0/XI0_59/d__3_ xsel_59_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_2 XI11_4/XI0/XI0_59/d__2_ xsel_59_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_1 XI11_4/XI0/XI0_59/d__1_ xsel_59_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_0 XI11_4/XI0/XI0_59/d__0_ xsel_59_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_15 XI11_4/net21_0_ xsel_58_ XI11_4/XI0/XI0_58/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_14 XI11_4/net21_1_ xsel_58_ XI11_4/XI0/XI0_58/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_13 XI11_4/net21_2_ xsel_58_ XI11_4/XI0/XI0_58/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_12 XI11_4/net21_3_ xsel_58_ XI11_4/XI0/XI0_58/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_11 XI11_4/net21_4_ xsel_58_ XI11_4/XI0/XI0_58/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_10 XI11_4/net21_5_ xsel_58_ XI11_4/XI0/XI0_58/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_9 XI11_4/net21_6_ xsel_58_ XI11_4/XI0/XI0_58/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_8 XI11_4/net21_7_ xsel_58_ XI11_4/XI0/XI0_58/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_7 XI11_4/net21_8_ xsel_58_ XI11_4/XI0/XI0_58/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_6 XI11_4/net21_9_ xsel_58_ XI11_4/XI0/XI0_58/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_5 XI11_4/net21_10_ xsel_58_ XI11_4/XI0/XI0_58/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_4 XI11_4/net21_11_ xsel_58_ XI11_4/XI0/XI0_58/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_3 XI11_4/net21_12_ xsel_58_ XI11_4/XI0/XI0_58/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_2 XI11_4/net21_13_ xsel_58_ XI11_4/XI0/XI0_58/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_1 XI11_4/net21_14_ xsel_58_ XI11_4/XI0/XI0_58/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_0 XI11_4/net21_15_ xsel_58_ XI11_4/XI0/XI0_58/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_15 XI11_4/XI0/XI0_58/d__15_ xsel_58_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_14 XI11_4/XI0/XI0_58/d__14_ xsel_58_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_13 XI11_4/XI0/XI0_58/d__13_ xsel_58_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_12 XI11_4/XI0/XI0_58/d__12_ xsel_58_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_11 XI11_4/XI0/XI0_58/d__11_ xsel_58_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_10 XI11_4/XI0/XI0_58/d__10_ xsel_58_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_9 XI11_4/XI0/XI0_58/d__9_ xsel_58_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_8 XI11_4/XI0/XI0_58/d__8_ xsel_58_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_7 XI11_4/XI0/XI0_58/d__7_ xsel_58_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_6 XI11_4/XI0/XI0_58/d__6_ xsel_58_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_5 XI11_4/XI0/XI0_58/d__5_ xsel_58_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_4 XI11_4/XI0/XI0_58/d__4_ xsel_58_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_3 XI11_4/XI0/XI0_58/d__3_ xsel_58_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_2 XI11_4/XI0/XI0_58/d__2_ xsel_58_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_1 XI11_4/XI0/XI0_58/d__1_ xsel_58_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_0 XI11_4/XI0/XI0_58/d__0_ xsel_58_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_15 XI11_4/net21_0_ xsel_57_ XI11_4/XI0/XI0_57/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_14 XI11_4/net21_1_ xsel_57_ XI11_4/XI0/XI0_57/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_13 XI11_4/net21_2_ xsel_57_ XI11_4/XI0/XI0_57/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_12 XI11_4/net21_3_ xsel_57_ XI11_4/XI0/XI0_57/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_11 XI11_4/net21_4_ xsel_57_ XI11_4/XI0/XI0_57/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_10 XI11_4/net21_5_ xsel_57_ XI11_4/XI0/XI0_57/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_9 XI11_4/net21_6_ xsel_57_ XI11_4/XI0/XI0_57/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_8 XI11_4/net21_7_ xsel_57_ XI11_4/XI0/XI0_57/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_7 XI11_4/net21_8_ xsel_57_ XI11_4/XI0/XI0_57/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_6 XI11_4/net21_9_ xsel_57_ XI11_4/XI0/XI0_57/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_5 XI11_4/net21_10_ xsel_57_ XI11_4/XI0/XI0_57/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_4 XI11_4/net21_11_ xsel_57_ XI11_4/XI0/XI0_57/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_3 XI11_4/net21_12_ xsel_57_ XI11_4/XI0/XI0_57/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_2 XI11_4/net21_13_ xsel_57_ XI11_4/XI0/XI0_57/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_1 XI11_4/net21_14_ xsel_57_ XI11_4/XI0/XI0_57/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_0 XI11_4/net21_15_ xsel_57_ XI11_4/XI0/XI0_57/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_15 XI11_4/XI0/XI0_57/d__15_ xsel_57_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_14 XI11_4/XI0/XI0_57/d__14_ xsel_57_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_13 XI11_4/XI0/XI0_57/d__13_ xsel_57_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_12 XI11_4/XI0/XI0_57/d__12_ xsel_57_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_11 XI11_4/XI0/XI0_57/d__11_ xsel_57_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_10 XI11_4/XI0/XI0_57/d__10_ xsel_57_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_9 XI11_4/XI0/XI0_57/d__9_ xsel_57_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_8 XI11_4/XI0/XI0_57/d__8_ xsel_57_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_7 XI11_4/XI0/XI0_57/d__7_ xsel_57_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_6 XI11_4/XI0/XI0_57/d__6_ xsel_57_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_5 XI11_4/XI0/XI0_57/d__5_ xsel_57_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_4 XI11_4/XI0/XI0_57/d__4_ xsel_57_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_3 XI11_4/XI0/XI0_57/d__3_ xsel_57_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_2 XI11_4/XI0/XI0_57/d__2_ xsel_57_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_1 XI11_4/XI0/XI0_57/d__1_ xsel_57_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_0 XI11_4/XI0/XI0_57/d__0_ xsel_57_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_15 XI11_4/net21_0_ xsel_56_ XI11_4/XI0/XI0_56/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_14 XI11_4/net21_1_ xsel_56_ XI11_4/XI0/XI0_56/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_13 XI11_4/net21_2_ xsel_56_ XI11_4/XI0/XI0_56/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_12 XI11_4/net21_3_ xsel_56_ XI11_4/XI0/XI0_56/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_11 XI11_4/net21_4_ xsel_56_ XI11_4/XI0/XI0_56/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_10 XI11_4/net21_5_ xsel_56_ XI11_4/XI0/XI0_56/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_9 XI11_4/net21_6_ xsel_56_ XI11_4/XI0/XI0_56/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_8 XI11_4/net21_7_ xsel_56_ XI11_4/XI0/XI0_56/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_7 XI11_4/net21_8_ xsel_56_ XI11_4/XI0/XI0_56/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_6 XI11_4/net21_9_ xsel_56_ XI11_4/XI0/XI0_56/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_5 XI11_4/net21_10_ xsel_56_ XI11_4/XI0/XI0_56/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_4 XI11_4/net21_11_ xsel_56_ XI11_4/XI0/XI0_56/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_3 XI11_4/net21_12_ xsel_56_ XI11_4/XI0/XI0_56/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_2 XI11_4/net21_13_ xsel_56_ XI11_4/XI0/XI0_56/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_1 XI11_4/net21_14_ xsel_56_ XI11_4/XI0/XI0_56/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_0 XI11_4/net21_15_ xsel_56_ XI11_4/XI0/XI0_56/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_15 XI11_4/XI0/XI0_56/d__15_ xsel_56_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_14 XI11_4/XI0/XI0_56/d__14_ xsel_56_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_13 XI11_4/XI0/XI0_56/d__13_ xsel_56_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_12 XI11_4/XI0/XI0_56/d__12_ xsel_56_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_11 XI11_4/XI0/XI0_56/d__11_ xsel_56_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_10 XI11_4/XI0/XI0_56/d__10_ xsel_56_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_9 XI11_4/XI0/XI0_56/d__9_ xsel_56_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_8 XI11_4/XI0/XI0_56/d__8_ xsel_56_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_7 XI11_4/XI0/XI0_56/d__7_ xsel_56_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_6 XI11_4/XI0/XI0_56/d__6_ xsel_56_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_5 XI11_4/XI0/XI0_56/d__5_ xsel_56_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_4 XI11_4/XI0/XI0_56/d__4_ xsel_56_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_3 XI11_4/XI0/XI0_56/d__3_ xsel_56_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_2 XI11_4/XI0/XI0_56/d__2_ xsel_56_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_1 XI11_4/XI0/XI0_56/d__1_ xsel_56_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_0 XI11_4/XI0/XI0_56/d__0_ xsel_56_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_15 XI11_4/net21_0_ xsel_55_ XI11_4/XI0/XI0_55/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_14 XI11_4/net21_1_ xsel_55_ XI11_4/XI0/XI0_55/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_13 XI11_4/net21_2_ xsel_55_ XI11_4/XI0/XI0_55/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_12 XI11_4/net21_3_ xsel_55_ XI11_4/XI0/XI0_55/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_11 XI11_4/net21_4_ xsel_55_ XI11_4/XI0/XI0_55/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_10 XI11_4/net21_5_ xsel_55_ XI11_4/XI0/XI0_55/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_9 XI11_4/net21_6_ xsel_55_ XI11_4/XI0/XI0_55/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_8 XI11_4/net21_7_ xsel_55_ XI11_4/XI0/XI0_55/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_7 XI11_4/net21_8_ xsel_55_ XI11_4/XI0/XI0_55/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_6 XI11_4/net21_9_ xsel_55_ XI11_4/XI0/XI0_55/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_5 XI11_4/net21_10_ xsel_55_ XI11_4/XI0/XI0_55/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_4 XI11_4/net21_11_ xsel_55_ XI11_4/XI0/XI0_55/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_3 XI11_4/net21_12_ xsel_55_ XI11_4/XI0/XI0_55/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_2 XI11_4/net21_13_ xsel_55_ XI11_4/XI0/XI0_55/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_1 XI11_4/net21_14_ xsel_55_ XI11_4/XI0/XI0_55/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_0 XI11_4/net21_15_ xsel_55_ XI11_4/XI0/XI0_55/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_15 XI11_4/XI0/XI0_55/d__15_ xsel_55_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_14 XI11_4/XI0/XI0_55/d__14_ xsel_55_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_13 XI11_4/XI0/XI0_55/d__13_ xsel_55_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_12 XI11_4/XI0/XI0_55/d__12_ xsel_55_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_11 XI11_4/XI0/XI0_55/d__11_ xsel_55_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_10 XI11_4/XI0/XI0_55/d__10_ xsel_55_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_9 XI11_4/XI0/XI0_55/d__9_ xsel_55_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_8 XI11_4/XI0/XI0_55/d__8_ xsel_55_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_7 XI11_4/XI0/XI0_55/d__7_ xsel_55_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_6 XI11_4/XI0/XI0_55/d__6_ xsel_55_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_5 XI11_4/XI0/XI0_55/d__5_ xsel_55_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_4 XI11_4/XI0/XI0_55/d__4_ xsel_55_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_3 XI11_4/XI0/XI0_55/d__3_ xsel_55_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_2 XI11_4/XI0/XI0_55/d__2_ xsel_55_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_1 XI11_4/XI0/XI0_55/d__1_ xsel_55_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_0 XI11_4/XI0/XI0_55/d__0_ xsel_55_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_15 XI11_4/net21_0_ xsel_54_ XI11_4/XI0/XI0_54/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_14 XI11_4/net21_1_ xsel_54_ XI11_4/XI0/XI0_54/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_13 XI11_4/net21_2_ xsel_54_ XI11_4/XI0/XI0_54/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_12 XI11_4/net21_3_ xsel_54_ XI11_4/XI0/XI0_54/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_11 XI11_4/net21_4_ xsel_54_ XI11_4/XI0/XI0_54/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_10 XI11_4/net21_5_ xsel_54_ XI11_4/XI0/XI0_54/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_9 XI11_4/net21_6_ xsel_54_ XI11_4/XI0/XI0_54/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_8 XI11_4/net21_7_ xsel_54_ XI11_4/XI0/XI0_54/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_7 XI11_4/net21_8_ xsel_54_ XI11_4/XI0/XI0_54/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_6 XI11_4/net21_9_ xsel_54_ XI11_4/XI0/XI0_54/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_5 XI11_4/net21_10_ xsel_54_ XI11_4/XI0/XI0_54/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_4 XI11_4/net21_11_ xsel_54_ XI11_4/XI0/XI0_54/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_3 XI11_4/net21_12_ xsel_54_ XI11_4/XI0/XI0_54/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_2 XI11_4/net21_13_ xsel_54_ XI11_4/XI0/XI0_54/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_1 XI11_4/net21_14_ xsel_54_ XI11_4/XI0/XI0_54/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_0 XI11_4/net21_15_ xsel_54_ XI11_4/XI0/XI0_54/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_15 XI11_4/XI0/XI0_54/d__15_ xsel_54_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_14 XI11_4/XI0/XI0_54/d__14_ xsel_54_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_13 XI11_4/XI0/XI0_54/d__13_ xsel_54_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_12 XI11_4/XI0/XI0_54/d__12_ xsel_54_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_11 XI11_4/XI0/XI0_54/d__11_ xsel_54_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_10 XI11_4/XI0/XI0_54/d__10_ xsel_54_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_9 XI11_4/XI0/XI0_54/d__9_ xsel_54_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_8 XI11_4/XI0/XI0_54/d__8_ xsel_54_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_7 XI11_4/XI0/XI0_54/d__7_ xsel_54_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_6 XI11_4/XI0/XI0_54/d__6_ xsel_54_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_5 XI11_4/XI0/XI0_54/d__5_ xsel_54_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_4 XI11_4/XI0/XI0_54/d__4_ xsel_54_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_3 XI11_4/XI0/XI0_54/d__3_ xsel_54_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_2 XI11_4/XI0/XI0_54/d__2_ xsel_54_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_1 XI11_4/XI0/XI0_54/d__1_ xsel_54_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_0 XI11_4/XI0/XI0_54/d__0_ xsel_54_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_15 XI11_4/net21_0_ xsel_53_ XI11_4/XI0/XI0_53/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_14 XI11_4/net21_1_ xsel_53_ XI11_4/XI0/XI0_53/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_13 XI11_4/net21_2_ xsel_53_ XI11_4/XI0/XI0_53/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_12 XI11_4/net21_3_ xsel_53_ XI11_4/XI0/XI0_53/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_11 XI11_4/net21_4_ xsel_53_ XI11_4/XI0/XI0_53/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_10 XI11_4/net21_5_ xsel_53_ XI11_4/XI0/XI0_53/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_9 XI11_4/net21_6_ xsel_53_ XI11_4/XI0/XI0_53/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_8 XI11_4/net21_7_ xsel_53_ XI11_4/XI0/XI0_53/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_7 XI11_4/net21_8_ xsel_53_ XI11_4/XI0/XI0_53/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_6 XI11_4/net21_9_ xsel_53_ XI11_4/XI0/XI0_53/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_5 XI11_4/net21_10_ xsel_53_ XI11_4/XI0/XI0_53/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_4 XI11_4/net21_11_ xsel_53_ XI11_4/XI0/XI0_53/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_3 XI11_4/net21_12_ xsel_53_ XI11_4/XI0/XI0_53/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_2 XI11_4/net21_13_ xsel_53_ XI11_4/XI0/XI0_53/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_1 XI11_4/net21_14_ xsel_53_ XI11_4/XI0/XI0_53/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_0 XI11_4/net21_15_ xsel_53_ XI11_4/XI0/XI0_53/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_15 XI11_4/XI0/XI0_53/d__15_ xsel_53_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_14 XI11_4/XI0/XI0_53/d__14_ xsel_53_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_13 XI11_4/XI0/XI0_53/d__13_ xsel_53_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_12 XI11_4/XI0/XI0_53/d__12_ xsel_53_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_11 XI11_4/XI0/XI0_53/d__11_ xsel_53_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_10 XI11_4/XI0/XI0_53/d__10_ xsel_53_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_9 XI11_4/XI0/XI0_53/d__9_ xsel_53_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_8 XI11_4/XI0/XI0_53/d__8_ xsel_53_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_7 XI11_4/XI0/XI0_53/d__7_ xsel_53_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_6 XI11_4/XI0/XI0_53/d__6_ xsel_53_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_5 XI11_4/XI0/XI0_53/d__5_ xsel_53_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_4 XI11_4/XI0/XI0_53/d__4_ xsel_53_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_3 XI11_4/XI0/XI0_53/d__3_ xsel_53_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_2 XI11_4/XI0/XI0_53/d__2_ xsel_53_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_1 XI11_4/XI0/XI0_53/d__1_ xsel_53_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_0 XI11_4/XI0/XI0_53/d__0_ xsel_53_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_15 XI11_4/net21_0_ xsel_52_ XI11_4/XI0/XI0_52/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_14 XI11_4/net21_1_ xsel_52_ XI11_4/XI0/XI0_52/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_13 XI11_4/net21_2_ xsel_52_ XI11_4/XI0/XI0_52/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_12 XI11_4/net21_3_ xsel_52_ XI11_4/XI0/XI0_52/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_11 XI11_4/net21_4_ xsel_52_ XI11_4/XI0/XI0_52/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_10 XI11_4/net21_5_ xsel_52_ XI11_4/XI0/XI0_52/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_9 XI11_4/net21_6_ xsel_52_ XI11_4/XI0/XI0_52/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_8 XI11_4/net21_7_ xsel_52_ XI11_4/XI0/XI0_52/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_7 XI11_4/net21_8_ xsel_52_ XI11_4/XI0/XI0_52/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_6 XI11_4/net21_9_ xsel_52_ XI11_4/XI0/XI0_52/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_5 XI11_4/net21_10_ xsel_52_ XI11_4/XI0/XI0_52/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_4 XI11_4/net21_11_ xsel_52_ XI11_4/XI0/XI0_52/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_3 XI11_4/net21_12_ xsel_52_ XI11_4/XI0/XI0_52/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_2 XI11_4/net21_13_ xsel_52_ XI11_4/XI0/XI0_52/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_1 XI11_4/net21_14_ xsel_52_ XI11_4/XI0/XI0_52/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_0 XI11_4/net21_15_ xsel_52_ XI11_4/XI0/XI0_52/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_15 XI11_4/XI0/XI0_52/d__15_ xsel_52_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_14 XI11_4/XI0/XI0_52/d__14_ xsel_52_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_13 XI11_4/XI0/XI0_52/d__13_ xsel_52_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_12 XI11_4/XI0/XI0_52/d__12_ xsel_52_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_11 XI11_4/XI0/XI0_52/d__11_ xsel_52_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_10 XI11_4/XI0/XI0_52/d__10_ xsel_52_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_9 XI11_4/XI0/XI0_52/d__9_ xsel_52_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_8 XI11_4/XI0/XI0_52/d__8_ xsel_52_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_7 XI11_4/XI0/XI0_52/d__7_ xsel_52_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_6 XI11_4/XI0/XI0_52/d__6_ xsel_52_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_5 XI11_4/XI0/XI0_52/d__5_ xsel_52_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_4 XI11_4/XI0/XI0_52/d__4_ xsel_52_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_3 XI11_4/XI0/XI0_52/d__3_ xsel_52_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_2 XI11_4/XI0/XI0_52/d__2_ xsel_52_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_1 XI11_4/XI0/XI0_52/d__1_ xsel_52_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_0 XI11_4/XI0/XI0_52/d__0_ xsel_52_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_15 XI11_4/net21_0_ xsel_51_ XI11_4/XI0/XI0_51/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_14 XI11_4/net21_1_ xsel_51_ XI11_4/XI0/XI0_51/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_13 XI11_4/net21_2_ xsel_51_ XI11_4/XI0/XI0_51/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_12 XI11_4/net21_3_ xsel_51_ XI11_4/XI0/XI0_51/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_11 XI11_4/net21_4_ xsel_51_ XI11_4/XI0/XI0_51/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_10 XI11_4/net21_5_ xsel_51_ XI11_4/XI0/XI0_51/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_9 XI11_4/net21_6_ xsel_51_ XI11_4/XI0/XI0_51/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_8 XI11_4/net21_7_ xsel_51_ XI11_4/XI0/XI0_51/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_7 XI11_4/net21_8_ xsel_51_ XI11_4/XI0/XI0_51/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_6 XI11_4/net21_9_ xsel_51_ XI11_4/XI0/XI0_51/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_5 XI11_4/net21_10_ xsel_51_ XI11_4/XI0/XI0_51/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_4 XI11_4/net21_11_ xsel_51_ XI11_4/XI0/XI0_51/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_3 XI11_4/net21_12_ xsel_51_ XI11_4/XI0/XI0_51/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_2 XI11_4/net21_13_ xsel_51_ XI11_4/XI0/XI0_51/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_1 XI11_4/net21_14_ xsel_51_ XI11_4/XI0/XI0_51/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_0 XI11_4/net21_15_ xsel_51_ XI11_4/XI0/XI0_51/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_15 XI11_4/XI0/XI0_51/d__15_ xsel_51_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_14 XI11_4/XI0/XI0_51/d__14_ xsel_51_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_13 XI11_4/XI0/XI0_51/d__13_ xsel_51_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_12 XI11_4/XI0/XI0_51/d__12_ xsel_51_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_11 XI11_4/XI0/XI0_51/d__11_ xsel_51_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_10 XI11_4/XI0/XI0_51/d__10_ xsel_51_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_9 XI11_4/XI0/XI0_51/d__9_ xsel_51_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_8 XI11_4/XI0/XI0_51/d__8_ xsel_51_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_7 XI11_4/XI0/XI0_51/d__7_ xsel_51_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_6 XI11_4/XI0/XI0_51/d__6_ xsel_51_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_5 XI11_4/XI0/XI0_51/d__5_ xsel_51_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_4 XI11_4/XI0/XI0_51/d__4_ xsel_51_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_3 XI11_4/XI0/XI0_51/d__3_ xsel_51_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_2 XI11_4/XI0/XI0_51/d__2_ xsel_51_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_1 XI11_4/XI0/XI0_51/d__1_ xsel_51_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_0 XI11_4/XI0/XI0_51/d__0_ xsel_51_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_15 XI11_4/net21_0_ xsel_50_ XI11_4/XI0/XI0_50/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_14 XI11_4/net21_1_ xsel_50_ XI11_4/XI0/XI0_50/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_13 XI11_4/net21_2_ xsel_50_ XI11_4/XI0/XI0_50/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_12 XI11_4/net21_3_ xsel_50_ XI11_4/XI0/XI0_50/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_11 XI11_4/net21_4_ xsel_50_ XI11_4/XI0/XI0_50/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_10 XI11_4/net21_5_ xsel_50_ XI11_4/XI0/XI0_50/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_9 XI11_4/net21_6_ xsel_50_ XI11_4/XI0/XI0_50/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_8 XI11_4/net21_7_ xsel_50_ XI11_4/XI0/XI0_50/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_7 XI11_4/net21_8_ xsel_50_ XI11_4/XI0/XI0_50/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_6 XI11_4/net21_9_ xsel_50_ XI11_4/XI0/XI0_50/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_5 XI11_4/net21_10_ xsel_50_ XI11_4/XI0/XI0_50/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_4 XI11_4/net21_11_ xsel_50_ XI11_4/XI0/XI0_50/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_3 XI11_4/net21_12_ xsel_50_ XI11_4/XI0/XI0_50/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_2 XI11_4/net21_13_ xsel_50_ XI11_4/XI0/XI0_50/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_1 XI11_4/net21_14_ xsel_50_ XI11_4/XI0/XI0_50/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_0 XI11_4/net21_15_ xsel_50_ XI11_4/XI0/XI0_50/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_15 XI11_4/XI0/XI0_50/d__15_ xsel_50_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_14 XI11_4/XI0/XI0_50/d__14_ xsel_50_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_13 XI11_4/XI0/XI0_50/d__13_ xsel_50_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_12 XI11_4/XI0/XI0_50/d__12_ xsel_50_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_11 XI11_4/XI0/XI0_50/d__11_ xsel_50_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_10 XI11_4/XI0/XI0_50/d__10_ xsel_50_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_9 XI11_4/XI0/XI0_50/d__9_ xsel_50_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_8 XI11_4/XI0/XI0_50/d__8_ xsel_50_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_7 XI11_4/XI0/XI0_50/d__7_ xsel_50_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_6 XI11_4/XI0/XI0_50/d__6_ xsel_50_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_5 XI11_4/XI0/XI0_50/d__5_ xsel_50_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_4 XI11_4/XI0/XI0_50/d__4_ xsel_50_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_3 XI11_4/XI0/XI0_50/d__3_ xsel_50_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_2 XI11_4/XI0/XI0_50/d__2_ xsel_50_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_1 XI11_4/XI0/XI0_50/d__1_ xsel_50_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_0 XI11_4/XI0/XI0_50/d__0_ xsel_50_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_15 XI11_4/net21_0_ xsel_49_ XI11_4/XI0/XI0_49/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_14 XI11_4/net21_1_ xsel_49_ XI11_4/XI0/XI0_49/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_13 XI11_4/net21_2_ xsel_49_ XI11_4/XI0/XI0_49/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_12 XI11_4/net21_3_ xsel_49_ XI11_4/XI0/XI0_49/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_11 XI11_4/net21_4_ xsel_49_ XI11_4/XI0/XI0_49/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_10 XI11_4/net21_5_ xsel_49_ XI11_4/XI0/XI0_49/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_9 XI11_4/net21_6_ xsel_49_ XI11_4/XI0/XI0_49/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_8 XI11_4/net21_7_ xsel_49_ XI11_4/XI0/XI0_49/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_7 XI11_4/net21_8_ xsel_49_ XI11_4/XI0/XI0_49/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_6 XI11_4/net21_9_ xsel_49_ XI11_4/XI0/XI0_49/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_5 XI11_4/net21_10_ xsel_49_ XI11_4/XI0/XI0_49/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_4 XI11_4/net21_11_ xsel_49_ XI11_4/XI0/XI0_49/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_3 XI11_4/net21_12_ xsel_49_ XI11_4/XI0/XI0_49/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_2 XI11_4/net21_13_ xsel_49_ XI11_4/XI0/XI0_49/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_1 XI11_4/net21_14_ xsel_49_ XI11_4/XI0/XI0_49/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_0 XI11_4/net21_15_ xsel_49_ XI11_4/XI0/XI0_49/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_15 XI11_4/XI0/XI0_49/d__15_ xsel_49_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_14 XI11_4/XI0/XI0_49/d__14_ xsel_49_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_13 XI11_4/XI0/XI0_49/d__13_ xsel_49_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_12 XI11_4/XI0/XI0_49/d__12_ xsel_49_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_11 XI11_4/XI0/XI0_49/d__11_ xsel_49_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_10 XI11_4/XI0/XI0_49/d__10_ xsel_49_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_9 XI11_4/XI0/XI0_49/d__9_ xsel_49_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_8 XI11_4/XI0/XI0_49/d__8_ xsel_49_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_7 XI11_4/XI0/XI0_49/d__7_ xsel_49_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_6 XI11_4/XI0/XI0_49/d__6_ xsel_49_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_5 XI11_4/XI0/XI0_49/d__5_ xsel_49_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_4 XI11_4/XI0/XI0_49/d__4_ xsel_49_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_3 XI11_4/XI0/XI0_49/d__3_ xsel_49_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_2 XI11_4/XI0/XI0_49/d__2_ xsel_49_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_1 XI11_4/XI0/XI0_49/d__1_ xsel_49_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_0 XI11_4/XI0/XI0_49/d__0_ xsel_49_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_15 XI11_4/net21_0_ xsel_48_ XI11_4/XI0/XI0_48/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_14 XI11_4/net21_1_ xsel_48_ XI11_4/XI0/XI0_48/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_13 XI11_4/net21_2_ xsel_48_ XI11_4/XI0/XI0_48/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_12 XI11_4/net21_3_ xsel_48_ XI11_4/XI0/XI0_48/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_11 XI11_4/net21_4_ xsel_48_ XI11_4/XI0/XI0_48/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_10 XI11_4/net21_5_ xsel_48_ XI11_4/XI0/XI0_48/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_9 XI11_4/net21_6_ xsel_48_ XI11_4/XI0/XI0_48/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_8 XI11_4/net21_7_ xsel_48_ XI11_4/XI0/XI0_48/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_7 XI11_4/net21_8_ xsel_48_ XI11_4/XI0/XI0_48/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_6 XI11_4/net21_9_ xsel_48_ XI11_4/XI0/XI0_48/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_5 XI11_4/net21_10_ xsel_48_ XI11_4/XI0/XI0_48/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_4 XI11_4/net21_11_ xsel_48_ XI11_4/XI0/XI0_48/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_3 XI11_4/net21_12_ xsel_48_ XI11_4/XI0/XI0_48/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_2 XI11_4/net21_13_ xsel_48_ XI11_4/XI0/XI0_48/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_1 XI11_4/net21_14_ xsel_48_ XI11_4/XI0/XI0_48/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_0 XI11_4/net21_15_ xsel_48_ XI11_4/XI0/XI0_48/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_15 XI11_4/XI0/XI0_48/d__15_ xsel_48_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_14 XI11_4/XI0/XI0_48/d__14_ xsel_48_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_13 XI11_4/XI0/XI0_48/d__13_ xsel_48_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_12 XI11_4/XI0/XI0_48/d__12_ xsel_48_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_11 XI11_4/XI0/XI0_48/d__11_ xsel_48_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_10 XI11_4/XI0/XI0_48/d__10_ xsel_48_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_9 XI11_4/XI0/XI0_48/d__9_ xsel_48_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_8 XI11_4/XI0/XI0_48/d__8_ xsel_48_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_7 XI11_4/XI0/XI0_48/d__7_ xsel_48_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_6 XI11_4/XI0/XI0_48/d__6_ xsel_48_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_5 XI11_4/XI0/XI0_48/d__5_ xsel_48_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_4 XI11_4/XI0/XI0_48/d__4_ xsel_48_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_3 XI11_4/XI0/XI0_48/d__3_ xsel_48_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_2 XI11_4/XI0/XI0_48/d__2_ xsel_48_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_1 XI11_4/XI0/XI0_48/d__1_ xsel_48_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_0 XI11_4/XI0/XI0_48/d__0_ xsel_48_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_15 XI11_4/net21_0_ xsel_47_ XI11_4/XI0/XI0_47/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_14 XI11_4/net21_1_ xsel_47_ XI11_4/XI0/XI0_47/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_13 XI11_4/net21_2_ xsel_47_ XI11_4/XI0/XI0_47/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_12 XI11_4/net21_3_ xsel_47_ XI11_4/XI0/XI0_47/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_11 XI11_4/net21_4_ xsel_47_ XI11_4/XI0/XI0_47/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_10 XI11_4/net21_5_ xsel_47_ XI11_4/XI0/XI0_47/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_9 XI11_4/net21_6_ xsel_47_ XI11_4/XI0/XI0_47/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_8 XI11_4/net21_7_ xsel_47_ XI11_4/XI0/XI0_47/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_7 XI11_4/net21_8_ xsel_47_ XI11_4/XI0/XI0_47/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_6 XI11_4/net21_9_ xsel_47_ XI11_4/XI0/XI0_47/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_5 XI11_4/net21_10_ xsel_47_ XI11_4/XI0/XI0_47/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_4 XI11_4/net21_11_ xsel_47_ XI11_4/XI0/XI0_47/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_3 XI11_4/net21_12_ xsel_47_ XI11_4/XI0/XI0_47/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_2 XI11_4/net21_13_ xsel_47_ XI11_4/XI0/XI0_47/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_1 XI11_4/net21_14_ xsel_47_ XI11_4/XI0/XI0_47/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_0 XI11_4/net21_15_ xsel_47_ XI11_4/XI0/XI0_47/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_15 XI11_4/XI0/XI0_47/d__15_ xsel_47_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_14 XI11_4/XI0/XI0_47/d__14_ xsel_47_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_13 XI11_4/XI0/XI0_47/d__13_ xsel_47_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_12 XI11_4/XI0/XI0_47/d__12_ xsel_47_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_11 XI11_4/XI0/XI0_47/d__11_ xsel_47_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_10 XI11_4/XI0/XI0_47/d__10_ xsel_47_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_9 XI11_4/XI0/XI0_47/d__9_ xsel_47_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_8 XI11_4/XI0/XI0_47/d__8_ xsel_47_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_7 XI11_4/XI0/XI0_47/d__7_ xsel_47_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_6 XI11_4/XI0/XI0_47/d__6_ xsel_47_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_5 XI11_4/XI0/XI0_47/d__5_ xsel_47_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_4 XI11_4/XI0/XI0_47/d__4_ xsel_47_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_3 XI11_4/XI0/XI0_47/d__3_ xsel_47_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_2 XI11_4/XI0/XI0_47/d__2_ xsel_47_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_1 XI11_4/XI0/XI0_47/d__1_ xsel_47_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_0 XI11_4/XI0/XI0_47/d__0_ xsel_47_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_15 XI11_4/net21_0_ xsel_46_ XI11_4/XI0/XI0_46/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_14 XI11_4/net21_1_ xsel_46_ XI11_4/XI0/XI0_46/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_13 XI11_4/net21_2_ xsel_46_ XI11_4/XI0/XI0_46/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_12 XI11_4/net21_3_ xsel_46_ XI11_4/XI0/XI0_46/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_11 XI11_4/net21_4_ xsel_46_ XI11_4/XI0/XI0_46/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_10 XI11_4/net21_5_ xsel_46_ XI11_4/XI0/XI0_46/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_9 XI11_4/net21_6_ xsel_46_ XI11_4/XI0/XI0_46/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_8 XI11_4/net21_7_ xsel_46_ XI11_4/XI0/XI0_46/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_7 XI11_4/net21_8_ xsel_46_ XI11_4/XI0/XI0_46/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_6 XI11_4/net21_9_ xsel_46_ XI11_4/XI0/XI0_46/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_5 XI11_4/net21_10_ xsel_46_ XI11_4/XI0/XI0_46/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_4 XI11_4/net21_11_ xsel_46_ XI11_4/XI0/XI0_46/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_3 XI11_4/net21_12_ xsel_46_ XI11_4/XI0/XI0_46/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_2 XI11_4/net21_13_ xsel_46_ XI11_4/XI0/XI0_46/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_1 XI11_4/net21_14_ xsel_46_ XI11_4/XI0/XI0_46/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_0 XI11_4/net21_15_ xsel_46_ XI11_4/XI0/XI0_46/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_15 XI11_4/XI0/XI0_46/d__15_ xsel_46_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_14 XI11_4/XI0/XI0_46/d__14_ xsel_46_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_13 XI11_4/XI0/XI0_46/d__13_ xsel_46_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_12 XI11_4/XI0/XI0_46/d__12_ xsel_46_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_11 XI11_4/XI0/XI0_46/d__11_ xsel_46_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_10 XI11_4/XI0/XI0_46/d__10_ xsel_46_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_9 XI11_4/XI0/XI0_46/d__9_ xsel_46_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_8 XI11_4/XI0/XI0_46/d__8_ xsel_46_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_7 XI11_4/XI0/XI0_46/d__7_ xsel_46_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_6 XI11_4/XI0/XI0_46/d__6_ xsel_46_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_5 XI11_4/XI0/XI0_46/d__5_ xsel_46_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_4 XI11_4/XI0/XI0_46/d__4_ xsel_46_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_3 XI11_4/XI0/XI0_46/d__3_ xsel_46_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_2 XI11_4/XI0/XI0_46/d__2_ xsel_46_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_1 XI11_4/XI0/XI0_46/d__1_ xsel_46_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_0 XI11_4/XI0/XI0_46/d__0_ xsel_46_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_15 XI11_4/net21_0_ xsel_45_ XI11_4/XI0/XI0_45/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_14 XI11_4/net21_1_ xsel_45_ XI11_4/XI0/XI0_45/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_13 XI11_4/net21_2_ xsel_45_ XI11_4/XI0/XI0_45/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_12 XI11_4/net21_3_ xsel_45_ XI11_4/XI0/XI0_45/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_11 XI11_4/net21_4_ xsel_45_ XI11_4/XI0/XI0_45/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_10 XI11_4/net21_5_ xsel_45_ XI11_4/XI0/XI0_45/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_9 XI11_4/net21_6_ xsel_45_ XI11_4/XI0/XI0_45/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_8 XI11_4/net21_7_ xsel_45_ XI11_4/XI0/XI0_45/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_7 XI11_4/net21_8_ xsel_45_ XI11_4/XI0/XI0_45/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_6 XI11_4/net21_9_ xsel_45_ XI11_4/XI0/XI0_45/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_5 XI11_4/net21_10_ xsel_45_ XI11_4/XI0/XI0_45/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_4 XI11_4/net21_11_ xsel_45_ XI11_4/XI0/XI0_45/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_3 XI11_4/net21_12_ xsel_45_ XI11_4/XI0/XI0_45/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_2 XI11_4/net21_13_ xsel_45_ XI11_4/XI0/XI0_45/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_1 XI11_4/net21_14_ xsel_45_ XI11_4/XI0/XI0_45/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_0 XI11_4/net21_15_ xsel_45_ XI11_4/XI0/XI0_45/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_15 XI11_4/XI0/XI0_45/d__15_ xsel_45_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_14 XI11_4/XI0/XI0_45/d__14_ xsel_45_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_13 XI11_4/XI0/XI0_45/d__13_ xsel_45_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_12 XI11_4/XI0/XI0_45/d__12_ xsel_45_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_11 XI11_4/XI0/XI0_45/d__11_ xsel_45_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_10 XI11_4/XI0/XI0_45/d__10_ xsel_45_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_9 XI11_4/XI0/XI0_45/d__9_ xsel_45_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_8 XI11_4/XI0/XI0_45/d__8_ xsel_45_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_7 XI11_4/XI0/XI0_45/d__7_ xsel_45_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_6 XI11_4/XI0/XI0_45/d__6_ xsel_45_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_5 XI11_4/XI0/XI0_45/d__5_ xsel_45_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_4 XI11_4/XI0/XI0_45/d__4_ xsel_45_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_3 XI11_4/XI0/XI0_45/d__3_ xsel_45_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_2 XI11_4/XI0/XI0_45/d__2_ xsel_45_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_1 XI11_4/XI0/XI0_45/d__1_ xsel_45_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_0 XI11_4/XI0/XI0_45/d__0_ xsel_45_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_15 XI11_4/net21_0_ xsel_44_ XI11_4/XI0/XI0_44/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_14 XI11_4/net21_1_ xsel_44_ XI11_4/XI0/XI0_44/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_13 XI11_4/net21_2_ xsel_44_ XI11_4/XI0/XI0_44/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_12 XI11_4/net21_3_ xsel_44_ XI11_4/XI0/XI0_44/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_11 XI11_4/net21_4_ xsel_44_ XI11_4/XI0/XI0_44/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_10 XI11_4/net21_5_ xsel_44_ XI11_4/XI0/XI0_44/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_9 XI11_4/net21_6_ xsel_44_ XI11_4/XI0/XI0_44/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_8 XI11_4/net21_7_ xsel_44_ XI11_4/XI0/XI0_44/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_7 XI11_4/net21_8_ xsel_44_ XI11_4/XI0/XI0_44/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_6 XI11_4/net21_9_ xsel_44_ XI11_4/XI0/XI0_44/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_5 XI11_4/net21_10_ xsel_44_ XI11_4/XI0/XI0_44/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_4 XI11_4/net21_11_ xsel_44_ XI11_4/XI0/XI0_44/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_3 XI11_4/net21_12_ xsel_44_ XI11_4/XI0/XI0_44/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_2 XI11_4/net21_13_ xsel_44_ XI11_4/XI0/XI0_44/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_1 XI11_4/net21_14_ xsel_44_ XI11_4/XI0/XI0_44/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_0 XI11_4/net21_15_ xsel_44_ XI11_4/XI0/XI0_44/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_15 XI11_4/XI0/XI0_44/d__15_ xsel_44_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_14 XI11_4/XI0/XI0_44/d__14_ xsel_44_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_13 XI11_4/XI0/XI0_44/d__13_ xsel_44_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_12 XI11_4/XI0/XI0_44/d__12_ xsel_44_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_11 XI11_4/XI0/XI0_44/d__11_ xsel_44_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_10 XI11_4/XI0/XI0_44/d__10_ xsel_44_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_9 XI11_4/XI0/XI0_44/d__9_ xsel_44_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_8 XI11_4/XI0/XI0_44/d__8_ xsel_44_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_7 XI11_4/XI0/XI0_44/d__7_ xsel_44_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_6 XI11_4/XI0/XI0_44/d__6_ xsel_44_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_5 XI11_4/XI0/XI0_44/d__5_ xsel_44_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_4 XI11_4/XI0/XI0_44/d__4_ xsel_44_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_3 XI11_4/XI0/XI0_44/d__3_ xsel_44_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_2 XI11_4/XI0/XI0_44/d__2_ xsel_44_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_1 XI11_4/XI0/XI0_44/d__1_ xsel_44_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_0 XI11_4/XI0/XI0_44/d__0_ xsel_44_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_15 XI11_4/net21_0_ xsel_43_ XI11_4/XI0/XI0_43/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_14 XI11_4/net21_1_ xsel_43_ XI11_4/XI0/XI0_43/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_13 XI11_4/net21_2_ xsel_43_ XI11_4/XI0/XI0_43/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_12 XI11_4/net21_3_ xsel_43_ XI11_4/XI0/XI0_43/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_11 XI11_4/net21_4_ xsel_43_ XI11_4/XI0/XI0_43/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_10 XI11_4/net21_5_ xsel_43_ XI11_4/XI0/XI0_43/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_9 XI11_4/net21_6_ xsel_43_ XI11_4/XI0/XI0_43/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_8 XI11_4/net21_7_ xsel_43_ XI11_4/XI0/XI0_43/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_7 XI11_4/net21_8_ xsel_43_ XI11_4/XI0/XI0_43/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_6 XI11_4/net21_9_ xsel_43_ XI11_4/XI0/XI0_43/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_5 XI11_4/net21_10_ xsel_43_ XI11_4/XI0/XI0_43/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_4 XI11_4/net21_11_ xsel_43_ XI11_4/XI0/XI0_43/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_3 XI11_4/net21_12_ xsel_43_ XI11_4/XI0/XI0_43/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_2 XI11_4/net21_13_ xsel_43_ XI11_4/XI0/XI0_43/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_1 XI11_4/net21_14_ xsel_43_ XI11_4/XI0/XI0_43/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_0 XI11_4/net21_15_ xsel_43_ XI11_4/XI0/XI0_43/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_15 XI11_4/XI0/XI0_43/d__15_ xsel_43_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_14 XI11_4/XI0/XI0_43/d__14_ xsel_43_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_13 XI11_4/XI0/XI0_43/d__13_ xsel_43_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_12 XI11_4/XI0/XI0_43/d__12_ xsel_43_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_11 XI11_4/XI0/XI0_43/d__11_ xsel_43_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_10 XI11_4/XI0/XI0_43/d__10_ xsel_43_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_9 XI11_4/XI0/XI0_43/d__9_ xsel_43_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_8 XI11_4/XI0/XI0_43/d__8_ xsel_43_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_7 XI11_4/XI0/XI0_43/d__7_ xsel_43_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_6 XI11_4/XI0/XI0_43/d__6_ xsel_43_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_5 XI11_4/XI0/XI0_43/d__5_ xsel_43_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_4 XI11_4/XI0/XI0_43/d__4_ xsel_43_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_3 XI11_4/XI0/XI0_43/d__3_ xsel_43_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_2 XI11_4/XI0/XI0_43/d__2_ xsel_43_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_1 XI11_4/XI0/XI0_43/d__1_ xsel_43_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_0 XI11_4/XI0/XI0_43/d__0_ xsel_43_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_15 XI11_4/net21_0_ xsel_42_ XI11_4/XI0/XI0_42/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_14 XI11_4/net21_1_ xsel_42_ XI11_4/XI0/XI0_42/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_13 XI11_4/net21_2_ xsel_42_ XI11_4/XI0/XI0_42/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_12 XI11_4/net21_3_ xsel_42_ XI11_4/XI0/XI0_42/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_11 XI11_4/net21_4_ xsel_42_ XI11_4/XI0/XI0_42/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_10 XI11_4/net21_5_ xsel_42_ XI11_4/XI0/XI0_42/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_9 XI11_4/net21_6_ xsel_42_ XI11_4/XI0/XI0_42/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_8 XI11_4/net21_7_ xsel_42_ XI11_4/XI0/XI0_42/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_7 XI11_4/net21_8_ xsel_42_ XI11_4/XI0/XI0_42/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_6 XI11_4/net21_9_ xsel_42_ XI11_4/XI0/XI0_42/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_5 XI11_4/net21_10_ xsel_42_ XI11_4/XI0/XI0_42/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_4 XI11_4/net21_11_ xsel_42_ XI11_4/XI0/XI0_42/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_3 XI11_4/net21_12_ xsel_42_ XI11_4/XI0/XI0_42/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_2 XI11_4/net21_13_ xsel_42_ XI11_4/XI0/XI0_42/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_1 XI11_4/net21_14_ xsel_42_ XI11_4/XI0/XI0_42/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_0 XI11_4/net21_15_ xsel_42_ XI11_4/XI0/XI0_42/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_15 XI11_4/XI0/XI0_42/d__15_ xsel_42_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_14 XI11_4/XI0/XI0_42/d__14_ xsel_42_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_13 XI11_4/XI0/XI0_42/d__13_ xsel_42_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_12 XI11_4/XI0/XI0_42/d__12_ xsel_42_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_11 XI11_4/XI0/XI0_42/d__11_ xsel_42_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_10 XI11_4/XI0/XI0_42/d__10_ xsel_42_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_9 XI11_4/XI0/XI0_42/d__9_ xsel_42_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_8 XI11_4/XI0/XI0_42/d__8_ xsel_42_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_7 XI11_4/XI0/XI0_42/d__7_ xsel_42_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_6 XI11_4/XI0/XI0_42/d__6_ xsel_42_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_5 XI11_4/XI0/XI0_42/d__5_ xsel_42_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_4 XI11_4/XI0/XI0_42/d__4_ xsel_42_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_3 XI11_4/XI0/XI0_42/d__3_ xsel_42_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_2 XI11_4/XI0/XI0_42/d__2_ xsel_42_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_1 XI11_4/XI0/XI0_42/d__1_ xsel_42_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_0 XI11_4/XI0/XI0_42/d__0_ xsel_42_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_15 XI11_4/net21_0_ xsel_41_ XI11_4/XI0/XI0_41/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_14 XI11_4/net21_1_ xsel_41_ XI11_4/XI0/XI0_41/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_13 XI11_4/net21_2_ xsel_41_ XI11_4/XI0/XI0_41/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_12 XI11_4/net21_3_ xsel_41_ XI11_4/XI0/XI0_41/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_11 XI11_4/net21_4_ xsel_41_ XI11_4/XI0/XI0_41/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_10 XI11_4/net21_5_ xsel_41_ XI11_4/XI0/XI0_41/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_9 XI11_4/net21_6_ xsel_41_ XI11_4/XI0/XI0_41/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_8 XI11_4/net21_7_ xsel_41_ XI11_4/XI0/XI0_41/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_7 XI11_4/net21_8_ xsel_41_ XI11_4/XI0/XI0_41/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_6 XI11_4/net21_9_ xsel_41_ XI11_4/XI0/XI0_41/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_5 XI11_4/net21_10_ xsel_41_ XI11_4/XI0/XI0_41/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_4 XI11_4/net21_11_ xsel_41_ XI11_4/XI0/XI0_41/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_3 XI11_4/net21_12_ xsel_41_ XI11_4/XI0/XI0_41/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_2 XI11_4/net21_13_ xsel_41_ XI11_4/XI0/XI0_41/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_1 XI11_4/net21_14_ xsel_41_ XI11_4/XI0/XI0_41/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_0 XI11_4/net21_15_ xsel_41_ XI11_4/XI0/XI0_41/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_15 XI11_4/XI0/XI0_41/d__15_ xsel_41_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_14 XI11_4/XI0/XI0_41/d__14_ xsel_41_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_13 XI11_4/XI0/XI0_41/d__13_ xsel_41_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_12 XI11_4/XI0/XI0_41/d__12_ xsel_41_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_11 XI11_4/XI0/XI0_41/d__11_ xsel_41_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_10 XI11_4/XI0/XI0_41/d__10_ xsel_41_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_9 XI11_4/XI0/XI0_41/d__9_ xsel_41_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_8 XI11_4/XI0/XI0_41/d__8_ xsel_41_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_7 XI11_4/XI0/XI0_41/d__7_ xsel_41_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_6 XI11_4/XI0/XI0_41/d__6_ xsel_41_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_5 XI11_4/XI0/XI0_41/d__5_ xsel_41_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_4 XI11_4/XI0/XI0_41/d__4_ xsel_41_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_3 XI11_4/XI0/XI0_41/d__3_ xsel_41_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_2 XI11_4/XI0/XI0_41/d__2_ xsel_41_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_1 XI11_4/XI0/XI0_41/d__1_ xsel_41_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_0 XI11_4/XI0/XI0_41/d__0_ xsel_41_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_15 XI11_4/net21_0_ xsel_40_ XI11_4/XI0/XI0_40/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_14 XI11_4/net21_1_ xsel_40_ XI11_4/XI0/XI0_40/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_13 XI11_4/net21_2_ xsel_40_ XI11_4/XI0/XI0_40/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_12 XI11_4/net21_3_ xsel_40_ XI11_4/XI0/XI0_40/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_11 XI11_4/net21_4_ xsel_40_ XI11_4/XI0/XI0_40/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_10 XI11_4/net21_5_ xsel_40_ XI11_4/XI0/XI0_40/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_9 XI11_4/net21_6_ xsel_40_ XI11_4/XI0/XI0_40/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_8 XI11_4/net21_7_ xsel_40_ XI11_4/XI0/XI0_40/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_7 XI11_4/net21_8_ xsel_40_ XI11_4/XI0/XI0_40/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_6 XI11_4/net21_9_ xsel_40_ XI11_4/XI0/XI0_40/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_5 XI11_4/net21_10_ xsel_40_ XI11_4/XI0/XI0_40/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_4 XI11_4/net21_11_ xsel_40_ XI11_4/XI0/XI0_40/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_3 XI11_4/net21_12_ xsel_40_ XI11_4/XI0/XI0_40/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_2 XI11_4/net21_13_ xsel_40_ XI11_4/XI0/XI0_40/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_1 XI11_4/net21_14_ xsel_40_ XI11_4/XI0/XI0_40/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_0 XI11_4/net21_15_ xsel_40_ XI11_4/XI0/XI0_40/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_15 XI11_4/XI0/XI0_40/d__15_ xsel_40_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_14 XI11_4/XI0/XI0_40/d__14_ xsel_40_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_13 XI11_4/XI0/XI0_40/d__13_ xsel_40_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_12 XI11_4/XI0/XI0_40/d__12_ xsel_40_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_11 XI11_4/XI0/XI0_40/d__11_ xsel_40_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_10 XI11_4/XI0/XI0_40/d__10_ xsel_40_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_9 XI11_4/XI0/XI0_40/d__9_ xsel_40_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_8 XI11_4/XI0/XI0_40/d__8_ xsel_40_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_7 XI11_4/XI0/XI0_40/d__7_ xsel_40_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_6 XI11_4/XI0/XI0_40/d__6_ xsel_40_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_5 XI11_4/XI0/XI0_40/d__5_ xsel_40_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_4 XI11_4/XI0/XI0_40/d__4_ xsel_40_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_3 XI11_4/XI0/XI0_40/d__3_ xsel_40_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_2 XI11_4/XI0/XI0_40/d__2_ xsel_40_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_1 XI11_4/XI0/XI0_40/d__1_ xsel_40_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_0 XI11_4/XI0/XI0_40/d__0_ xsel_40_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_15 XI11_4/net21_0_ xsel_39_ XI11_4/XI0/XI0_39/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_14 XI11_4/net21_1_ xsel_39_ XI11_4/XI0/XI0_39/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_13 XI11_4/net21_2_ xsel_39_ XI11_4/XI0/XI0_39/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_12 XI11_4/net21_3_ xsel_39_ XI11_4/XI0/XI0_39/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_11 XI11_4/net21_4_ xsel_39_ XI11_4/XI0/XI0_39/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_10 XI11_4/net21_5_ xsel_39_ XI11_4/XI0/XI0_39/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_9 XI11_4/net21_6_ xsel_39_ XI11_4/XI0/XI0_39/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_8 XI11_4/net21_7_ xsel_39_ XI11_4/XI0/XI0_39/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_7 XI11_4/net21_8_ xsel_39_ XI11_4/XI0/XI0_39/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_6 XI11_4/net21_9_ xsel_39_ XI11_4/XI0/XI0_39/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_5 XI11_4/net21_10_ xsel_39_ XI11_4/XI0/XI0_39/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_4 XI11_4/net21_11_ xsel_39_ XI11_4/XI0/XI0_39/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_3 XI11_4/net21_12_ xsel_39_ XI11_4/XI0/XI0_39/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_2 XI11_4/net21_13_ xsel_39_ XI11_4/XI0/XI0_39/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_1 XI11_4/net21_14_ xsel_39_ XI11_4/XI0/XI0_39/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_0 XI11_4/net21_15_ xsel_39_ XI11_4/XI0/XI0_39/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_15 XI11_4/XI0/XI0_39/d__15_ xsel_39_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_14 XI11_4/XI0/XI0_39/d__14_ xsel_39_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_13 XI11_4/XI0/XI0_39/d__13_ xsel_39_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_12 XI11_4/XI0/XI0_39/d__12_ xsel_39_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_11 XI11_4/XI0/XI0_39/d__11_ xsel_39_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_10 XI11_4/XI0/XI0_39/d__10_ xsel_39_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_9 XI11_4/XI0/XI0_39/d__9_ xsel_39_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_8 XI11_4/XI0/XI0_39/d__8_ xsel_39_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_7 XI11_4/XI0/XI0_39/d__7_ xsel_39_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_6 XI11_4/XI0/XI0_39/d__6_ xsel_39_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_5 XI11_4/XI0/XI0_39/d__5_ xsel_39_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_4 XI11_4/XI0/XI0_39/d__4_ xsel_39_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_3 XI11_4/XI0/XI0_39/d__3_ xsel_39_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_2 XI11_4/XI0/XI0_39/d__2_ xsel_39_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_1 XI11_4/XI0/XI0_39/d__1_ xsel_39_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_0 XI11_4/XI0/XI0_39/d__0_ xsel_39_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_15 XI11_4/net21_0_ xsel_38_ XI11_4/XI0/XI0_38/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_14 XI11_4/net21_1_ xsel_38_ XI11_4/XI0/XI0_38/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_13 XI11_4/net21_2_ xsel_38_ XI11_4/XI0/XI0_38/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_12 XI11_4/net21_3_ xsel_38_ XI11_4/XI0/XI0_38/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_11 XI11_4/net21_4_ xsel_38_ XI11_4/XI0/XI0_38/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_10 XI11_4/net21_5_ xsel_38_ XI11_4/XI0/XI0_38/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_9 XI11_4/net21_6_ xsel_38_ XI11_4/XI0/XI0_38/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_8 XI11_4/net21_7_ xsel_38_ XI11_4/XI0/XI0_38/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_7 XI11_4/net21_8_ xsel_38_ XI11_4/XI0/XI0_38/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_6 XI11_4/net21_9_ xsel_38_ XI11_4/XI0/XI0_38/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_5 XI11_4/net21_10_ xsel_38_ XI11_4/XI0/XI0_38/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_4 XI11_4/net21_11_ xsel_38_ XI11_4/XI0/XI0_38/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_3 XI11_4/net21_12_ xsel_38_ XI11_4/XI0/XI0_38/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_2 XI11_4/net21_13_ xsel_38_ XI11_4/XI0/XI0_38/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_1 XI11_4/net21_14_ xsel_38_ XI11_4/XI0/XI0_38/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_0 XI11_4/net21_15_ xsel_38_ XI11_4/XI0/XI0_38/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_15 XI11_4/XI0/XI0_38/d__15_ xsel_38_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_14 XI11_4/XI0/XI0_38/d__14_ xsel_38_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_13 XI11_4/XI0/XI0_38/d__13_ xsel_38_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_12 XI11_4/XI0/XI0_38/d__12_ xsel_38_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_11 XI11_4/XI0/XI0_38/d__11_ xsel_38_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_10 XI11_4/XI0/XI0_38/d__10_ xsel_38_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_9 XI11_4/XI0/XI0_38/d__9_ xsel_38_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_8 XI11_4/XI0/XI0_38/d__8_ xsel_38_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_7 XI11_4/XI0/XI0_38/d__7_ xsel_38_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_6 XI11_4/XI0/XI0_38/d__6_ xsel_38_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_5 XI11_4/XI0/XI0_38/d__5_ xsel_38_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_4 XI11_4/XI0/XI0_38/d__4_ xsel_38_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_3 XI11_4/XI0/XI0_38/d__3_ xsel_38_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_2 XI11_4/XI0/XI0_38/d__2_ xsel_38_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_1 XI11_4/XI0/XI0_38/d__1_ xsel_38_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_0 XI11_4/XI0/XI0_38/d__0_ xsel_38_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_15 XI11_4/net21_0_ xsel_37_ XI11_4/XI0/XI0_37/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_14 XI11_4/net21_1_ xsel_37_ XI11_4/XI0/XI0_37/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_13 XI11_4/net21_2_ xsel_37_ XI11_4/XI0/XI0_37/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_12 XI11_4/net21_3_ xsel_37_ XI11_4/XI0/XI0_37/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_11 XI11_4/net21_4_ xsel_37_ XI11_4/XI0/XI0_37/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_10 XI11_4/net21_5_ xsel_37_ XI11_4/XI0/XI0_37/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_9 XI11_4/net21_6_ xsel_37_ XI11_4/XI0/XI0_37/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_8 XI11_4/net21_7_ xsel_37_ XI11_4/XI0/XI0_37/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_7 XI11_4/net21_8_ xsel_37_ XI11_4/XI0/XI0_37/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_6 XI11_4/net21_9_ xsel_37_ XI11_4/XI0/XI0_37/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_5 XI11_4/net21_10_ xsel_37_ XI11_4/XI0/XI0_37/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_4 XI11_4/net21_11_ xsel_37_ XI11_4/XI0/XI0_37/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_3 XI11_4/net21_12_ xsel_37_ XI11_4/XI0/XI0_37/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_2 XI11_4/net21_13_ xsel_37_ XI11_4/XI0/XI0_37/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_1 XI11_4/net21_14_ xsel_37_ XI11_4/XI0/XI0_37/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_0 XI11_4/net21_15_ xsel_37_ XI11_4/XI0/XI0_37/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_15 XI11_4/XI0/XI0_37/d__15_ xsel_37_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_14 XI11_4/XI0/XI0_37/d__14_ xsel_37_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_13 XI11_4/XI0/XI0_37/d__13_ xsel_37_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_12 XI11_4/XI0/XI0_37/d__12_ xsel_37_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_11 XI11_4/XI0/XI0_37/d__11_ xsel_37_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_10 XI11_4/XI0/XI0_37/d__10_ xsel_37_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_9 XI11_4/XI0/XI0_37/d__9_ xsel_37_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_8 XI11_4/XI0/XI0_37/d__8_ xsel_37_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_7 XI11_4/XI0/XI0_37/d__7_ xsel_37_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_6 XI11_4/XI0/XI0_37/d__6_ xsel_37_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_5 XI11_4/XI0/XI0_37/d__5_ xsel_37_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_4 XI11_4/XI0/XI0_37/d__4_ xsel_37_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_3 XI11_4/XI0/XI0_37/d__3_ xsel_37_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_2 XI11_4/XI0/XI0_37/d__2_ xsel_37_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_1 XI11_4/XI0/XI0_37/d__1_ xsel_37_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_0 XI11_4/XI0/XI0_37/d__0_ xsel_37_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_15 XI11_4/net21_0_ xsel_36_ XI11_4/XI0/XI0_36/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_14 XI11_4/net21_1_ xsel_36_ XI11_4/XI0/XI0_36/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_13 XI11_4/net21_2_ xsel_36_ XI11_4/XI0/XI0_36/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_12 XI11_4/net21_3_ xsel_36_ XI11_4/XI0/XI0_36/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_11 XI11_4/net21_4_ xsel_36_ XI11_4/XI0/XI0_36/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_10 XI11_4/net21_5_ xsel_36_ XI11_4/XI0/XI0_36/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_9 XI11_4/net21_6_ xsel_36_ XI11_4/XI0/XI0_36/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_8 XI11_4/net21_7_ xsel_36_ XI11_4/XI0/XI0_36/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_7 XI11_4/net21_8_ xsel_36_ XI11_4/XI0/XI0_36/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_6 XI11_4/net21_9_ xsel_36_ XI11_4/XI0/XI0_36/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_5 XI11_4/net21_10_ xsel_36_ XI11_4/XI0/XI0_36/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_4 XI11_4/net21_11_ xsel_36_ XI11_4/XI0/XI0_36/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_3 XI11_4/net21_12_ xsel_36_ XI11_4/XI0/XI0_36/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_2 XI11_4/net21_13_ xsel_36_ XI11_4/XI0/XI0_36/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_1 XI11_4/net21_14_ xsel_36_ XI11_4/XI0/XI0_36/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_0 XI11_4/net21_15_ xsel_36_ XI11_4/XI0/XI0_36/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_15 XI11_4/XI0/XI0_36/d__15_ xsel_36_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_14 XI11_4/XI0/XI0_36/d__14_ xsel_36_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_13 XI11_4/XI0/XI0_36/d__13_ xsel_36_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_12 XI11_4/XI0/XI0_36/d__12_ xsel_36_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_11 XI11_4/XI0/XI0_36/d__11_ xsel_36_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_10 XI11_4/XI0/XI0_36/d__10_ xsel_36_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_9 XI11_4/XI0/XI0_36/d__9_ xsel_36_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_8 XI11_4/XI0/XI0_36/d__8_ xsel_36_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_7 XI11_4/XI0/XI0_36/d__7_ xsel_36_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_6 XI11_4/XI0/XI0_36/d__6_ xsel_36_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_5 XI11_4/XI0/XI0_36/d__5_ xsel_36_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_4 XI11_4/XI0/XI0_36/d__4_ xsel_36_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_3 XI11_4/XI0/XI0_36/d__3_ xsel_36_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_2 XI11_4/XI0/XI0_36/d__2_ xsel_36_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_1 XI11_4/XI0/XI0_36/d__1_ xsel_36_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_0 XI11_4/XI0/XI0_36/d__0_ xsel_36_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_15 XI11_4/net21_0_ xsel_35_ XI11_4/XI0/XI0_35/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_14 XI11_4/net21_1_ xsel_35_ XI11_4/XI0/XI0_35/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_13 XI11_4/net21_2_ xsel_35_ XI11_4/XI0/XI0_35/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_12 XI11_4/net21_3_ xsel_35_ XI11_4/XI0/XI0_35/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_11 XI11_4/net21_4_ xsel_35_ XI11_4/XI0/XI0_35/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_10 XI11_4/net21_5_ xsel_35_ XI11_4/XI0/XI0_35/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_9 XI11_4/net21_6_ xsel_35_ XI11_4/XI0/XI0_35/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_8 XI11_4/net21_7_ xsel_35_ XI11_4/XI0/XI0_35/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_7 XI11_4/net21_8_ xsel_35_ XI11_4/XI0/XI0_35/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_6 XI11_4/net21_9_ xsel_35_ XI11_4/XI0/XI0_35/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_5 XI11_4/net21_10_ xsel_35_ XI11_4/XI0/XI0_35/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_4 XI11_4/net21_11_ xsel_35_ XI11_4/XI0/XI0_35/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_3 XI11_4/net21_12_ xsel_35_ XI11_4/XI0/XI0_35/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_2 XI11_4/net21_13_ xsel_35_ XI11_4/XI0/XI0_35/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_1 XI11_4/net21_14_ xsel_35_ XI11_4/XI0/XI0_35/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_0 XI11_4/net21_15_ xsel_35_ XI11_4/XI0/XI0_35/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_15 XI11_4/XI0/XI0_35/d__15_ xsel_35_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_14 XI11_4/XI0/XI0_35/d__14_ xsel_35_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_13 XI11_4/XI0/XI0_35/d__13_ xsel_35_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_12 XI11_4/XI0/XI0_35/d__12_ xsel_35_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_11 XI11_4/XI0/XI0_35/d__11_ xsel_35_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_10 XI11_4/XI0/XI0_35/d__10_ xsel_35_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_9 XI11_4/XI0/XI0_35/d__9_ xsel_35_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_8 XI11_4/XI0/XI0_35/d__8_ xsel_35_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_7 XI11_4/XI0/XI0_35/d__7_ xsel_35_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_6 XI11_4/XI0/XI0_35/d__6_ xsel_35_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_5 XI11_4/XI0/XI0_35/d__5_ xsel_35_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_4 XI11_4/XI0/XI0_35/d__4_ xsel_35_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_3 XI11_4/XI0/XI0_35/d__3_ xsel_35_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_2 XI11_4/XI0/XI0_35/d__2_ xsel_35_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_1 XI11_4/XI0/XI0_35/d__1_ xsel_35_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_0 XI11_4/XI0/XI0_35/d__0_ xsel_35_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_15 XI11_4/net21_0_ xsel_34_ XI11_4/XI0/XI0_34/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_14 XI11_4/net21_1_ xsel_34_ XI11_4/XI0/XI0_34/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_13 XI11_4/net21_2_ xsel_34_ XI11_4/XI0/XI0_34/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_12 XI11_4/net21_3_ xsel_34_ XI11_4/XI0/XI0_34/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_11 XI11_4/net21_4_ xsel_34_ XI11_4/XI0/XI0_34/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_10 XI11_4/net21_5_ xsel_34_ XI11_4/XI0/XI0_34/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_9 XI11_4/net21_6_ xsel_34_ XI11_4/XI0/XI0_34/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_8 XI11_4/net21_7_ xsel_34_ XI11_4/XI0/XI0_34/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_7 XI11_4/net21_8_ xsel_34_ XI11_4/XI0/XI0_34/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_6 XI11_4/net21_9_ xsel_34_ XI11_4/XI0/XI0_34/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_5 XI11_4/net21_10_ xsel_34_ XI11_4/XI0/XI0_34/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_4 XI11_4/net21_11_ xsel_34_ XI11_4/XI0/XI0_34/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_3 XI11_4/net21_12_ xsel_34_ XI11_4/XI0/XI0_34/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_2 XI11_4/net21_13_ xsel_34_ XI11_4/XI0/XI0_34/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_1 XI11_4/net21_14_ xsel_34_ XI11_4/XI0/XI0_34/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_0 XI11_4/net21_15_ xsel_34_ XI11_4/XI0/XI0_34/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_15 XI11_4/XI0/XI0_34/d__15_ xsel_34_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_14 XI11_4/XI0/XI0_34/d__14_ xsel_34_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_13 XI11_4/XI0/XI0_34/d__13_ xsel_34_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_12 XI11_4/XI0/XI0_34/d__12_ xsel_34_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_11 XI11_4/XI0/XI0_34/d__11_ xsel_34_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_10 XI11_4/XI0/XI0_34/d__10_ xsel_34_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_9 XI11_4/XI0/XI0_34/d__9_ xsel_34_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_8 XI11_4/XI0/XI0_34/d__8_ xsel_34_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_7 XI11_4/XI0/XI0_34/d__7_ xsel_34_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_6 XI11_4/XI0/XI0_34/d__6_ xsel_34_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_5 XI11_4/XI0/XI0_34/d__5_ xsel_34_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_4 XI11_4/XI0/XI0_34/d__4_ xsel_34_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_3 XI11_4/XI0/XI0_34/d__3_ xsel_34_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_2 XI11_4/XI0/XI0_34/d__2_ xsel_34_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_1 XI11_4/XI0/XI0_34/d__1_ xsel_34_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_0 XI11_4/XI0/XI0_34/d__0_ xsel_34_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_15 XI11_4/net21_0_ xsel_33_ XI11_4/XI0/XI0_33/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_14 XI11_4/net21_1_ xsel_33_ XI11_4/XI0/XI0_33/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_13 XI11_4/net21_2_ xsel_33_ XI11_4/XI0/XI0_33/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_12 XI11_4/net21_3_ xsel_33_ XI11_4/XI0/XI0_33/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_11 XI11_4/net21_4_ xsel_33_ XI11_4/XI0/XI0_33/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_10 XI11_4/net21_5_ xsel_33_ XI11_4/XI0/XI0_33/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_9 XI11_4/net21_6_ xsel_33_ XI11_4/XI0/XI0_33/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_8 XI11_4/net21_7_ xsel_33_ XI11_4/XI0/XI0_33/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_7 XI11_4/net21_8_ xsel_33_ XI11_4/XI0/XI0_33/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_6 XI11_4/net21_9_ xsel_33_ XI11_4/XI0/XI0_33/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_5 XI11_4/net21_10_ xsel_33_ XI11_4/XI0/XI0_33/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_4 XI11_4/net21_11_ xsel_33_ XI11_4/XI0/XI0_33/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_3 XI11_4/net21_12_ xsel_33_ XI11_4/XI0/XI0_33/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_2 XI11_4/net21_13_ xsel_33_ XI11_4/XI0/XI0_33/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_1 XI11_4/net21_14_ xsel_33_ XI11_4/XI0/XI0_33/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_0 XI11_4/net21_15_ xsel_33_ XI11_4/XI0/XI0_33/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_15 XI11_4/XI0/XI0_33/d__15_ xsel_33_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_14 XI11_4/XI0/XI0_33/d__14_ xsel_33_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_13 XI11_4/XI0/XI0_33/d__13_ xsel_33_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_12 XI11_4/XI0/XI0_33/d__12_ xsel_33_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_11 XI11_4/XI0/XI0_33/d__11_ xsel_33_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_10 XI11_4/XI0/XI0_33/d__10_ xsel_33_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_9 XI11_4/XI0/XI0_33/d__9_ xsel_33_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_8 XI11_4/XI0/XI0_33/d__8_ xsel_33_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_7 XI11_4/XI0/XI0_33/d__7_ xsel_33_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_6 XI11_4/XI0/XI0_33/d__6_ xsel_33_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_5 XI11_4/XI0/XI0_33/d__5_ xsel_33_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_4 XI11_4/XI0/XI0_33/d__4_ xsel_33_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_3 XI11_4/XI0/XI0_33/d__3_ xsel_33_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_2 XI11_4/XI0/XI0_33/d__2_ xsel_33_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_1 XI11_4/XI0/XI0_33/d__1_ xsel_33_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_0 XI11_4/XI0/XI0_33/d__0_ xsel_33_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_15 XI11_4/net21_0_ xsel_32_ XI11_4/XI0/XI0_32/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_14 XI11_4/net21_1_ xsel_32_ XI11_4/XI0/XI0_32/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_13 XI11_4/net21_2_ xsel_32_ XI11_4/XI0/XI0_32/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_12 XI11_4/net21_3_ xsel_32_ XI11_4/XI0/XI0_32/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_11 XI11_4/net21_4_ xsel_32_ XI11_4/XI0/XI0_32/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_10 XI11_4/net21_5_ xsel_32_ XI11_4/XI0/XI0_32/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_9 XI11_4/net21_6_ xsel_32_ XI11_4/XI0/XI0_32/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_8 XI11_4/net21_7_ xsel_32_ XI11_4/XI0/XI0_32/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_7 XI11_4/net21_8_ xsel_32_ XI11_4/XI0/XI0_32/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_6 XI11_4/net21_9_ xsel_32_ XI11_4/XI0/XI0_32/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_5 XI11_4/net21_10_ xsel_32_ XI11_4/XI0/XI0_32/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_4 XI11_4/net21_11_ xsel_32_ XI11_4/XI0/XI0_32/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_3 XI11_4/net21_12_ xsel_32_ XI11_4/XI0/XI0_32/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_2 XI11_4/net21_13_ xsel_32_ XI11_4/XI0/XI0_32/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_1 XI11_4/net21_14_ xsel_32_ XI11_4/XI0/XI0_32/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_0 XI11_4/net21_15_ xsel_32_ XI11_4/XI0/XI0_32/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_15 XI11_4/XI0/XI0_32/d__15_ xsel_32_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_14 XI11_4/XI0/XI0_32/d__14_ xsel_32_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_13 XI11_4/XI0/XI0_32/d__13_ xsel_32_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_12 XI11_4/XI0/XI0_32/d__12_ xsel_32_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_11 XI11_4/XI0/XI0_32/d__11_ xsel_32_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_10 XI11_4/XI0/XI0_32/d__10_ xsel_32_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_9 XI11_4/XI0/XI0_32/d__9_ xsel_32_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_8 XI11_4/XI0/XI0_32/d__8_ xsel_32_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_7 XI11_4/XI0/XI0_32/d__7_ xsel_32_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_6 XI11_4/XI0/XI0_32/d__6_ xsel_32_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_5 XI11_4/XI0/XI0_32/d__5_ xsel_32_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_4 XI11_4/XI0/XI0_32/d__4_ xsel_32_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_3 XI11_4/XI0/XI0_32/d__3_ xsel_32_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_2 XI11_4/XI0/XI0_32/d__2_ xsel_32_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_1 XI11_4/XI0/XI0_32/d__1_ xsel_32_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_0 XI11_4/XI0/XI0_32/d__0_ xsel_32_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_15 XI11_4/net21_0_ xsel_31_ XI11_4/XI0/XI0_31/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_14 XI11_4/net21_1_ xsel_31_ XI11_4/XI0/XI0_31/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_13 XI11_4/net21_2_ xsel_31_ XI11_4/XI0/XI0_31/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_12 XI11_4/net21_3_ xsel_31_ XI11_4/XI0/XI0_31/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_11 XI11_4/net21_4_ xsel_31_ XI11_4/XI0/XI0_31/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_10 XI11_4/net21_5_ xsel_31_ XI11_4/XI0/XI0_31/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_9 XI11_4/net21_6_ xsel_31_ XI11_4/XI0/XI0_31/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_8 XI11_4/net21_7_ xsel_31_ XI11_4/XI0/XI0_31/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_7 XI11_4/net21_8_ xsel_31_ XI11_4/XI0/XI0_31/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_6 XI11_4/net21_9_ xsel_31_ XI11_4/XI0/XI0_31/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_5 XI11_4/net21_10_ xsel_31_ XI11_4/XI0/XI0_31/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_4 XI11_4/net21_11_ xsel_31_ XI11_4/XI0/XI0_31/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_3 XI11_4/net21_12_ xsel_31_ XI11_4/XI0/XI0_31/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_2 XI11_4/net21_13_ xsel_31_ XI11_4/XI0/XI0_31/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_1 XI11_4/net21_14_ xsel_31_ XI11_4/XI0/XI0_31/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_0 XI11_4/net21_15_ xsel_31_ XI11_4/XI0/XI0_31/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_15 XI11_4/XI0/XI0_31/d__15_ xsel_31_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_14 XI11_4/XI0/XI0_31/d__14_ xsel_31_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_13 XI11_4/XI0/XI0_31/d__13_ xsel_31_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_12 XI11_4/XI0/XI0_31/d__12_ xsel_31_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_11 XI11_4/XI0/XI0_31/d__11_ xsel_31_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_10 XI11_4/XI0/XI0_31/d__10_ xsel_31_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_9 XI11_4/XI0/XI0_31/d__9_ xsel_31_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_8 XI11_4/XI0/XI0_31/d__8_ xsel_31_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_7 XI11_4/XI0/XI0_31/d__7_ xsel_31_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_6 XI11_4/XI0/XI0_31/d__6_ xsel_31_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_5 XI11_4/XI0/XI0_31/d__5_ xsel_31_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_4 XI11_4/XI0/XI0_31/d__4_ xsel_31_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_3 XI11_4/XI0/XI0_31/d__3_ xsel_31_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_2 XI11_4/XI0/XI0_31/d__2_ xsel_31_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_1 XI11_4/XI0/XI0_31/d__1_ xsel_31_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_0 XI11_4/XI0/XI0_31/d__0_ xsel_31_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_15 XI11_4/net21_0_ xsel_30_ XI11_4/XI0/XI0_30/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_14 XI11_4/net21_1_ xsel_30_ XI11_4/XI0/XI0_30/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_13 XI11_4/net21_2_ xsel_30_ XI11_4/XI0/XI0_30/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_12 XI11_4/net21_3_ xsel_30_ XI11_4/XI0/XI0_30/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_11 XI11_4/net21_4_ xsel_30_ XI11_4/XI0/XI0_30/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_10 XI11_4/net21_5_ xsel_30_ XI11_4/XI0/XI0_30/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_9 XI11_4/net21_6_ xsel_30_ XI11_4/XI0/XI0_30/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_8 XI11_4/net21_7_ xsel_30_ XI11_4/XI0/XI0_30/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_7 XI11_4/net21_8_ xsel_30_ XI11_4/XI0/XI0_30/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_6 XI11_4/net21_9_ xsel_30_ XI11_4/XI0/XI0_30/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_5 XI11_4/net21_10_ xsel_30_ XI11_4/XI0/XI0_30/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_4 XI11_4/net21_11_ xsel_30_ XI11_4/XI0/XI0_30/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_3 XI11_4/net21_12_ xsel_30_ XI11_4/XI0/XI0_30/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_2 XI11_4/net21_13_ xsel_30_ XI11_4/XI0/XI0_30/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_1 XI11_4/net21_14_ xsel_30_ XI11_4/XI0/XI0_30/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_0 XI11_4/net21_15_ xsel_30_ XI11_4/XI0/XI0_30/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_15 XI11_4/XI0/XI0_30/d__15_ xsel_30_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_14 XI11_4/XI0/XI0_30/d__14_ xsel_30_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_13 XI11_4/XI0/XI0_30/d__13_ xsel_30_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_12 XI11_4/XI0/XI0_30/d__12_ xsel_30_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_11 XI11_4/XI0/XI0_30/d__11_ xsel_30_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_10 XI11_4/XI0/XI0_30/d__10_ xsel_30_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_9 XI11_4/XI0/XI0_30/d__9_ xsel_30_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_8 XI11_4/XI0/XI0_30/d__8_ xsel_30_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_7 XI11_4/XI0/XI0_30/d__7_ xsel_30_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_6 XI11_4/XI0/XI0_30/d__6_ xsel_30_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_5 XI11_4/XI0/XI0_30/d__5_ xsel_30_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_4 XI11_4/XI0/XI0_30/d__4_ xsel_30_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_3 XI11_4/XI0/XI0_30/d__3_ xsel_30_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_2 XI11_4/XI0/XI0_30/d__2_ xsel_30_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_1 XI11_4/XI0/XI0_30/d__1_ xsel_30_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_0 XI11_4/XI0/XI0_30/d__0_ xsel_30_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_15 XI11_4/net21_0_ xsel_29_ XI11_4/XI0/XI0_29/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_14 XI11_4/net21_1_ xsel_29_ XI11_4/XI0/XI0_29/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_13 XI11_4/net21_2_ xsel_29_ XI11_4/XI0/XI0_29/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_12 XI11_4/net21_3_ xsel_29_ XI11_4/XI0/XI0_29/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_11 XI11_4/net21_4_ xsel_29_ XI11_4/XI0/XI0_29/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_10 XI11_4/net21_5_ xsel_29_ XI11_4/XI0/XI0_29/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_9 XI11_4/net21_6_ xsel_29_ XI11_4/XI0/XI0_29/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_8 XI11_4/net21_7_ xsel_29_ XI11_4/XI0/XI0_29/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_7 XI11_4/net21_8_ xsel_29_ XI11_4/XI0/XI0_29/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_6 XI11_4/net21_9_ xsel_29_ XI11_4/XI0/XI0_29/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_5 XI11_4/net21_10_ xsel_29_ XI11_4/XI0/XI0_29/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_4 XI11_4/net21_11_ xsel_29_ XI11_4/XI0/XI0_29/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_3 XI11_4/net21_12_ xsel_29_ XI11_4/XI0/XI0_29/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_2 XI11_4/net21_13_ xsel_29_ XI11_4/XI0/XI0_29/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_1 XI11_4/net21_14_ xsel_29_ XI11_4/XI0/XI0_29/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_0 XI11_4/net21_15_ xsel_29_ XI11_4/XI0/XI0_29/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_15 XI11_4/XI0/XI0_29/d__15_ xsel_29_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_14 XI11_4/XI0/XI0_29/d__14_ xsel_29_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_13 XI11_4/XI0/XI0_29/d__13_ xsel_29_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_12 XI11_4/XI0/XI0_29/d__12_ xsel_29_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_11 XI11_4/XI0/XI0_29/d__11_ xsel_29_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_10 XI11_4/XI0/XI0_29/d__10_ xsel_29_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_9 XI11_4/XI0/XI0_29/d__9_ xsel_29_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_8 XI11_4/XI0/XI0_29/d__8_ xsel_29_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_7 XI11_4/XI0/XI0_29/d__7_ xsel_29_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_6 XI11_4/XI0/XI0_29/d__6_ xsel_29_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_5 XI11_4/XI0/XI0_29/d__5_ xsel_29_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_4 XI11_4/XI0/XI0_29/d__4_ xsel_29_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_3 XI11_4/XI0/XI0_29/d__3_ xsel_29_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_2 XI11_4/XI0/XI0_29/d__2_ xsel_29_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_1 XI11_4/XI0/XI0_29/d__1_ xsel_29_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_0 XI11_4/XI0/XI0_29/d__0_ xsel_29_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_15 XI11_4/net21_0_ xsel_28_ XI11_4/XI0/XI0_28/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_14 XI11_4/net21_1_ xsel_28_ XI11_4/XI0/XI0_28/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_13 XI11_4/net21_2_ xsel_28_ XI11_4/XI0/XI0_28/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_12 XI11_4/net21_3_ xsel_28_ XI11_4/XI0/XI0_28/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_11 XI11_4/net21_4_ xsel_28_ XI11_4/XI0/XI0_28/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_10 XI11_4/net21_5_ xsel_28_ XI11_4/XI0/XI0_28/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_9 XI11_4/net21_6_ xsel_28_ XI11_4/XI0/XI0_28/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_8 XI11_4/net21_7_ xsel_28_ XI11_4/XI0/XI0_28/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_7 XI11_4/net21_8_ xsel_28_ XI11_4/XI0/XI0_28/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_6 XI11_4/net21_9_ xsel_28_ XI11_4/XI0/XI0_28/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_5 XI11_4/net21_10_ xsel_28_ XI11_4/XI0/XI0_28/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_4 XI11_4/net21_11_ xsel_28_ XI11_4/XI0/XI0_28/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_3 XI11_4/net21_12_ xsel_28_ XI11_4/XI0/XI0_28/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_2 XI11_4/net21_13_ xsel_28_ XI11_4/XI0/XI0_28/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_1 XI11_4/net21_14_ xsel_28_ XI11_4/XI0/XI0_28/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_0 XI11_4/net21_15_ xsel_28_ XI11_4/XI0/XI0_28/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_15 XI11_4/XI0/XI0_28/d__15_ xsel_28_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_14 XI11_4/XI0/XI0_28/d__14_ xsel_28_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_13 XI11_4/XI0/XI0_28/d__13_ xsel_28_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_12 XI11_4/XI0/XI0_28/d__12_ xsel_28_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_11 XI11_4/XI0/XI0_28/d__11_ xsel_28_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_10 XI11_4/XI0/XI0_28/d__10_ xsel_28_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_9 XI11_4/XI0/XI0_28/d__9_ xsel_28_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_8 XI11_4/XI0/XI0_28/d__8_ xsel_28_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_7 XI11_4/XI0/XI0_28/d__7_ xsel_28_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_6 XI11_4/XI0/XI0_28/d__6_ xsel_28_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_5 XI11_4/XI0/XI0_28/d__5_ xsel_28_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_4 XI11_4/XI0/XI0_28/d__4_ xsel_28_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_3 XI11_4/XI0/XI0_28/d__3_ xsel_28_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_2 XI11_4/XI0/XI0_28/d__2_ xsel_28_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_1 XI11_4/XI0/XI0_28/d__1_ xsel_28_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_0 XI11_4/XI0/XI0_28/d__0_ xsel_28_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_15 XI11_4/net21_0_ xsel_27_ XI11_4/XI0/XI0_27/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_14 XI11_4/net21_1_ xsel_27_ XI11_4/XI0/XI0_27/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_13 XI11_4/net21_2_ xsel_27_ XI11_4/XI0/XI0_27/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_12 XI11_4/net21_3_ xsel_27_ XI11_4/XI0/XI0_27/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_11 XI11_4/net21_4_ xsel_27_ XI11_4/XI0/XI0_27/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_10 XI11_4/net21_5_ xsel_27_ XI11_4/XI0/XI0_27/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_9 XI11_4/net21_6_ xsel_27_ XI11_4/XI0/XI0_27/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_8 XI11_4/net21_7_ xsel_27_ XI11_4/XI0/XI0_27/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_7 XI11_4/net21_8_ xsel_27_ XI11_4/XI0/XI0_27/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_6 XI11_4/net21_9_ xsel_27_ XI11_4/XI0/XI0_27/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_5 XI11_4/net21_10_ xsel_27_ XI11_4/XI0/XI0_27/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_4 XI11_4/net21_11_ xsel_27_ XI11_4/XI0/XI0_27/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_3 XI11_4/net21_12_ xsel_27_ XI11_4/XI0/XI0_27/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_2 XI11_4/net21_13_ xsel_27_ XI11_4/XI0/XI0_27/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_1 XI11_4/net21_14_ xsel_27_ XI11_4/XI0/XI0_27/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_0 XI11_4/net21_15_ xsel_27_ XI11_4/XI0/XI0_27/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_15 XI11_4/XI0/XI0_27/d__15_ xsel_27_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_14 XI11_4/XI0/XI0_27/d__14_ xsel_27_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_13 XI11_4/XI0/XI0_27/d__13_ xsel_27_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_12 XI11_4/XI0/XI0_27/d__12_ xsel_27_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_11 XI11_4/XI0/XI0_27/d__11_ xsel_27_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_10 XI11_4/XI0/XI0_27/d__10_ xsel_27_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_9 XI11_4/XI0/XI0_27/d__9_ xsel_27_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_8 XI11_4/XI0/XI0_27/d__8_ xsel_27_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_7 XI11_4/XI0/XI0_27/d__7_ xsel_27_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_6 XI11_4/XI0/XI0_27/d__6_ xsel_27_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_5 XI11_4/XI0/XI0_27/d__5_ xsel_27_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_4 XI11_4/XI0/XI0_27/d__4_ xsel_27_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_3 XI11_4/XI0/XI0_27/d__3_ xsel_27_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_2 XI11_4/XI0/XI0_27/d__2_ xsel_27_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_1 XI11_4/XI0/XI0_27/d__1_ xsel_27_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_0 XI11_4/XI0/XI0_27/d__0_ xsel_27_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_15 XI11_4/net21_0_ xsel_26_ XI11_4/XI0/XI0_26/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_14 XI11_4/net21_1_ xsel_26_ XI11_4/XI0/XI0_26/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_13 XI11_4/net21_2_ xsel_26_ XI11_4/XI0/XI0_26/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_12 XI11_4/net21_3_ xsel_26_ XI11_4/XI0/XI0_26/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_11 XI11_4/net21_4_ xsel_26_ XI11_4/XI0/XI0_26/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_10 XI11_4/net21_5_ xsel_26_ XI11_4/XI0/XI0_26/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_9 XI11_4/net21_6_ xsel_26_ XI11_4/XI0/XI0_26/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_8 XI11_4/net21_7_ xsel_26_ XI11_4/XI0/XI0_26/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_7 XI11_4/net21_8_ xsel_26_ XI11_4/XI0/XI0_26/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_6 XI11_4/net21_9_ xsel_26_ XI11_4/XI0/XI0_26/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_5 XI11_4/net21_10_ xsel_26_ XI11_4/XI0/XI0_26/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_4 XI11_4/net21_11_ xsel_26_ XI11_4/XI0/XI0_26/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_3 XI11_4/net21_12_ xsel_26_ XI11_4/XI0/XI0_26/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_2 XI11_4/net21_13_ xsel_26_ XI11_4/XI0/XI0_26/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_1 XI11_4/net21_14_ xsel_26_ XI11_4/XI0/XI0_26/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_0 XI11_4/net21_15_ xsel_26_ XI11_4/XI0/XI0_26/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_15 XI11_4/XI0/XI0_26/d__15_ xsel_26_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_14 XI11_4/XI0/XI0_26/d__14_ xsel_26_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_13 XI11_4/XI0/XI0_26/d__13_ xsel_26_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_12 XI11_4/XI0/XI0_26/d__12_ xsel_26_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_11 XI11_4/XI0/XI0_26/d__11_ xsel_26_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_10 XI11_4/XI0/XI0_26/d__10_ xsel_26_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_9 XI11_4/XI0/XI0_26/d__9_ xsel_26_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_8 XI11_4/XI0/XI0_26/d__8_ xsel_26_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_7 XI11_4/XI0/XI0_26/d__7_ xsel_26_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_6 XI11_4/XI0/XI0_26/d__6_ xsel_26_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_5 XI11_4/XI0/XI0_26/d__5_ xsel_26_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_4 XI11_4/XI0/XI0_26/d__4_ xsel_26_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_3 XI11_4/XI0/XI0_26/d__3_ xsel_26_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_2 XI11_4/XI0/XI0_26/d__2_ xsel_26_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_1 XI11_4/XI0/XI0_26/d__1_ xsel_26_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_0 XI11_4/XI0/XI0_26/d__0_ xsel_26_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_15 XI11_4/net21_0_ xsel_25_ XI11_4/XI0/XI0_25/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_14 XI11_4/net21_1_ xsel_25_ XI11_4/XI0/XI0_25/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_13 XI11_4/net21_2_ xsel_25_ XI11_4/XI0/XI0_25/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_12 XI11_4/net21_3_ xsel_25_ XI11_4/XI0/XI0_25/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_11 XI11_4/net21_4_ xsel_25_ XI11_4/XI0/XI0_25/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_10 XI11_4/net21_5_ xsel_25_ XI11_4/XI0/XI0_25/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_9 XI11_4/net21_6_ xsel_25_ XI11_4/XI0/XI0_25/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_8 XI11_4/net21_7_ xsel_25_ XI11_4/XI0/XI0_25/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_7 XI11_4/net21_8_ xsel_25_ XI11_4/XI0/XI0_25/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_6 XI11_4/net21_9_ xsel_25_ XI11_4/XI0/XI0_25/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_5 XI11_4/net21_10_ xsel_25_ XI11_4/XI0/XI0_25/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_4 XI11_4/net21_11_ xsel_25_ XI11_4/XI0/XI0_25/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_3 XI11_4/net21_12_ xsel_25_ XI11_4/XI0/XI0_25/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_2 XI11_4/net21_13_ xsel_25_ XI11_4/XI0/XI0_25/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_1 XI11_4/net21_14_ xsel_25_ XI11_4/XI0/XI0_25/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_0 XI11_4/net21_15_ xsel_25_ XI11_4/XI0/XI0_25/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_15 XI11_4/XI0/XI0_25/d__15_ xsel_25_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_14 XI11_4/XI0/XI0_25/d__14_ xsel_25_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_13 XI11_4/XI0/XI0_25/d__13_ xsel_25_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_12 XI11_4/XI0/XI0_25/d__12_ xsel_25_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_11 XI11_4/XI0/XI0_25/d__11_ xsel_25_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_10 XI11_4/XI0/XI0_25/d__10_ xsel_25_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_9 XI11_4/XI0/XI0_25/d__9_ xsel_25_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_8 XI11_4/XI0/XI0_25/d__8_ xsel_25_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_7 XI11_4/XI0/XI0_25/d__7_ xsel_25_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_6 XI11_4/XI0/XI0_25/d__6_ xsel_25_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_5 XI11_4/XI0/XI0_25/d__5_ xsel_25_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_4 XI11_4/XI0/XI0_25/d__4_ xsel_25_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_3 XI11_4/XI0/XI0_25/d__3_ xsel_25_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_2 XI11_4/XI0/XI0_25/d__2_ xsel_25_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_1 XI11_4/XI0/XI0_25/d__1_ xsel_25_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_0 XI11_4/XI0/XI0_25/d__0_ xsel_25_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_15 XI11_4/net21_0_ xsel_24_ XI11_4/XI0/XI0_24/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_14 XI11_4/net21_1_ xsel_24_ XI11_4/XI0/XI0_24/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_13 XI11_4/net21_2_ xsel_24_ XI11_4/XI0/XI0_24/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_12 XI11_4/net21_3_ xsel_24_ XI11_4/XI0/XI0_24/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_11 XI11_4/net21_4_ xsel_24_ XI11_4/XI0/XI0_24/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_10 XI11_4/net21_5_ xsel_24_ XI11_4/XI0/XI0_24/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_9 XI11_4/net21_6_ xsel_24_ XI11_4/XI0/XI0_24/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_8 XI11_4/net21_7_ xsel_24_ XI11_4/XI0/XI0_24/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_7 XI11_4/net21_8_ xsel_24_ XI11_4/XI0/XI0_24/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_6 XI11_4/net21_9_ xsel_24_ XI11_4/XI0/XI0_24/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_5 XI11_4/net21_10_ xsel_24_ XI11_4/XI0/XI0_24/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_4 XI11_4/net21_11_ xsel_24_ XI11_4/XI0/XI0_24/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_3 XI11_4/net21_12_ xsel_24_ XI11_4/XI0/XI0_24/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_2 XI11_4/net21_13_ xsel_24_ XI11_4/XI0/XI0_24/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_1 XI11_4/net21_14_ xsel_24_ XI11_4/XI0/XI0_24/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_0 XI11_4/net21_15_ xsel_24_ XI11_4/XI0/XI0_24/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_15 XI11_4/XI0/XI0_24/d__15_ xsel_24_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_14 XI11_4/XI0/XI0_24/d__14_ xsel_24_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_13 XI11_4/XI0/XI0_24/d__13_ xsel_24_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_12 XI11_4/XI0/XI0_24/d__12_ xsel_24_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_11 XI11_4/XI0/XI0_24/d__11_ xsel_24_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_10 XI11_4/XI0/XI0_24/d__10_ xsel_24_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_9 XI11_4/XI0/XI0_24/d__9_ xsel_24_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_8 XI11_4/XI0/XI0_24/d__8_ xsel_24_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_7 XI11_4/XI0/XI0_24/d__7_ xsel_24_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_6 XI11_4/XI0/XI0_24/d__6_ xsel_24_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_5 XI11_4/XI0/XI0_24/d__5_ xsel_24_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_4 XI11_4/XI0/XI0_24/d__4_ xsel_24_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_3 XI11_4/XI0/XI0_24/d__3_ xsel_24_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_2 XI11_4/XI0/XI0_24/d__2_ xsel_24_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_1 XI11_4/XI0/XI0_24/d__1_ xsel_24_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_0 XI11_4/XI0/XI0_24/d__0_ xsel_24_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_15 XI11_4/net21_0_ xsel_23_ XI11_4/XI0/XI0_23/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_14 XI11_4/net21_1_ xsel_23_ XI11_4/XI0/XI0_23/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_13 XI11_4/net21_2_ xsel_23_ XI11_4/XI0/XI0_23/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_12 XI11_4/net21_3_ xsel_23_ XI11_4/XI0/XI0_23/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_11 XI11_4/net21_4_ xsel_23_ XI11_4/XI0/XI0_23/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_10 XI11_4/net21_5_ xsel_23_ XI11_4/XI0/XI0_23/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_9 XI11_4/net21_6_ xsel_23_ XI11_4/XI0/XI0_23/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_8 XI11_4/net21_7_ xsel_23_ XI11_4/XI0/XI0_23/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_7 XI11_4/net21_8_ xsel_23_ XI11_4/XI0/XI0_23/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_6 XI11_4/net21_9_ xsel_23_ XI11_4/XI0/XI0_23/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_5 XI11_4/net21_10_ xsel_23_ XI11_4/XI0/XI0_23/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_4 XI11_4/net21_11_ xsel_23_ XI11_4/XI0/XI0_23/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_3 XI11_4/net21_12_ xsel_23_ XI11_4/XI0/XI0_23/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_2 XI11_4/net21_13_ xsel_23_ XI11_4/XI0/XI0_23/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_1 XI11_4/net21_14_ xsel_23_ XI11_4/XI0/XI0_23/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_0 XI11_4/net21_15_ xsel_23_ XI11_4/XI0/XI0_23/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_15 XI11_4/XI0/XI0_23/d__15_ xsel_23_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_14 XI11_4/XI0/XI0_23/d__14_ xsel_23_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_13 XI11_4/XI0/XI0_23/d__13_ xsel_23_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_12 XI11_4/XI0/XI0_23/d__12_ xsel_23_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_11 XI11_4/XI0/XI0_23/d__11_ xsel_23_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_10 XI11_4/XI0/XI0_23/d__10_ xsel_23_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_9 XI11_4/XI0/XI0_23/d__9_ xsel_23_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_8 XI11_4/XI0/XI0_23/d__8_ xsel_23_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_7 XI11_4/XI0/XI0_23/d__7_ xsel_23_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_6 XI11_4/XI0/XI0_23/d__6_ xsel_23_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_5 XI11_4/XI0/XI0_23/d__5_ xsel_23_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_4 XI11_4/XI0/XI0_23/d__4_ xsel_23_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_3 XI11_4/XI0/XI0_23/d__3_ xsel_23_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_2 XI11_4/XI0/XI0_23/d__2_ xsel_23_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_1 XI11_4/XI0/XI0_23/d__1_ xsel_23_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_0 XI11_4/XI0/XI0_23/d__0_ xsel_23_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_15 XI11_4/net21_0_ xsel_22_ XI11_4/XI0/XI0_22/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_14 XI11_4/net21_1_ xsel_22_ XI11_4/XI0/XI0_22/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_13 XI11_4/net21_2_ xsel_22_ XI11_4/XI0/XI0_22/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_12 XI11_4/net21_3_ xsel_22_ XI11_4/XI0/XI0_22/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_11 XI11_4/net21_4_ xsel_22_ XI11_4/XI0/XI0_22/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_10 XI11_4/net21_5_ xsel_22_ XI11_4/XI0/XI0_22/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_9 XI11_4/net21_6_ xsel_22_ XI11_4/XI0/XI0_22/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_8 XI11_4/net21_7_ xsel_22_ XI11_4/XI0/XI0_22/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_7 XI11_4/net21_8_ xsel_22_ XI11_4/XI0/XI0_22/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_6 XI11_4/net21_9_ xsel_22_ XI11_4/XI0/XI0_22/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_5 XI11_4/net21_10_ xsel_22_ XI11_4/XI0/XI0_22/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_4 XI11_4/net21_11_ xsel_22_ XI11_4/XI0/XI0_22/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_3 XI11_4/net21_12_ xsel_22_ XI11_4/XI0/XI0_22/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_2 XI11_4/net21_13_ xsel_22_ XI11_4/XI0/XI0_22/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_1 XI11_4/net21_14_ xsel_22_ XI11_4/XI0/XI0_22/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_0 XI11_4/net21_15_ xsel_22_ XI11_4/XI0/XI0_22/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_15 XI11_4/XI0/XI0_22/d__15_ xsel_22_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_14 XI11_4/XI0/XI0_22/d__14_ xsel_22_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_13 XI11_4/XI0/XI0_22/d__13_ xsel_22_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_12 XI11_4/XI0/XI0_22/d__12_ xsel_22_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_11 XI11_4/XI0/XI0_22/d__11_ xsel_22_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_10 XI11_4/XI0/XI0_22/d__10_ xsel_22_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_9 XI11_4/XI0/XI0_22/d__9_ xsel_22_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_8 XI11_4/XI0/XI0_22/d__8_ xsel_22_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_7 XI11_4/XI0/XI0_22/d__7_ xsel_22_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_6 XI11_4/XI0/XI0_22/d__6_ xsel_22_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_5 XI11_4/XI0/XI0_22/d__5_ xsel_22_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_4 XI11_4/XI0/XI0_22/d__4_ xsel_22_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_3 XI11_4/XI0/XI0_22/d__3_ xsel_22_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_2 XI11_4/XI0/XI0_22/d__2_ xsel_22_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_1 XI11_4/XI0/XI0_22/d__1_ xsel_22_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_0 XI11_4/XI0/XI0_22/d__0_ xsel_22_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_15 XI11_4/net21_0_ xsel_21_ XI11_4/XI0/XI0_21/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_14 XI11_4/net21_1_ xsel_21_ XI11_4/XI0/XI0_21/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_13 XI11_4/net21_2_ xsel_21_ XI11_4/XI0/XI0_21/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_12 XI11_4/net21_3_ xsel_21_ XI11_4/XI0/XI0_21/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_11 XI11_4/net21_4_ xsel_21_ XI11_4/XI0/XI0_21/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_10 XI11_4/net21_5_ xsel_21_ XI11_4/XI0/XI0_21/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_9 XI11_4/net21_6_ xsel_21_ XI11_4/XI0/XI0_21/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_8 XI11_4/net21_7_ xsel_21_ XI11_4/XI0/XI0_21/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_7 XI11_4/net21_8_ xsel_21_ XI11_4/XI0/XI0_21/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_6 XI11_4/net21_9_ xsel_21_ XI11_4/XI0/XI0_21/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_5 XI11_4/net21_10_ xsel_21_ XI11_4/XI0/XI0_21/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_4 XI11_4/net21_11_ xsel_21_ XI11_4/XI0/XI0_21/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_3 XI11_4/net21_12_ xsel_21_ XI11_4/XI0/XI0_21/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_2 XI11_4/net21_13_ xsel_21_ XI11_4/XI0/XI0_21/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_1 XI11_4/net21_14_ xsel_21_ XI11_4/XI0/XI0_21/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_0 XI11_4/net21_15_ xsel_21_ XI11_4/XI0/XI0_21/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_15 XI11_4/XI0/XI0_21/d__15_ xsel_21_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_14 XI11_4/XI0/XI0_21/d__14_ xsel_21_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_13 XI11_4/XI0/XI0_21/d__13_ xsel_21_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_12 XI11_4/XI0/XI0_21/d__12_ xsel_21_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_11 XI11_4/XI0/XI0_21/d__11_ xsel_21_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_10 XI11_4/XI0/XI0_21/d__10_ xsel_21_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_9 XI11_4/XI0/XI0_21/d__9_ xsel_21_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_8 XI11_4/XI0/XI0_21/d__8_ xsel_21_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_7 XI11_4/XI0/XI0_21/d__7_ xsel_21_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_6 XI11_4/XI0/XI0_21/d__6_ xsel_21_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_5 XI11_4/XI0/XI0_21/d__5_ xsel_21_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_4 XI11_4/XI0/XI0_21/d__4_ xsel_21_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_3 XI11_4/XI0/XI0_21/d__3_ xsel_21_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_2 XI11_4/XI0/XI0_21/d__2_ xsel_21_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_1 XI11_4/XI0/XI0_21/d__1_ xsel_21_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_0 XI11_4/XI0/XI0_21/d__0_ xsel_21_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_15 XI11_4/net21_0_ xsel_20_ XI11_4/XI0/XI0_20/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_14 XI11_4/net21_1_ xsel_20_ XI11_4/XI0/XI0_20/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_13 XI11_4/net21_2_ xsel_20_ XI11_4/XI0/XI0_20/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_12 XI11_4/net21_3_ xsel_20_ XI11_4/XI0/XI0_20/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_11 XI11_4/net21_4_ xsel_20_ XI11_4/XI0/XI0_20/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_10 XI11_4/net21_5_ xsel_20_ XI11_4/XI0/XI0_20/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_9 XI11_4/net21_6_ xsel_20_ XI11_4/XI0/XI0_20/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_8 XI11_4/net21_7_ xsel_20_ XI11_4/XI0/XI0_20/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_7 XI11_4/net21_8_ xsel_20_ XI11_4/XI0/XI0_20/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_6 XI11_4/net21_9_ xsel_20_ XI11_4/XI0/XI0_20/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_5 XI11_4/net21_10_ xsel_20_ XI11_4/XI0/XI0_20/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_4 XI11_4/net21_11_ xsel_20_ XI11_4/XI0/XI0_20/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_3 XI11_4/net21_12_ xsel_20_ XI11_4/XI0/XI0_20/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_2 XI11_4/net21_13_ xsel_20_ XI11_4/XI0/XI0_20/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_1 XI11_4/net21_14_ xsel_20_ XI11_4/XI0/XI0_20/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_0 XI11_4/net21_15_ xsel_20_ XI11_4/XI0/XI0_20/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_15 XI11_4/XI0/XI0_20/d__15_ xsel_20_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_14 XI11_4/XI0/XI0_20/d__14_ xsel_20_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_13 XI11_4/XI0/XI0_20/d__13_ xsel_20_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_12 XI11_4/XI0/XI0_20/d__12_ xsel_20_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_11 XI11_4/XI0/XI0_20/d__11_ xsel_20_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_10 XI11_4/XI0/XI0_20/d__10_ xsel_20_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_9 XI11_4/XI0/XI0_20/d__9_ xsel_20_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_8 XI11_4/XI0/XI0_20/d__8_ xsel_20_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_7 XI11_4/XI0/XI0_20/d__7_ xsel_20_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_6 XI11_4/XI0/XI0_20/d__6_ xsel_20_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_5 XI11_4/XI0/XI0_20/d__5_ xsel_20_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_4 XI11_4/XI0/XI0_20/d__4_ xsel_20_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_3 XI11_4/XI0/XI0_20/d__3_ xsel_20_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_2 XI11_4/XI0/XI0_20/d__2_ xsel_20_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_1 XI11_4/XI0/XI0_20/d__1_ xsel_20_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_0 XI11_4/XI0/XI0_20/d__0_ xsel_20_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_15 XI11_4/net21_0_ xsel_19_ XI11_4/XI0/XI0_19/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_14 XI11_4/net21_1_ xsel_19_ XI11_4/XI0/XI0_19/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_13 XI11_4/net21_2_ xsel_19_ XI11_4/XI0/XI0_19/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_12 XI11_4/net21_3_ xsel_19_ XI11_4/XI0/XI0_19/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_11 XI11_4/net21_4_ xsel_19_ XI11_4/XI0/XI0_19/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_10 XI11_4/net21_5_ xsel_19_ XI11_4/XI0/XI0_19/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_9 XI11_4/net21_6_ xsel_19_ XI11_4/XI0/XI0_19/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_8 XI11_4/net21_7_ xsel_19_ XI11_4/XI0/XI0_19/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_7 XI11_4/net21_8_ xsel_19_ XI11_4/XI0/XI0_19/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_6 XI11_4/net21_9_ xsel_19_ XI11_4/XI0/XI0_19/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_5 XI11_4/net21_10_ xsel_19_ XI11_4/XI0/XI0_19/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_4 XI11_4/net21_11_ xsel_19_ XI11_4/XI0/XI0_19/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_3 XI11_4/net21_12_ xsel_19_ XI11_4/XI0/XI0_19/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_2 XI11_4/net21_13_ xsel_19_ XI11_4/XI0/XI0_19/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_1 XI11_4/net21_14_ xsel_19_ XI11_4/XI0/XI0_19/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_0 XI11_4/net21_15_ xsel_19_ XI11_4/XI0/XI0_19/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_15 XI11_4/XI0/XI0_19/d__15_ xsel_19_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_14 XI11_4/XI0/XI0_19/d__14_ xsel_19_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_13 XI11_4/XI0/XI0_19/d__13_ xsel_19_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_12 XI11_4/XI0/XI0_19/d__12_ xsel_19_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_11 XI11_4/XI0/XI0_19/d__11_ xsel_19_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_10 XI11_4/XI0/XI0_19/d__10_ xsel_19_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_9 XI11_4/XI0/XI0_19/d__9_ xsel_19_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_8 XI11_4/XI0/XI0_19/d__8_ xsel_19_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_7 XI11_4/XI0/XI0_19/d__7_ xsel_19_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_6 XI11_4/XI0/XI0_19/d__6_ xsel_19_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_5 XI11_4/XI0/XI0_19/d__5_ xsel_19_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_4 XI11_4/XI0/XI0_19/d__4_ xsel_19_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_3 XI11_4/XI0/XI0_19/d__3_ xsel_19_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_2 XI11_4/XI0/XI0_19/d__2_ xsel_19_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_1 XI11_4/XI0/XI0_19/d__1_ xsel_19_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_0 XI11_4/XI0/XI0_19/d__0_ xsel_19_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_15 XI11_4/net21_0_ xsel_18_ XI11_4/XI0/XI0_18/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_14 XI11_4/net21_1_ xsel_18_ XI11_4/XI0/XI0_18/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_13 XI11_4/net21_2_ xsel_18_ XI11_4/XI0/XI0_18/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_12 XI11_4/net21_3_ xsel_18_ XI11_4/XI0/XI0_18/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_11 XI11_4/net21_4_ xsel_18_ XI11_4/XI0/XI0_18/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_10 XI11_4/net21_5_ xsel_18_ XI11_4/XI0/XI0_18/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_9 XI11_4/net21_6_ xsel_18_ XI11_4/XI0/XI0_18/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_8 XI11_4/net21_7_ xsel_18_ XI11_4/XI0/XI0_18/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_7 XI11_4/net21_8_ xsel_18_ XI11_4/XI0/XI0_18/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_6 XI11_4/net21_9_ xsel_18_ XI11_4/XI0/XI0_18/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_5 XI11_4/net21_10_ xsel_18_ XI11_4/XI0/XI0_18/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_4 XI11_4/net21_11_ xsel_18_ XI11_4/XI0/XI0_18/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_3 XI11_4/net21_12_ xsel_18_ XI11_4/XI0/XI0_18/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_2 XI11_4/net21_13_ xsel_18_ XI11_4/XI0/XI0_18/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_1 XI11_4/net21_14_ xsel_18_ XI11_4/XI0/XI0_18/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_0 XI11_4/net21_15_ xsel_18_ XI11_4/XI0/XI0_18/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_15 XI11_4/XI0/XI0_18/d__15_ xsel_18_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_14 XI11_4/XI0/XI0_18/d__14_ xsel_18_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_13 XI11_4/XI0/XI0_18/d__13_ xsel_18_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_12 XI11_4/XI0/XI0_18/d__12_ xsel_18_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_11 XI11_4/XI0/XI0_18/d__11_ xsel_18_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_10 XI11_4/XI0/XI0_18/d__10_ xsel_18_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_9 XI11_4/XI0/XI0_18/d__9_ xsel_18_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_8 XI11_4/XI0/XI0_18/d__8_ xsel_18_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_7 XI11_4/XI0/XI0_18/d__7_ xsel_18_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_6 XI11_4/XI0/XI0_18/d__6_ xsel_18_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_5 XI11_4/XI0/XI0_18/d__5_ xsel_18_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_4 XI11_4/XI0/XI0_18/d__4_ xsel_18_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_3 XI11_4/XI0/XI0_18/d__3_ xsel_18_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_2 XI11_4/XI0/XI0_18/d__2_ xsel_18_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_1 XI11_4/XI0/XI0_18/d__1_ xsel_18_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_0 XI11_4/XI0/XI0_18/d__0_ xsel_18_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_15 XI11_4/net21_0_ xsel_17_ XI11_4/XI0/XI0_17/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_14 XI11_4/net21_1_ xsel_17_ XI11_4/XI0/XI0_17/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_13 XI11_4/net21_2_ xsel_17_ XI11_4/XI0/XI0_17/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_12 XI11_4/net21_3_ xsel_17_ XI11_4/XI0/XI0_17/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_11 XI11_4/net21_4_ xsel_17_ XI11_4/XI0/XI0_17/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_10 XI11_4/net21_5_ xsel_17_ XI11_4/XI0/XI0_17/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_9 XI11_4/net21_6_ xsel_17_ XI11_4/XI0/XI0_17/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_8 XI11_4/net21_7_ xsel_17_ XI11_4/XI0/XI0_17/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_7 XI11_4/net21_8_ xsel_17_ XI11_4/XI0/XI0_17/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_6 XI11_4/net21_9_ xsel_17_ XI11_4/XI0/XI0_17/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_5 XI11_4/net21_10_ xsel_17_ XI11_4/XI0/XI0_17/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_4 XI11_4/net21_11_ xsel_17_ XI11_4/XI0/XI0_17/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_3 XI11_4/net21_12_ xsel_17_ XI11_4/XI0/XI0_17/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_2 XI11_4/net21_13_ xsel_17_ XI11_4/XI0/XI0_17/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_1 XI11_4/net21_14_ xsel_17_ XI11_4/XI0/XI0_17/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_0 XI11_4/net21_15_ xsel_17_ XI11_4/XI0/XI0_17/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_15 XI11_4/XI0/XI0_17/d__15_ xsel_17_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_14 XI11_4/XI0/XI0_17/d__14_ xsel_17_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_13 XI11_4/XI0/XI0_17/d__13_ xsel_17_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_12 XI11_4/XI0/XI0_17/d__12_ xsel_17_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_11 XI11_4/XI0/XI0_17/d__11_ xsel_17_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_10 XI11_4/XI0/XI0_17/d__10_ xsel_17_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_9 XI11_4/XI0/XI0_17/d__9_ xsel_17_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_8 XI11_4/XI0/XI0_17/d__8_ xsel_17_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_7 XI11_4/XI0/XI0_17/d__7_ xsel_17_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_6 XI11_4/XI0/XI0_17/d__6_ xsel_17_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_5 XI11_4/XI0/XI0_17/d__5_ xsel_17_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_4 XI11_4/XI0/XI0_17/d__4_ xsel_17_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_3 XI11_4/XI0/XI0_17/d__3_ xsel_17_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_2 XI11_4/XI0/XI0_17/d__2_ xsel_17_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_1 XI11_4/XI0/XI0_17/d__1_ xsel_17_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_0 XI11_4/XI0/XI0_17/d__0_ xsel_17_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_15 XI11_4/net21_0_ xsel_16_ XI11_4/XI0/XI0_16/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_14 XI11_4/net21_1_ xsel_16_ XI11_4/XI0/XI0_16/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_13 XI11_4/net21_2_ xsel_16_ XI11_4/XI0/XI0_16/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_12 XI11_4/net21_3_ xsel_16_ XI11_4/XI0/XI0_16/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_11 XI11_4/net21_4_ xsel_16_ XI11_4/XI0/XI0_16/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_10 XI11_4/net21_5_ xsel_16_ XI11_4/XI0/XI0_16/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_9 XI11_4/net21_6_ xsel_16_ XI11_4/XI0/XI0_16/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_8 XI11_4/net21_7_ xsel_16_ XI11_4/XI0/XI0_16/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_7 XI11_4/net21_8_ xsel_16_ XI11_4/XI0/XI0_16/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_6 XI11_4/net21_9_ xsel_16_ XI11_4/XI0/XI0_16/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_5 XI11_4/net21_10_ xsel_16_ XI11_4/XI0/XI0_16/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_4 XI11_4/net21_11_ xsel_16_ XI11_4/XI0/XI0_16/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_3 XI11_4/net21_12_ xsel_16_ XI11_4/XI0/XI0_16/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_2 XI11_4/net21_13_ xsel_16_ XI11_4/XI0/XI0_16/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_1 XI11_4/net21_14_ xsel_16_ XI11_4/XI0/XI0_16/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_0 XI11_4/net21_15_ xsel_16_ XI11_4/XI0/XI0_16/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_15 XI11_4/XI0/XI0_16/d__15_ xsel_16_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_14 XI11_4/XI0/XI0_16/d__14_ xsel_16_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_13 XI11_4/XI0/XI0_16/d__13_ xsel_16_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_12 XI11_4/XI0/XI0_16/d__12_ xsel_16_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_11 XI11_4/XI0/XI0_16/d__11_ xsel_16_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_10 XI11_4/XI0/XI0_16/d__10_ xsel_16_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_9 XI11_4/XI0/XI0_16/d__9_ xsel_16_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_8 XI11_4/XI0/XI0_16/d__8_ xsel_16_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_7 XI11_4/XI0/XI0_16/d__7_ xsel_16_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_6 XI11_4/XI0/XI0_16/d__6_ xsel_16_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_5 XI11_4/XI0/XI0_16/d__5_ xsel_16_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_4 XI11_4/XI0/XI0_16/d__4_ xsel_16_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_3 XI11_4/XI0/XI0_16/d__3_ xsel_16_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_2 XI11_4/XI0/XI0_16/d__2_ xsel_16_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_1 XI11_4/XI0/XI0_16/d__1_ xsel_16_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_0 XI11_4/XI0/XI0_16/d__0_ xsel_16_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_15 XI11_4/net21_0_ xsel_15_ XI11_4/XI0/XI0_15/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_14 XI11_4/net21_1_ xsel_15_ XI11_4/XI0/XI0_15/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_13 XI11_4/net21_2_ xsel_15_ XI11_4/XI0/XI0_15/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_12 XI11_4/net21_3_ xsel_15_ XI11_4/XI0/XI0_15/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_11 XI11_4/net21_4_ xsel_15_ XI11_4/XI0/XI0_15/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_10 XI11_4/net21_5_ xsel_15_ XI11_4/XI0/XI0_15/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_9 XI11_4/net21_6_ xsel_15_ XI11_4/XI0/XI0_15/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_8 XI11_4/net21_7_ xsel_15_ XI11_4/XI0/XI0_15/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_7 XI11_4/net21_8_ xsel_15_ XI11_4/XI0/XI0_15/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_6 XI11_4/net21_9_ xsel_15_ XI11_4/XI0/XI0_15/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_5 XI11_4/net21_10_ xsel_15_ XI11_4/XI0/XI0_15/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_4 XI11_4/net21_11_ xsel_15_ XI11_4/XI0/XI0_15/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_3 XI11_4/net21_12_ xsel_15_ XI11_4/XI0/XI0_15/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_2 XI11_4/net21_13_ xsel_15_ XI11_4/XI0/XI0_15/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_1 XI11_4/net21_14_ xsel_15_ XI11_4/XI0/XI0_15/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_0 XI11_4/net21_15_ xsel_15_ XI11_4/XI0/XI0_15/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_15 XI11_4/XI0/XI0_15/d__15_ xsel_15_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_14 XI11_4/XI0/XI0_15/d__14_ xsel_15_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_13 XI11_4/XI0/XI0_15/d__13_ xsel_15_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_12 XI11_4/XI0/XI0_15/d__12_ xsel_15_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_11 XI11_4/XI0/XI0_15/d__11_ xsel_15_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_10 XI11_4/XI0/XI0_15/d__10_ xsel_15_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_9 XI11_4/XI0/XI0_15/d__9_ xsel_15_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_8 XI11_4/XI0/XI0_15/d__8_ xsel_15_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_7 XI11_4/XI0/XI0_15/d__7_ xsel_15_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_6 XI11_4/XI0/XI0_15/d__6_ xsel_15_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_5 XI11_4/XI0/XI0_15/d__5_ xsel_15_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_4 XI11_4/XI0/XI0_15/d__4_ xsel_15_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_3 XI11_4/XI0/XI0_15/d__3_ xsel_15_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_2 XI11_4/XI0/XI0_15/d__2_ xsel_15_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_1 XI11_4/XI0/XI0_15/d__1_ xsel_15_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_0 XI11_4/XI0/XI0_15/d__0_ xsel_15_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_15 XI11_4/net21_0_ xsel_14_ XI11_4/XI0/XI0_14/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_14 XI11_4/net21_1_ xsel_14_ XI11_4/XI0/XI0_14/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_13 XI11_4/net21_2_ xsel_14_ XI11_4/XI0/XI0_14/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_12 XI11_4/net21_3_ xsel_14_ XI11_4/XI0/XI0_14/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_11 XI11_4/net21_4_ xsel_14_ XI11_4/XI0/XI0_14/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_10 XI11_4/net21_5_ xsel_14_ XI11_4/XI0/XI0_14/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_9 XI11_4/net21_6_ xsel_14_ XI11_4/XI0/XI0_14/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_8 XI11_4/net21_7_ xsel_14_ XI11_4/XI0/XI0_14/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_7 XI11_4/net21_8_ xsel_14_ XI11_4/XI0/XI0_14/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_6 XI11_4/net21_9_ xsel_14_ XI11_4/XI0/XI0_14/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_5 XI11_4/net21_10_ xsel_14_ XI11_4/XI0/XI0_14/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_4 XI11_4/net21_11_ xsel_14_ XI11_4/XI0/XI0_14/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_3 XI11_4/net21_12_ xsel_14_ XI11_4/XI0/XI0_14/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_2 XI11_4/net21_13_ xsel_14_ XI11_4/XI0/XI0_14/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_1 XI11_4/net21_14_ xsel_14_ XI11_4/XI0/XI0_14/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_0 XI11_4/net21_15_ xsel_14_ XI11_4/XI0/XI0_14/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_15 XI11_4/XI0/XI0_14/d__15_ xsel_14_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_14 XI11_4/XI0/XI0_14/d__14_ xsel_14_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_13 XI11_4/XI0/XI0_14/d__13_ xsel_14_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_12 XI11_4/XI0/XI0_14/d__12_ xsel_14_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_11 XI11_4/XI0/XI0_14/d__11_ xsel_14_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_10 XI11_4/XI0/XI0_14/d__10_ xsel_14_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_9 XI11_4/XI0/XI0_14/d__9_ xsel_14_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_8 XI11_4/XI0/XI0_14/d__8_ xsel_14_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_7 XI11_4/XI0/XI0_14/d__7_ xsel_14_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_6 XI11_4/XI0/XI0_14/d__6_ xsel_14_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_5 XI11_4/XI0/XI0_14/d__5_ xsel_14_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_4 XI11_4/XI0/XI0_14/d__4_ xsel_14_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_3 XI11_4/XI0/XI0_14/d__3_ xsel_14_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_2 XI11_4/XI0/XI0_14/d__2_ xsel_14_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_1 XI11_4/XI0/XI0_14/d__1_ xsel_14_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_0 XI11_4/XI0/XI0_14/d__0_ xsel_14_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_15 XI11_4/net21_0_ xsel_13_ XI11_4/XI0/XI0_13/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_14 XI11_4/net21_1_ xsel_13_ XI11_4/XI0/XI0_13/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_13 XI11_4/net21_2_ xsel_13_ XI11_4/XI0/XI0_13/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_12 XI11_4/net21_3_ xsel_13_ XI11_4/XI0/XI0_13/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_11 XI11_4/net21_4_ xsel_13_ XI11_4/XI0/XI0_13/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_10 XI11_4/net21_5_ xsel_13_ XI11_4/XI0/XI0_13/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_9 XI11_4/net21_6_ xsel_13_ XI11_4/XI0/XI0_13/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_8 XI11_4/net21_7_ xsel_13_ XI11_4/XI0/XI0_13/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_7 XI11_4/net21_8_ xsel_13_ XI11_4/XI0/XI0_13/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_6 XI11_4/net21_9_ xsel_13_ XI11_4/XI0/XI0_13/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_5 XI11_4/net21_10_ xsel_13_ XI11_4/XI0/XI0_13/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_4 XI11_4/net21_11_ xsel_13_ XI11_4/XI0/XI0_13/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_3 XI11_4/net21_12_ xsel_13_ XI11_4/XI0/XI0_13/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_2 XI11_4/net21_13_ xsel_13_ XI11_4/XI0/XI0_13/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_1 XI11_4/net21_14_ xsel_13_ XI11_4/XI0/XI0_13/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_0 XI11_4/net21_15_ xsel_13_ XI11_4/XI0/XI0_13/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_15 XI11_4/XI0/XI0_13/d__15_ xsel_13_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_14 XI11_4/XI0/XI0_13/d__14_ xsel_13_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_13 XI11_4/XI0/XI0_13/d__13_ xsel_13_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_12 XI11_4/XI0/XI0_13/d__12_ xsel_13_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_11 XI11_4/XI0/XI0_13/d__11_ xsel_13_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_10 XI11_4/XI0/XI0_13/d__10_ xsel_13_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_9 XI11_4/XI0/XI0_13/d__9_ xsel_13_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_8 XI11_4/XI0/XI0_13/d__8_ xsel_13_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_7 XI11_4/XI0/XI0_13/d__7_ xsel_13_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_6 XI11_4/XI0/XI0_13/d__6_ xsel_13_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_5 XI11_4/XI0/XI0_13/d__5_ xsel_13_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_4 XI11_4/XI0/XI0_13/d__4_ xsel_13_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_3 XI11_4/XI0/XI0_13/d__3_ xsel_13_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_2 XI11_4/XI0/XI0_13/d__2_ xsel_13_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_1 XI11_4/XI0/XI0_13/d__1_ xsel_13_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_0 XI11_4/XI0/XI0_13/d__0_ xsel_13_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_15 XI11_4/net21_0_ xsel_12_ XI11_4/XI0/XI0_12/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_14 XI11_4/net21_1_ xsel_12_ XI11_4/XI0/XI0_12/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_13 XI11_4/net21_2_ xsel_12_ XI11_4/XI0/XI0_12/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_12 XI11_4/net21_3_ xsel_12_ XI11_4/XI0/XI0_12/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_11 XI11_4/net21_4_ xsel_12_ XI11_4/XI0/XI0_12/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_10 XI11_4/net21_5_ xsel_12_ XI11_4/XI0/XI0_12/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_9 XI11_4/net21_6_ xsel_12_ XI11_4/XI0/XI0_12/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_8 XI11_4/net21_7_ xsel_12_ XI11_4/XI0/XI0_12/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_7 XI11_4/net21_8_ xsel_12_ XI11_4/XI0/XI0_12/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_6 XI11_4/net21_9_ xsel_12_ XI11_4/XI0/XI0_12/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_5 XI11_4/net21_10_ xsel_12_ XI11_4/XI0/XI0_12/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_4 XI11_4/net21_11_ xsel_12_ XI11_4/XI0/XI0_12/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_3 XI11_4/net21_12_ xsel_12_ XI11_4/XI0/XI0_12/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_2 XI11_4/net21_13_ xsel_12_ XI11_4/XI0/XI0_12/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_1 XI11_4/net21_14_ xsel_12_ XI11_4/XI0/XI0_12/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_0 XI11_4/net21_15_ xsel_12_ XI11_4/XI0/XI0_12/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_15 XI11_4/XI0/XI0_12/d__15_ xsel_12_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_14 XI11_4/XI0/XI0_12/d__14_ xsel_12_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_13 XI11_4/XI0/XI0_12/d__13_ xsel_12_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_12 XI11_4/XI0/XI0_12/d__12_ xsel_12_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_11 XI11_4/XI0/XI0_12/d__11_ xsel_12_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_10 XI11_4/XI0/XI0_12/d__10_ xsel_12_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_9 XI11_4/XI0/XI0_12/d__9_ xsel_12_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_8 XI11_4/XI0/XI0_12/d__8_ xsel_12_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_7 XI11_4/XI0/XI0_12/d__7_ xsel_12_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_6 XI11_4/XI0/XI0_12/d__6_ xsel_12_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_5 XI11_4/XI0/XI0_12/d__5_ xsel_12_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_4 XI11_4/XI0/XI0_12/d__4_ xsel_12_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_3 XI11_4/XI0/XI0_12/d__3_ xsel_12_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_2 XI11_4/XI0/XI0_12/d__2_ xsel_12_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_1 XI11_4/XI0/XI0_12/d__1_ xsel_12_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_0 XI11_4/XI0/XI0_12/d__0_ xsel_12_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_15 XI11_4/net21_0_ xsel_11_ XI11_4/XI0/XI0_11/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_14 XI11_4/net21_1_ xsel_11_ XI11_4/XI0/XI0_11/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_13 XI11_4/net21_2_ xsel_11_ XI11_4/XI0/XI0_11/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_12 XI11_4/net21_3_ xsel_11_ XI11_4/XI0/XI0_11/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_11 XI11_4/net21_4_ xsel_11_ XI11_4/XI0/XI0_11/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_10 XI11_4/net21_5_ xsel_11_ XI11_4/XI0/XI0_11/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_9 XI11_4/net21_6_ xsel_11_ XI11_4/XI0/XI0_11/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_8 XI11_4/net21_7_ xsel_11_ XI11_4/XI0/XI0_11/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_7 XI11_4/net21_8_ xsel_11_ XI11_4/XI0/XI0_11/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_6 XI11_4/net21_9_ xsel_11_ XI11_4/XI0/XI0_11/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_5 XI11_4/net21_10_ xsel_11_ XI11_4/XI0/XI0_11/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_4 XI11_4/net21_11_ xsel_11_ XI11_4/XI0/XI0_11/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_3 XI11_4/net21_12_ xsel_11_ XI11_4/XI0/XI0_11/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_2 XI11_4/net21_13_ xsel_11_ XI11_4/XI0/XI0_11/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_1 XI11_4/net21_14_ xsel_11_ XI11_4/XI0/XI0_11/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_0 XI11_4/net21_15_ xsel_11_ XI11_4/XI0/XI0_11/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_15 XI11_4/XI0/XI0_11/d__15_ xsel_11_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_14 XI11_4/XI0/XI0_11/d__14_ xsel_11_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_13 XI11_4/XI0/XI0_11/d__13_ xsel_11_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_12 XI11_4/XI0/XI0_11/d__12_ xsel_11_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_11 XI11_4/XI0/XI0_11/d__11_ xsel_11_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_10 XI11_4/XI0/XI0_11/d__10_ xsel_11_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_9 XI11_4/XI0/XI0_11/d__9_ xsel_11_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_8 XI11_4/XI0/XI0_11/d__8_ xsel_11_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_7 XI11_4/XI0/XI0_11/d__7_ xsel_11_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_6 XI11_4/XI0/XI0_11/d__6_ xsel_11_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_5 XI11_4/XI0/XI0_11/d__5_ xsel_11_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_4 XI11_4/XI0/XI0_11/d__4_ xsel_11_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_3 XI11_4/XI0/XI0_11/d__3_ xsel_11_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_2 XI11_4/XI0/XI0_11/d__2_ xsel_11_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_1 XI11_4/XI0/XI0_11/d__1_ xsel_11_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_0 XI11_4/XI0/XI0_11/d__0_ xsel_11_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_15 XI11_4/net21_0_ xsel_10_ XI11_4/XI0/XI0_10/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_14 XI11_4/net21_1_ xsel_10_ XI11_4/XI0/XI0_10/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_13 XI11_4/net21_2_ xsel_10_ XI11_4/XI0/XI0_10/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_12 XI11_4/net21_3_ xsel_10_ XI11_4/XI0/XI0_10/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_11 XI11_4/net21_4_ xsel_10_ XI11_4/XI0/XI0_10/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_10 XI11_4/net21_5_ xsel_10_ XI11_4/XI0/XI0_10/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_9 XI11_4/net21_6_ xsel_10_ XI11_4/XI0/XI0_10/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_8 XI11_4/net21_7_ xsel_10_ XI11_4/XI0/XI0_10/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_7 XI11_4/net21_8_ xsel_10_ XI11_4/XI0/XI0_10/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_6 XI11_4/net21_9_ xsel_10_ XI11_4/XI0/XI0_10/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_5 XI11_4/net21_10_ xsel_10_ XI11_4/XI0/XI0_10/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_4 XI11_4/net21_11_ xsel_10_ XI11_4/XI0/XI0_10/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_3 XI11_4/net21_12_ xsel_10_ XI11_4/XI0/XI0_10/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_2 XI11_4/net21_13_ xsel_10_ XI11_4/XI0/XI0_10/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_1 XI11_4/net21_14_ xsel_10_ XI11_4/XI0/XI0_10/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_0 XI11_4/net21_15_ xsel_10_ XI11_4/XI0/XI0_10/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_15 XI11_4/XI0/XI0_10/d__15_ xsel_10_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_14 XI11_4/XI0/XI0_10/d__14_ xsel_10_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_13 XI11_4/XI0/XI0_10/d__13_ xsel_10_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_12 XI11_4/XI0/XI0_10/d__12_ xsel_10_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_11 XI11_4/XI0/XI0_10/d__11_ xsel_10_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_10 XI11_4/XI0/XI0_10/d__10_ xsel_10_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_9 XI11_4/XI0/XI0_10/d__9_ xsel_10_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_8 XI11_4/XI0/XI0_10/d__8_ xsel_10_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_7 XI11_4/XI0/XI0_10/d__7_ xsel_10_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_6 XI11_4/XI0/XI0_10/d__6_ xsel_10_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_5 XI11_4/XI0/XI0_10/d__5_ xsel_10_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_4 XI11_4/XI0/XI0_10/d__4_ xsel_10_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_3 XI11_4/XI0/XI0_10/d__3_ xsel_10_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_2 XI11_4/XI0/XI0_10/d__2_ xsel_10_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_1 XI11_4/XI0/XI0_10/d__1_ xsel_10_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_0 XI11_4/XI0/XI0_10/d__0_ xsel_10_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_15 XI11_4/net21_0_ xsel_9_ XI11_4/XI0/XI0_9/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_14 XI11_4/net21_1_ xsel_9_ XI11_4/XI0/XI0_9/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_13 XI11_4/net21_2_ xsel_9_ XI11_4/XI0/XI0_9/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_12 XI11_4/net21_3_ xsel_9_ XI11_4/XI0/XI0_9/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_11 XI11_4/net21_4_ xsel_9_ XI11_4/XI0/XI0_9/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_10 XI11_4/net21_5_ xsel_9_ XI11_4/XI0/XI0_9/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_9 XI11_4/net21_6_ xsel_9_ XI11_4/XI0/XI0_9/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_8 XI11_4/net21_7_ xsel_9_ XI11_4/XI0/XI0_9/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_7 XI11_4/net21_8_ xsel_9_ XI11_4/XI0/XI0_9/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_6 XI11_4/net21_9_ xsel_9_ XI11_4/XI0/XI0_9/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_5 XI11_4/net21_10_ xsel_9_ XI11_4/XI0/XI0_9/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_4 XI11_4/net21_11_ xsel_9_ XI11_4/XI0/XI0_9/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_3 XI11_4/net21_12_ xsel_9_ XI11_4/XI0/XI0_9/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_2 XI11_4/net21_13_ xsel_9_ XI11_4/XI0/XI0_9/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_1 XI11_4/net21_14_ xsel_9_ XI11_4/XI0/XI0_9/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_0 XI11_4/net21_15_ xsel_9_ XI11_4/XI0/XI0_9/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_15 XI11_4/XI0/XI0_9/d__15_ xsel_9_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_14 XI11_4/XI0/XI0_9/d__14_ xsel_9_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_13 XI11_4/XI0/XI0_9/d__13_ xsel_9_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_12 XI11_4/XI0/XI0_9/d__12_ xsel_9_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_11 XI11_4/XI0/XI0_9/d__11_ xsel_9_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_10 XI11_4/XI0/XI0_9/d__10_ xsel_9_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_9 XI11_4/XI0/XI0_9/d__9_ xsel_9_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_8 XI11_4/XI0/XI0_9/d__8_ xsel_9_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_7 XI11_4/XI0/XI0_9/d__7_ xsel_9_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_6 XI11_4/XI0/XI0_9/d__6_ xsel_9_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_5 XI11_4/XI0/XI0_9/d__5_ xsel_9_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_4 XI11_4/XI0/XI0_9/d__4_ xsel_9_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_3 XI11_4/XI0/XI0_9/d__3_ xsel_9_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_2 XI11_4/XI0/XI0_9/d__2_ xsel_9_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_1 XI11_4/XI0/XI0_9/d__1_ xsel_9_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_0 XI11_4/XI0/XI0_9/d__0_ xsel_9_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_15 XI11_4/net21_0_ xsel_8_ XI11_4/XI0/XI0_8/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_14 XI11_4/net21_1_ xsel_8_ XI11_4/XI0/XI0_8/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_13 XI11_4/net21_2_ xsel_8_ XI11_4/XI0/XI0_8/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_12 XI11_4/net21_3_ xsel_8_ XI11_4/XI0/XI0_8/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_11 XI11_4/net21_4_ xsel_8_ XI11_4/XI0/XI0_8/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_10 XI11_4/net21_5_ xsel_8_ XI11_4/XI0/XI0_8/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_9 XI11_4/net21_6_ xsel_8_ XI11_4/XI0/XI0_8/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_8 XI11_4/net21_7_ xsel_8_ XI11_4/XI0/XI0_8/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_7 XI11_4/net21_8_ xsel_8_ XI11_4/XI0/XI0_8/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_6 XI11_4/net21_9_ xsel_8_ XI11_4/XI0/XI0_8/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_5 XI11_4/net21_10_ xsel_8_ XI11_4/XI0/XI0_8/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_4 XI11_4/net21_11_ xsel_8_ XI11_4/XI0/XI0_8/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_3 XI11_4/net21_12_ xsel_8_ XI11_4/XI0/XI0_8/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_2 XI11_4/net21_13_ xsel_8_ XI11_4/XI0/XI0_8/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_1 XI11_4/net21_14_ xsel_8_ XI11_4/XI0/XI0_8/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_0 XI11_4/net21_15_ xsel_8_ XI11_4/XI0/XI0_8/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_15 XI11_4/XI0/XI0_8/d__15_ xsel_8_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_14 XI11_4/XI0/XI0_8/d__14_ xsel_8_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_13 XI11_4/XI0/XI0_8/d__13_ xsel_8_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_12 XI11_4/XI0/XI0_8/d__12_ xsel_8_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_11 XI11_4/XI0/XI0_8/d__11_ xsel_8_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_10 XI11_4/XI0/XI0_8/d__10_ xsel_8_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_9 XI11_4/XI0/XI0_8/d__9_ xsel_8_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_8 XI11_4/XI0/XI0_8/d__8_ xsel_8_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_7 XI11_4/XI0/XI0_8/d__7_ xsel_8_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_6 XI11_4/XI0/XI0_8/d__6_ xsel_8_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_5 XI11_4/XI0/XI0_8/d__5_ xsel_8_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_4 XI11_4/XI0/XI0_8/d__4_ xsel_8_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_3 XI11_4/XI0/XI0_8/d__3_ xsel_8_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_2 XI11_4/XI0/XI0_8/d__2_ xsel_8_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_1 XI11_4/XI0/XI0_8/d__1_ xsel_8_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_0 XI11_4/XI0/XI0_8/d__0_ xsel_8_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_15 XI11_4/net21_0_ xsel_7_ XI11_4/XI0/XI0_7/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_14 XI11_4/net21_1_ xsel_7_ XI11_4/XI0/XI0_7/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_13 XI11_4/net21_2_ xsel_7_ XI11_4/XI0/XI0_7/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_12 XI11_4/net21_3_ xsel_7_ XI11_4/XI0/XI0_7/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_11 XI11_4/net21_4_ xsel_7_ XI11_4/XI0/XI0_7/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_10 XI11_4/net21_5_ xsel_7_ XI11_4/XI0/XI0_7/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_9 XI11_4/net21_6_ xsel_7_ XI11_4/XI0/XI0_7/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_8 XI11_4/net21_7_ xsel_7_ XI11_4/XI0/XI0_7/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_7 XI11_4/net21_8_ xsel_7_ XI11_4/XI0/XI0_7/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_6 XI11_4/net21_9_ xsel_7_ XI11_4/XI0/XI0_7/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_5 XI11_4/net21_10_ xsel_7_ XI11_4/XI0/XI0_7/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_4 XI11_4/net21_11_ xsel_7_ XI11_4/XI0/XI0_7/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_3 XI11_4/net21_12_ xsel_7_ XI11_4/XI0/XI0_7/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_2 XI11_4/net21_13_ xsel_7_ XI11_4/XI0/XI0_7/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_1 XI11_4/net21_14_ xsel_7_ XI11_4/XI0/XI0_7/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_0 XI11_4/net21_15_ xsel_7_ XI11_4/XI0/XI0_7/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_15 XI11_4/XI0/XI0_7/d__15_ xsel_7_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_14 XI11_4/XI0/XI0_7/d__14_ xsel_7_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_13 XI11_4/XI0/XI0_7/d__13_ xsel_7_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_12 XI11_4/XI0/XI0_7/d__12_ xsel_7_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_11 XI11_4/XI0/XI0_7/d__11_ xsel_7_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_10 XI11_4/XI0/XI0_7/d__10_ xsel_7_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_9 XI11_4/XI0/XI0_7/d__9_ xsel_7_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_8 XI11_4/XI0/XI0_7/d__8_ xsel_7_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_7 XI11_4/XI0/XI0_7/d__7_ xsel_7_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_6 XI11_4/XI0/XI0_7/d__6_ xsel_7_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_5 XI11_4/XI0/XI0_7/d__5_ xsel_7_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_4 XI11_4/XI0/XI0_7/d__4_ xsel_7_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_3 XI11_4/XI0/XI0_7/d__3_ xsel_7_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_2 XI11_4/XI0/XI0_7/d__2_ xsel_7_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_1 XI11_4/XI0/XI0_7/d__1_ xsel_7_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_0 XI11_4/XI0/XI0_7/d__0_ xsel_7_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_15 XI11_4/net21_0_ xsel_6_ XI11_4/XI0/XI0_6/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_14 XI11_4/net21_1_ xsel_6_ XI11_4/XI0/XI0_6/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_13 XI11_4/net21_2_ xsel_6_ XI11_4/XI0/XI0_6/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_12 XI11_4/net21_3_ xsel_6_ XI11_4/XI0/XI0_6/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_11 XI11_4/net21_4_ xsel_6_ XI11_4/XI0/XI0_6/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_10 XI11_4/net21_5_ xsel_6_ XI11_4/XI0/XI0_6/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_9 XI11_4/net21_6_ xsel_6_ XI11_4/XI0/XI0_6/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_8 XI11_4/net21_7_ xsel_6_ XI11_4/XI0/XI0_6/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_7 XI11_4/net21_8_ xsel_6_ XI11_4/XI0/XI0_6/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_6 XI11_4/net21_9_ xsel_6_ XI11_4/XI0/XI0_6/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_5 XI11_4/net21_10_ xsel_6_ XI11_4/XI0/XI0_6/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_4 XI11_4/net21_11_ xsel_6_ XI11_4/XI0/XI0_6/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_3 XI11_4/net21_12_ xsel_6_ XI11_4/XI0/XI0_6/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_2 XI11_4/net21_13_ xsel_6_ XI11_4/XI0/XI0_6/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_1 XI11_4/net21_14_ xsel_6_ XI11_4/XI0/XI0_6/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_0 XI11_4/net21_15_ xsel_6_ XI11_4/XI0/XI0_6/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_15 XI11_4/XI0/XI0_6/d__15_ xsel_6_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_14 XI11_4/XI0/XI0_6/d__14_ xsel_6_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_13 XI11_4/XI0/XI0_6/d__13_ xsel_6_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_12 XI11_4/XI0/XI0_6/d__12_ xsel_6_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_11 XI11_4/XI0/XI0_6/d__11_ xsel_6_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_10 XI11_4/XI0/XI0_6/d__10_ xsel_6_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_9 XI11_4/XI0/XI0_6/d__9_ xsel_6_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_8 XI11_4/XI0/XI0_6/d__8_ xsel_6_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_7 XI11_4/XI0/XI0_6/d__7_ xsel_6_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_6 XI11_4/XI0/XI0_6/d__6_ xsel_6_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_5 XI11_4/XI0/XI0_6/d__5_ xsel_6_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_4 XI11_4/XI0/XI0_6/d__4_ xsel_6_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_3 XI11_4/XI0/XI0_6/d__3_ xsel_6_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_2 XI11_4/XI0/XI0_6/d__2_ xsel_6_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_1 XI11_4/XI0/XI0_6/d__1_ xsel_6_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_0 XI11_4/XI0/XI0_6/d__0_ xsel_6_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_15 XI11_4/net21_0_ xsel_5_ XI11_4/XI0/XI0_5/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_14 XI11_4/net21_1_ xsel_5_ XI11_4/XI0/XI0_5/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_13 XI11_4/net21_2_ xsel_5_ XI11_4/XI0/XI0_5/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_12 XI11_4/net21_3_ xsel_5_ XI11_4/XI0/XI0_5/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_11 XI11_4/net21_4_ xsel_5_ XI11_4/XI0/XI0_5/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_10 XI11_4/net21_5_ xsel_5_ XI11_4/XI0/XI0_5/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_9 XI11_4/net21_6_ xsel_5_ XI11_4/XI0/XI0_5/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_8 XI11_4/net21_7_ xsel_5_ XI11_4/XI0/XI0_5/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_7 XI11_4/net21_8_ xsel_5_ XI11_4/XI0/XI0_5/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_6 XI11_4/net21_9_ xsel_5_ XI11_4/XI0/XI0_5/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_5 XI11_4/net21_10_ xsel_5_ XI11_4/XI0/XI0_5/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_4 XI11_4/net21_11_ xsel_5_ XI11_4/XI0/XI0_5/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_3 XI11_4/net21_12_ xsel_5_ XI11_4/XI0/XI0_5/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_2 XI11_4/net21_13_ xsel_5_ XI11_4/XI0/XI0_5/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_1 XI11_4/net21_14_ xsel_5_ XI11_4/XI0/XI0_5/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_0 XI11_4/net21_15_ xsel_5_ XI11_4/XI0/XI0_5/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_15 XI11_4/XI0/XI0_5/d__15_ xsel_5_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_14 XI11_4/XI0/XI0_5/d__14_ xsel_5_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_13 XI11_4/XI0/XI0_5/d__13_ xsel_5_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_12 XI11_4/XI0/XI0_5/d__12_ xsel_5_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_11 XI11_4/XI0/XI0_5/d__11_ xsel_5_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_10 XI11_4/XI0/XI0_5/d__10_ xsel_5_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_9 XI11_4/XI0/XI0_5/d__9_ xsel_5_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_8 XI11_4/XI0/XI0_5/d__8_ xsel_5_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_7 XI11_4/XI0/XI0_5/d__7_ xsel_5_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_6 XI11_4/XI0/XI0_5/d__6_ xsel_5_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_5 XI11_4/XI0/XI0_5/d__5_ xsel_5_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_4 XI11_4/XI0/XI0_5/d__4_ xsel_5_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_3 XI11_4/XI0/XI0_5/d__3_ xsel_5_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_2 XI11_4/XI0/XI0_5/d__2_ xsel_5_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_1 XI11_4/XI0/XI0_5/d__1_ xsel_5_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_0 XI11_4/XI0/XI0_5/d__0_ xsel_5_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_15 XI11_4/net21_0_ xsel_4_ XI11_4/XI0/XI0_4/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_14 XI11_4/net21_1_ xsel_4_ XI11_4/XI0/XI0_4/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_13 XI11_4/net21_2_ xsel_4_ XI11_4/XI0/XI0_4/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_12 XI11_4/net21_3_ xsel_4_ XI11_4/XI0/XI0_4/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_11 XI11_4/net21_4_ xsel_4_ XI11_4/XI0/XI0_4/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_10 XI11_4/net21_5_ xsel_4_ XI11_4/XI0/XI0_4/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_9 XI11_4/net21_6_ xsel_4_ XI11_4/XI0/XI0_4/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_8 XI11_4/net21_7_ xsel_4_ XI11_4/XI0/XI0_4/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_7 XI11_4/net21_8_ xsel_4_ XI11_4/XI0/XI0_4/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_6 XI11_4/net21_9_ xsel_4_ XI11_4/XI0/XI0_4/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_5 XI11_4/net21_10_ xsel_4_ XI11_4/XI0/XI0_4/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_4 XI11_4/net21_11_ xsel_4_ XI11_4/XI0/XI0_4/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_3 XI11_4/net21_12_ xsel_4_ XI11_4/XI0/XI0_4/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_2 XI11_4/net21_13_ xsel_4_ XI11_4/XI0/XI0_4/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_1 XI11_4/net21_14_ xsel_4_ XI11_4/XI0/XI0_4/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_0 XI11_4/net21_15_ xsel_4_ XI11_4/XI0/XI0_4/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_15 XI11_4/XI0/XI0_4/d__15_ xsel_4_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_14 XI11_4/XI0/XI0_4/d__14_ xsel_4_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_13 XI11_4/XI0/XI0_4/d__13_ xsel_4_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_12 XI11_4/XI0/XI0_4/d__12_ xsel_4_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_11 XI11_4/XI0/XI0_4/d__11_ xsel_4_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_10 XI11_4/XI0/XI0_4/d__10_ xsel_4_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_9 XI11_4/XI0/XI0_4/d__9_ xsel_4_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_8 XI11_4/XI0/XI0_4/d__8_ xsel_4_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_7 XI11_4/XI0/XI0_4/d__7_ xsel_4_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_6 XI11_4/XI0/XI0_4/d__6_ xsel_4_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_5 XI11_4/XI0/XI0_4/d__5_ xsel_4_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_4 XI11_4/XI0/XI0_4/d__4_ xsel_4_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_3 XI11_4/XI0/XI0_4/d__3_ xsel_4_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_2 XI11_4/XI0/XI0_4/d__2_ xsel_4_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_1 XI11_4/XI0/XI0_4/d__1_ xsel_4_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_0 XI11_4/XI0/XI0_4/d__0_ xsel_4_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_15 XI11_4/net21_0_ xsel_3_ XI11_4/XI0/XI0_3/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_14 XI11_4/net21_1_ xsel_3_ XI11_4/XI0/XI0_3/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_13 XI11_4/net21_2_ xsel_3_ XI11_4/XI0/XI0_3/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_12 XI11_4/net21_3_ xsel_3_ XI11_4/XI0/XI0_3/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_11 XI11_4/net21_4_ xsel_3_ XI11_4/XI0/XI0_3/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_10 XI11_4/net21_5_ xsel_3_ XI11_4/XI0/XI0_3/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_9 XI11_4/net21_6_ xsel_3_ XI11_4/XI0/XI0_3/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_8 XI11_4/net21_7_ xsel_3_ XI11_4/XI0/XI0_3/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_7 XI11_4/net21_8_ xsel_3_ XI11_4/XI0/XI0_3/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_6 XI11_4/net21_9_ xsel_3_ XI11_4/XI0/XI0_3/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_5 XI11_4/net21_10_ xsel_3_ XI11_4/XI0/XI0_3/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_4 XI11_4/net21_11_ xsel_3_ XI11_4/XI0/XI0_3/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_3 XI11_4/net21_12_ xsel_3_ XI11_4/XI0/XI0_3/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_2 XI11_4/net21_13_ xsel_3_ XI11_4/XI0/XI0_3/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_1 XI11_4/net21_14_ xsel_3_ XI11_4/XI0/XI0_3/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_0 XI11_4/net21_15_ xsel_3_ XI11_4/XI0/XI0_3/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_15 XI11_4/XI0/XI0_3/d__15_ xsel_3_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_14 XI11_4/XI0/XI0_3/d__14_ xsel_3_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_13 XI11_4/XI0/XI0_3/d__13_ xsel_3_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_12 XI11_4/XI0/XI0_3/d__12_ xsel_3_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_11 XI11_4/XI0/XI0_3/d__11_ xsel_3_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_10 XI11_4/XI0/XI0_3/d__10_ xsel_3_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_9 XI11_4/XI0/XI0_3/d__9_ xsel_3_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_8 XI11_4/XI0/XI0_3/d__8_ xsel_3_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_7 XI11_4/XI0/XI0_3/d__7_ xsel_3_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_6 XI11_4/XI0/XI0_3/d__6_ xsel_3_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_5 XI11_4/XI0/XI0_3/d__5_ xsel_3_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_4 XI11_4/XI0/XI0_3/d__4_ xsel_3_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_3 XI11_4/XI0/XI0_3/d__3_ xsel_3_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_2 XI11_4/XI0/XI0_3/d__2_ xsel_3_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_1 XI11_4/XI0/XI0_3/d__1_ xsel_3_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_0 XI11_4/XI0/XI0_3/d__0_ xsel_3_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_15 XI11_4/net21_0_ xsel_2_ XI11_4/XI0/XI0_2/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_14 XI11_4/net21_1_ xsel_2_ XI11_4/XI0/XI0_2/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_13 XI11_4/net21_2_ xsel_2_ XI11_4/XI0/XI0_2/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_12 XI11_4/net21_3_ xsel_2_ XI11_4/XI0/XI0_2/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_11 XI11_4/net21_4_ xsel_2_ XI11_4/XI0/XI0_2/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_10 XI11_4/net21_5_ xsel_2_ XI11_4/XI0/XI0_2/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_9 XI11_4/net21_6_ xsel_2_ XI11_4/XI0/XI0_2/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_8 XI11_4/net21_7_ xsel_2_ XI11_4/XI0/XI0_2/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_7 XI11_4/net21_8_ xsel_2_ XI11_4/XI0/XI0_2/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_6 XI11_4/net21_9_ xsel_2_ XI11_4/XI0/XI0_2/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_5 XI11_4/net21_10_ xsel_2_ XI11_4/XI0/XI0_2/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_4 XI11_4/net21_11_ xsel_2_ XI11_4/XI0/XI0_2/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_3 XI11_4/net21_12_ xsel_2_ XI11_4/XI0/XI0_2/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_2 XI11_4/net21_13_ xsel_2_ XI11_4/XI0/XI0_2/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_1 XI11_4/net21_14_ xsel_2_ XI11_4/XI0/XI0_2/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_0 XI11_4/net21_15_ xsel_2_ XI11_4/XI0/XI0_2/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_15 XI11_4/XI0/XI0_2/d__15_ xsel_2_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_14 XI11_4/XI0/XI0_2/d__14_ xsel_2_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_13 XI11_4/XI0/XI0_2/d__13_ xsel_2_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_12 XI11_4/XI0/XI0_2/d__12_ xsel_2_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_11 XI11_4/XI0/XI0_2/d__11_ xsel_2_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_10 XI11_4/XI0/XI0_2/d__10_ xsel_2_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_9 XI11_4/XI0/XI0_2/d__9_ xsel_2_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_8 XI11_4/XI0/XI0_2/d__8_ xsel_2_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_7 XI11_4/XI0/XI0_2/d__7_ xsel_2_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_6 XI11_4/XI0/XI0_2/d__6_ xsel_2_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_5 XI11_4/XI0/XI0_2/d__5_ xsel_2_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_4 XI11_4/XI0/XI0_2/d__4_ xsel_2_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_3 XI11_4/XI0/XI0_2/d__3_ xsel_2_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_2 XI11_4/XI0/XI0_2/d__2_ xsel_2_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_1 XI11_4/XI0/XI0_2/d__1_ xsel_2_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_0 XI11_4/XI0/XI0_2/d__0_ xsel_2_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_15 XI11_4/net21_0_ xsel_1_ XI11_4/XI0/XI0_1/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_14 XI11_4/net21_1_ xsel_1_ XI11_4/XI0/XI0_1/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_13 XI11_4/net21_2_ xsel_1_ XI11_4/XI0/XI0_1/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_12 XI11_4/net21_3_ xsel_1_ XI11_4/XI0/XI0_1/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_11 XI11_4/net21_4_ xsel_1_ XI11_4/XI0/XI0_1/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_10 XI11_4/net21_5_ xsel_1_ XI11_4/XI0/XI0_1/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_9 XI11_4/net21_6_ xsel_1_ XI11_4/XI0/XI0_1/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_8 XI11_4/net21_7_ xsel_1_ XI11_4/XI0/XI0_1/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_7 XI11_4/net21_8_ xsel_1_ XI11_4/XI0/XI0_1/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_6 XI11_4/net21_9_ xsel_1_ XI11_4/XI0/XI0_1/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_5 XI11_4/net21_10_ xsel_1_ XI11_4/XI0/XI0_1/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_4 XI11_4/net21_11_ xsel_1_ XI11_4/XI0/XI0_1/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_3 XI11_4/net21_12_ xsel_1_ XI11_4/XI0/XI0_1/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_2 XI11_4/net21_13_ xsel_1_ XI11_4/XI0/XI0_1/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_1 XI11_4/net21_14_ xsel_1_ XI11_4/XI0/XI0_1/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_0 XI11_4/net21_15_ xsel_1_ XI11_4/XI0/XI0_1/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_15 XI11_4/XI0/XI0_1/d__15_ xsel_1_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_14 XI11_4/XI0/XI0_1/d__14_ xsel_1_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_13 XI11_4/XI0/XI0_1/d__13_ xsel_1_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_12 XI11_4/XI0/XI0_1/d__12_ xsel_1_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_11 XI11_4/XI0/XI0_1/d__11_ xsel_1_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_10 XI11_4/XI0/XI0_1/d__10_ xsel_1_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_9 XI11_4/XI0/XI0_1/d__9_ xsel_1_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_8 XI11_4/XI0/XI0_1/d__8_ xsel_1_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_7 XI11_4/XI0/XI0_1/d__7_ xsel_1_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_6 XI11_4/XI0/XI0_1/d__6_ xsel_1_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_5 XI11_4/XI0/XI0_1/d__5_ xsel_1_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_4 XI11_4/XI0/XI0_1/d__4_ xsel_1_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_3 XI11_4/XI0/XI0_1/d__3_ xsel_1_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_2 XI11_4/XI0/XI0_1/d__2_ xsel_1_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_1 XI11_4/XI0/XI0_1/d__1_ xsel_1_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_0 XI11_4/XI0/XI0_1/d__0_ xsel_1_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_15 XI11_4/net21_0_ xsel_0_ XI11_4/XI0/XI0_0/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_14 XI11_4/net21_1_ xsel_0_ XI11_4/XI0/XI0_0/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_13 XI11_4/net21_2_ xsel_0_ XI11_4/XI0/XI0_0/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_12 XI11_4/net21_3_ xsel_0_ XI11_4/XI0/XI0_0/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_11 XI11_4/net21_4_ xsel_0_ XI11_4/XI0/XI0_0/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_10 XI11_4/net21_5_ xsel_0_ XI11_4/XI0/XI0_0/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_9 XI11_4/net21_6_ xsel_0_ XI11_4/XI0/XI0_0/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_8 XI11_4/net21_7_ xsel_0_ XI11_4/XI0/XI0_0/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_7 XI11_4/net21_8_ xsel_0_ XI11_4/XI0/XI0_0/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_6 XI11_4/net21_9_ xsel_0_ XI11_4/XI0/XI0_0/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_5 XI11_4/net21_10_ xsel_0_ XI11_4/XI0/XI0_0/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_4 XI11_4/net21_11_ xsel_0_ XI11_4/XI0/XI0_0/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_3 XI11_4/net21_12_ xsel_0_ XI11_4/XI0/XI0_0/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_2 XI11_4/net21_13_ xsel_0_ XI11_4/XI0/XI0_0/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_1 XI11_4/net21_14_ xsel_0_ XI11_4/XI0/XI0_0/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_0 XI11_4/net21_15_ xsel_0_ XI11_4/XI0/XI0_0/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_15 XI11_4/XI0/XI0_0/d__15_ xsel_0_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_14 XI11_4/XI0/XI0_0/d__14_ xsel_0_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_13 XI11_4/XI0/XI0_0/d__13_ xsel_0_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_12 XI11_4/XI0/XI0_0/d__12_ xsel_0_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_11 XI11_4/XI0/XI0_0/d__11_ xsel_0_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_10 XI11_4/XI0/XI0_0/d__10_ xsel_0_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_9 XI11_4/XI0/XI0_0/d__9_ xsel_0_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_8 XI11_4/XI0/XI0_0/d__8_ xsel_0_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_7 XI11_4/XI0/XI0_0/d__7_ xsel_0_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_6 XI11_4/XI0/XI0_0/d__6_ xsel_0_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_5 XI11_4/XI0/XI0_0/d__5_ xsel_0_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_4 XI11_4/XI0/XI0_0/d__4_ xsel_0_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_3 XI11_4/XI0/XI0_0/d__3_ xsel_0_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_2 XI11_4/XI0/XI0_0/d__2_ xsel_0_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_1 XI11_4/XI0/XI0_0/d__1_ xsel_0_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_0 XI11_4/XI0/XI0_0/d__0_ xsel_0_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI2/MN0_15 XI11_3/net21_0_ ysel_15_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_14 XI11_3/net21_1_ ysel_14_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_13 XI11_3/net21_2_ ysel_13_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_12 XI11_3/net21_3_ ysel_12_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_11 XI11_3/net21_4_ ysel_11_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_10 XI11_3/net21_5_ ysel_10_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_9 XI11_3/net21_6_ ysel_9_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_8 XI11_3/net21_7_ ysel_8_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_7 XI11_3/net21_8_ ysel_7_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_6 XI11_3/net21_9_ ysel_6_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_5 XI11_3/net21_10_ ysel_5_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_4 XI11_3/net21_11_ ysel_4_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_3 XI11_3/net21_12_ ysel_3_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_2 XI11_3/net21_13_ ysel_2_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_1 XI11_3/net21_14_ ysel_1_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_0 XI11_3/net21_15_ ysel_0_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_15 XI11_3/net20_0_ ysel_15_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_14 XI11_3/net20_1_ ysel_14_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_13 XI11_3/net20_2_ ysel_13_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_12 XI11_3/net20_3_ ysel_12_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_11 XI11_3/net20_4_ ysel_11_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_10 XI11_3/net20_5_ ysel_10_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_9 XI11_3/net20_6_ ysel_9_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_8 XI11_3/net20_7_ ysel_8_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_7 XI11_3/net20_8_ ysel_7_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_6 XI11_3/net20_9_ ysel_6_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_5 XI11_3/net20_10_ ysel_5_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_4 XI11_3/net20_11_ ysel_4_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_3 XI11_3/net20_12_ ysel_3_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_2 XI11_3/net20_13_ ysel_2_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_1 XI11_3/net20_14_ ysel_1_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_0 XI11_3/net20_15_ ysel_0_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI4/MN8 vdd XI11_3/XI4/net8 XI11_3/net12 vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_3/XI4/MP0 XI11_3/net9 XI11_3/XI4/net23 vdd vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_3/XI4/MP4 XI11_3/net12 XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI4/MP1 XI11_3/net9 XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI4/MP5 XI11_3/net12 XI11_3/preck XI11_3/net9 vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI4/MN7 vdd XI11_3/XI4/net090 DOUT_3_ vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_3/XI4/MP3 gnd XI11_3/XI4/net089 XI11_3/net12 gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_3/XI4/MN5 XI11_3/net9 XI11_3/XI4/net0103 gnd gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_3/XI4/MN4 XI11_3/XI4/data_out_ XI11_3/XI4/net32 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_3/XI4/MN0 XI11_3/XI4/data_out XI11_3/XI4/net52 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_3/XI4/MN9 gnd XI11_3/XI4/net0112 DOUT_3_ gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_3/XI1_15/MP2 XI11_3/net20_0_ XI11_3/preck XI11_3/net21_0_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_15/MP1 XI11_3/net20_0_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_15/MP0 XI11_3/net21_0_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_14/MP2 XI11_3/net20_1_ XI11_3/preck XI11_3/net21_1_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_14/MP1 XI11_3/net20_1_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_14/MP0 XI11_3/net21_1_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_13/MP2 XI11_3/net20_2_ XI11_3/preck XI11_3/net21_2_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_13/MP1 XI11_3/net20_2_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_13/MP0 XI11_3/net21_2_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_12/MP2 XI11_3/net20_3_ XI11_3/preck XI11_3/net21_3_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_12/MP1 XI11_3/net20_3_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_12/MP0 XI11_3/net21_3_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_11/MP2 XI11_3/net20_4_ XI11_3/preck XI11_3/net21_4_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_11/MP1 XI11_3/net20_4_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_11/MP0 XI11_3/net21_4_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_10/MP2 XI11_3/net20_5_ XI11_3/preck XI11_3/net21_5_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_10/MP1 XI11_3/net20_5_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_10/MP0 XI11_3/net21_5_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_9/MP2 XI11_3/net20_6_ XI11_3/preck XI11_3/net21_6_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_9/MP1 XI11_3/net20_6_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_9/MP0 XI11_3/net21_6_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_8/MP2 XI11_3/net20_7_ XI11_3/preck XI11_3/net21_7_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_8/MP1 XI11_3/net20_7_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_8/MP0 XI11_3/net21_7_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_7/MP2 XI11_3/net20_8_ XI11_3/preck XI11_3/net21_8_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_7/MP1 XI11_3/net20_8_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_7/MP0 XI11_3/net21_8_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_6/MP2 XI11_3/net20_9_ XI11_3/preck XI11_3/net21_9_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_6/MP1 XI11_3/net20_9_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_6/MP0 XI11_3/net21_9_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_5/MP2 XI11_3/net20_10_ XI11_3/preck XI11_3/net21_10_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_5/MP1 XI11_3/net20_10_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_5/MP0 XI11_3/net21_10_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_4/MP2 XI11_3/net20_11_ XI11_3/preck XI11_3/net21_11_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_4/MP1 XI11_3/net20_11_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_4/MP0 XI11_3/net21_11_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_3/MP2 XI11_3/net20_12_ XI11_3/preck XI11_3/net21_12_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_3/MP1 XI11_3/net20_12_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_3/MP0 XI11_3/net21_12_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_2/MP2 XI11_3/net20_13_ XI11_3/preck XI11_3/net21_13_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_2/MP1 XI11_3/net20_13_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_2/MP0 XI11_3/net21_13_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_1/MP2 XI11_3/net20_14_ XI11_3/preck XI11_3/net21_14_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_1/MP1 XI11_3/net20_14_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_1/MP0 XI11_3/net21_14_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_0/MP2 XI11_3/net20_15_ XI11_3/preck XI11_3/net21_15_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_0/MP1 XI11_3/net20_15_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_0/MP0 XI11_3/net21_15_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI0/MN0_15 gnd gnd XI11_3/net21_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_14 gnd gnd XI11_3/net21_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_13 gnd gnd XI11_3/net21_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_12 gnd gnd XI11_3/net21_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_11 gnd gnd XI11_3/net21_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_10 gnd gnd XI11_3/net21_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_9 gnd gnd XI11_3/net21_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_8 gnd gnd XI11_3/net21_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_7 gnd gnd XI11_3/net21_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_6 gnd gnd XI11_3/net21_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_5 gnd gnd XI11_3/net21_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_4 gnd gnd XI11_3/net21_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_3 gnd gnd XI11_3/net21_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_2 gnd gnd XI11_3/net21_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_1 gnd gnd XI11_3/net21_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_0 gnd gnd XI11_3/net21_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_15 gnd gnd XI11_3/net20_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_14 gnd gnd XI11_3/net20_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_13 gnd gnd XI11_3/net20_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_12 gnd gnd XI11_3/net20_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_11 gnd gnd XI11_3/net20_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_10 gnd gnd XI11_3/net20_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_9 gnd gnd XI11_3/net20_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_8 gnd gnd XI11_3/net20_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_7 gnd gnd XI11_3/net20_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_6 gnd gnd XI11_3/net20_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_5 gnd gnd XI11_3/net20_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_4 gnd gnd XI11_3/net20_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_3 gnd gnd XI11_3/net20_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_2 gnd gnd XI11_3/net20_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_1 gnd gnd XI11_3/net20_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_0 gnd gnd XI11_3/net20_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_15 XI11_3/net21_0_ xsel_63_ XI11_3/XI0/XI0_63/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_14 XI11_3/net21_1_ xsel_63_ XI11_3/XI0/XI0_63/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_13 XI11_3/net21_2_ xsel_63_ XI11_3/XI0/XI0_63/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_12 XI11_3/net21_3_ xsel_63_ XI11_3/XI0/XI0_63/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_11 XI11_3/net21_4_ xsel_63_ XI11_3/XI0/XI0_63/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_10 XI11_3/net21_5_ xsel_63_ XI11_3/XI0/XI0_63/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_9 XI11_3/net21_6_ xsel_63_ XI11_3/XI0/XI0_63/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_8 XI11_3/net21_7_ xsel_63_ XI11_3/XI0/XI0_63/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_7 XI11_3/net21_8_ xsel_63_ XI11_3/XI0/XI0_63/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_6 XI11_3/net21_9_ xsel_63_ XI11_3/XI0/XI0_63/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_5 XI11_3/net21_10_ xsel_63_ XI11_3/XI0/XI0_63/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_4 XI11_3/net21_11_ xsel_63_ XI11_3/XI0/XI0_63/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_3 XI11_3/net21_12_ xsel_63_ XI11_3/XI0/XI0_63/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_2 XI11_3/net21_13_ xsel_63_ XI11_3/XI0/XI0_63/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_1 XI11_3/net21_14_ xsel_63_ XI11_3/XI0/XI0_63/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_0 XI11_3/net21_15_ xsel_63_ XI11_3/XI0/XI0_63/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_15 XI11_3/XI0/XI0_63/d__15_ xsel_63_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_14 XI11_3/XI0/XI0_63/d__14_ xsel_63_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_13 XI11_3/XI0/XI0_63/d__13_ xsel_63_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_12 XI11_3/XI0/XI0_63/d__12_ xsel_63_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_11 XI11_3/XI0/XI0_63/d__11_ xsel_63_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_10 XI11_3/XI0/XI0_63/d__10_ xsel_63_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_9 XI11_3/XI0/XI0_63/d__9_ xsel_63_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_8 XI11_3/XI0/XI0_63/d__8_ xsel_63_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_7 XI11_3/XI0/XI0_63/d__7_ xsel_63_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_6 XI11_3/XI0/XI0_63/d__6_ xsel_63_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_5 XI11_3/XI0/XI0_63/d__5_ xsel_63_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_4 XI11_3/XI0/XI0_63/d__4_ xsel_63_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_3 XI11_3/XI0/XI0_63/d__3_ xsel_63_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_2 XI11_3/XI0/XI0_63/d__2_ xsel_63_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_1 XI11_3/XI0/XI0_63/d__1_ xsel_63_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_0 XI11_3/XI0/XI0_63/d__0_ xsel_63_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_15 XI11_3/net21_0_ xsel_62_ XI11_3/XI0/XI0_62/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_14 XI11_3/net21_1_ xsel_62_ XI11_3/XI0/XI0_62/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_13 XI11_3/net21_2_ xsel_62_ XI11_3/XI0/XI0_62/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_12 XI11_3/net21_3_ xsel_62_ XI11_3/XI0/XI0_62/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_11 XI11_3/net21_4_ xsel_62_ XI11_3/XI0/XI0_62/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_10 XI11_3/net21_5_ xsel_62_ XI11_3/XI0/XI0_62/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_9 XI11_3/net21_6_ xsel_62_ XI11_3/XI0/XI0_62/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_8 XI11_3/net21_7_ xsel_62_ XI11_3/XI0/XI0_62/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_7 XI11_3/net21_8_ xsel_62_ XI11_3/XI0/XI0_62/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_6 XI11_3/net21_9_ xsel_62_ XI11_3/XI0/XI0_62/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_5 XI11_3/net21_10_ xsel_62_ XI11_3/XI0/XI0_62/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_4 XI11_3/net21_11_ xsel_62_ XI11_3/XI0/XI0_62/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_3 XI11_3/net21_12_ xsel_62_ XI11_3/XI0/XI0_62/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_2 XI11_3/net21_13_ xsel_62_ XI11_3/XI0/XI0_62/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_1 XI11_3/net21_14_ xsel_62_ XI11_3/XI0/XI0_62/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_0 XI11_3/net21_15_ xsel_62_ XI11_3/XI0/XI0_62/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_15 XI11_3/XI0/XI0_62/d__15_ xsel_62_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_14 XI11_3/XI0/XI0_62/d__14_ xsel_62_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_13 XI11_3/XI0/XI0_62/d__13_ xsel_62_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_12 XI11_3/XI0/XI0_62/d__12_ xsel_62_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_11 XI11_3/XI0/XI0_62/d__11_ xsel_62_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_10 XI11_3/XI0/XI0_62/d__10_ xsel_62_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_9 XI11_3/XI0/XI0_62/d__9_ xsel_62_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_8 XI11_3/XI0/XI0_62/d__8_ xsel_62_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_7 XI11_3/XI0/XI0_62/d__7_ xsel_62_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_6 XI11_3/XI0/XI0_62/d__6_ xsel_62_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_5 XI11_3/XI0/XI0_62/d__5_ xsel_62_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_4 XI11_3/XI0/XI0_62/d__4_ xsel_62_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_3 XI11_3/XI0/XI0_62/d__3_ xsel_62_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_2 XI11_3/XI0/XI0_62/d__2_ xsel_62_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_1 XI11_3/XI0/XI0_62/d__1_ xsel_62_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_0 XI11_3/XI0/XI0_62/d__0_ xsel_62_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_15 XI11_3/net21_0_ xsel_61_ XI11_3/XI0/XI0_61/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_14 XI11_3/net21_1_ xsel_61_ XI11_3/XI0/XI0_61/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_13 XI11_3/net21_2_ xsel_61_ XI11_3/XI0/XI0_61/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_12 XI11_3/net21_3_ xsel_61_ XI11_3/XI0/XI0_61/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_11 XI11_3/net21_4_ xsel_61_ XI11_3/XI0/XI0_61/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_10 XI11_3/net21_5_ xsel_61_ XI11_3/XI0/XI0_61/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_9 XI11_3/net21_6_ xsel_61_ XI11_3/XI0/XI0_61/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_8 XI11_3/net21_7_ xsel_61_ XI11_3/XI0/XI0_61/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_7 XI11_3/net21_8_ xsel_61_ XI11_3/XI0/XI0_61/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_6 XI11_3/net21_9_ xsel_61_ XI11_3/XI0/XI0_61/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_5 XI11_3/net21_10_ xsel_61_ XI11_3/XI0/XI0_61/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_4 XI11_3/net21_11_ xsel_61_ XI11_3/XI0/XI0_61/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_3 XI11_3/net21_12_ xsel_61_ XI11_3/XI0/XI0_61/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_2 XI11_3/net21_13_ xsel_61_ XI11_3/XI0/XI0_61/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_1 XI11_3/net21_14_ xsel_61_ XI11_3/XI0/XI0_61/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_0 XI11_3/net21_15_ xsel_61_ XI11_3/XI0/XI0_61/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_15 XI11_3/XI0/XI0_61/d__15_ xsel_61_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_14 XI11_3/XI0/XI0_61/d__14_ xsel_61_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_13 XI11_3/XI0/XI0_61/d__13_ xsel_61_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_12 XI11_3/XI0/XI0_61/d__12_ xsel_61_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_11 XI11_3/XI0/XI0_61/d__11_ xsel_61_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_10 XI11_3/XI0/XI0_61/d__10_ xsel_61_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_9 XI11_3/XI0/XI0_61/d__9_ xsel_61_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_8 XI11_3/XI0/XI0_61/d__8_ xsel_61_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_7 XI11_3/XI0/XI0_61/d__7_ xsel_61_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_6 XI11_3/XI0/XI0_61/d__6_ xsel_61_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_5 XI11_3/XI0/XI0_61/d__5_ xsel_61_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_4 XI11_3/XI0/XI0_61/d__4_ xsel_61_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_3 XI11_3/XI0/XI0_61/d__3_ xsel_61_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_2 XI11_3/XI0/XI0_61/d__2_ xsel_61_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_1 XI11_3/XI0/XI0_61/d__1_ xsel_61_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_0 XI11_3/XI0/XI0_61/d__0_ xsel_61_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_15 XI11_3/net21_0_ xsel_60_ XI11_3/XI0/XI0_60/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_14 XI11_3/net21_1_ xsel_60_ XI11_3/XI0/XI0_60/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_13 XI11_3/net21_2_ xsel_60_ XI11_3/XI0/XI0_60/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_12 XI11_3/net21_3_ xsel_60_ XI11_3/XI0/XI0_60/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_11 XI11_3/net21_4_ xsel_60_ XI11_3/XI0/XI0_60/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_10 XI11_3/net21_5_ xsel_60_ XI11_3/XI0/XI0_60/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_9 XI11_3/net21_6_ xsel_60_ XI11_3/XI0/XI0_60/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_8 XI11_3/net21_7_ xsel_60_ XI11_3/XI0/XI0_60/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_7 XI11_3/net21_8_ xsel_60_ XI11_3/XI0/XI0_60/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_6 XI11_3/net21_9_ xsel_60_ XI11_3/XI0/XI0_60/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_5 XI11_3/net21_10_ xsel_60_ XI11_3/XI0/XI0_60/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_4 XI11_3/net21_11_ xsel_60_ XI11_3/XI0/XI0_60/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_3 XI11_3/net21_12_ xsel_60_ XI11_3/XI0/XI0_60/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_2 XI11_3/net21_13_ xsel_60_ XI11_3/XI0/XI0_60/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_1 XI11_3/net21_14_ xsel_60_ XI11_3/XI0/XI0_60/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_0 XI11_3/net21_15_ xsel_60_ XI11_3/XI0/XI0_60/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_15 XI11_3/XI0/XI0_60/d__15_ xsel_60_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_14 XI11_3/XI0/XI0_60/d__14_ xsel_60_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_13 XI11_3/XI0/XI0_60/d__13_ xsel_60_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_12 XI11_3/XI0/XI0_60/d__12_ xsel_60_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_11 XI11_3/XI0/XI0_60/d__11_ xsel_60_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_10 XI11_3/XI0/XI0_60/d__10_ xsel_60_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_9 XI11_3/XI0/XI0_60/d__9_ xsel_60_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_8 XI11_3/XI0/XI0_60/d__8_ xsel_60_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_7 XI11_3/XI0/XI0_60/d__7_ xsel_60_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_6 XI11_3/XI0/XI0_60/d__6_ xsel_60_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_5 XI11_3/XI0/XI0_60/d__5_ xsel_60_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_4 XI11_3/XI0/XI0_60/d__4_ xsel_60_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_3 XI11_3/XI0/XI0_60/d__3_ xsel_60_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_2 XI11_3/XI0/XI0_60/d__2_ xsel_60_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_1 XI11_3/XI0/XI0_60/d__1_ xsel_60_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_0 XI11_3/XI0/XI0_60/d__0_ xsel_60_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_15 XI11_3/net21_0_ xsel_59_ XI11_3/XI0/XI0_59/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_14 XI11_3/net21_1_ xsel_59_ XI11_3/XI0/XI0_59/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_13 XI11_3/net21_2_ xsel_59_ XI11_3/XI0/XI0_59/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_12 XI11_3/net21_3_ xsel_59_ XI11_3/XI0/XI0_59/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_11 XI11_3/net21_4_ xsel_59_ XI11_3/XI0/XI0_59/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_10 XI11_3/net21_5_ xsel_59_ XI11_3/XI0/XI0_59/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_9 XI11_3/net21_6_ xsel_59_ XI11_3/XI0/XI0_59/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_8 XI11_3/net21_7_ xsel_59_ XI11_3/XI0/XI0_59/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_7 XI11_3/net21_8_ xsel_59_ XI11_3/XI0/XI0_59/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_6 XI11_3/net21_9_ xsel_59_ XI11_3/XI0/XI0_59/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_5 XI11_3/net21_10_ xsel_59_ XI11_3/XI0/XI0_59/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_4 XI11_3/net21_11_ xsel_59_ XI11_3/XI0/XI0_59/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_3 XI11_3/net21_12_ xsel_59_ XI11_3/XI0/XI0_59/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_2 XI11_3/net21_13_ xsel_59_ XI11_3/XI0/XI0_59/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_1 XI11_3/net21_14_ xsel_59_ XI11_3/XI0/XI0_59/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_0 XI11_3/net21_15_ xsel_59_ XI11_3/XI0/XI0_59/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_15 XI11_3/XI0/XI0_59/d__15_ xsel_59_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_14 XI11_3/XI0/XI0_59/d__14_ xsel_59_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_13 XI11_3/XI0/XI0_59/d__13_ xsel_59_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_12 XI11_3/XI0/XI0_59/d__12_ xsel_59_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_11 XI11_3/XI0/XI0_59/d__11_ xsel_59_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_10 XI11_3/XI0/XI0_59/d__10_ xsel_59_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_9 XI11_3/XI0/XI0_59/d__9_ xsel_59_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_8 XI11_3/XI0/XI0_59/d__8_ xsel_59_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_7 XI11_3/XI0/XI0_59/d__7_ xsel_59_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_6 XI11_3/XI0/XI0_59/d__6_ xsel_59_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_5 XI11_3/XI0/XI0_59/d__5_ xsel_59_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_4 XI11_3/XI0/XI0_59/d__4_ xsel_59_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_3 XI11_3/XI0/XI0_59/d__3_ xsel_59_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_2 XI11_3/XI0/XI0_59/d__2_ xsel_59_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_1 XI11_3/XI0/XI0_59/d__1_ xsel_59_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_0 XI11_3/XI0/XI0_59/d__0_ xsel_59_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_15 XI11_3/net21_0_ xsel_58_ XI11_3/XI0/XI0_58/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_14 XI11_3/net21_1_ xsel_58_ XI11_3/XI0/XI0_58/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_13 XI11_3/net21_2_ xsel_58_ XI11_3/XI0/XI0_58/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_12 XI11_3/net21_3_ xsel_58_ XI11_3/XI0/XI0_58/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_11 XI11_3/net21_4_ xsel_58_ XI11_3/XI0/XI0_58/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_10 XI11_3/net21_5_ xsel_58_ XI11_3/XI0/XI0_58/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_9 XI11_3/net21_6_ xsel_58_ XI11_3/XI0/XI0_58/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_8 XI11_3/net21_7_ xsel_58_ XI11_3/XI0/XI0_58/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_7 XI11_3/net21_8_ xsel_58_ XI11_3/XI0/XI0_58/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_6 XI11_3/net21_9_ xsel_58_ XI11_3/XI0/XI0_58/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_5 XI11_3/net21_10_ xsel_58_ XI11_3/XI0/XI0_58/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_4 XI11_3/net21_11_ xsel_58_ XI11_3/XI0/XI0_58/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_3 XI11_3/net21_12_ xsel_58_ XI11_3/XI0/XI0_58/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_2 XI11_3/net21_13_ xsel_58_ XI11_3/XI0/XI0_58/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_1 XI11_3/net21_14_ xsel_58_ XI11_3/XI0/XI0_58/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_0 XI11_3/net21_15_ xsel_58_ XI11_3/XI0/XI0_58/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_15 XI11_3/XI0/XI0_58/d__15_ xsel_58_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_14 XI11_3/XI0/XI0_58/d__14_ xsel_58_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_13 XI11_3/XI0/XI0_58/d__13_ xsel_58_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_12 XI11_3/XI0/XI0_58/d__12_ xsel_58_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_11 XI11_3/XI0/XI0_58/d__11_ xsel_58_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_10 XI11_3/XI0/XI0_58/d__10_ xsel_58_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_9 XI11_3/XI0/XI0_58/d__9_ xsel_58_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_8 XI11_3/XI0/XI0_58/d__8_ xsel_58_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_7 XI11_3/XI0/XI0_58/d__7_ xsel_58_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_6 XI11_3/XI0/XI0_58/d__6_ xsel_58_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_5 XI11_3/XI0/XI0_58/d__5_ xsel_58_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_4 XI11_3/XI0/XI0_58/d__4_ xsel_58_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_3 XI11_3/XI0/XI0_58/d__3_ xsel_58_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_2 XI11_3/XI0/XI0_58/d__2_ xsel_58_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_1 XI11_3/XI0/XI0_58/d__1_ xsel_58_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_0 XI11_3/XI0/XI0_58/d__0_ xsel_58_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_15 XI11_3/net21_0_ xsel_57_ XI11_3/XI0/XI0_57/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_14 XI11_3/net21_1_ xsel_57_ XI11_3/XI0/XI0_57/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_13 XI11_3/net21_2_ xsel_57_ XI11_3/XI0/XI0_57/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_12 XI11_3/net21_3_ xsel_57_ XI11_3/XI0/XI0_57/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_11 XI11_3/net21_4_ xsel_57_ XI11_3/XI0/XI0_57/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_10 XI11_3/net21_5_ xsel_57_ XI11_3/XI0/XI0_57/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_9 XI11_3/net21_6_ xsel_57_ XI11_3/XI0/XI0_57/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_8 XI11_3/net21_7_ xsel_57_ XI11_3/XI0/XI0_57/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_7 XI11_3/net21_8_ xsel_57_ XI11_3/XI0/XI0_57/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_6 XI11_3/net21_9_ xsel_57_ XI11_3/XI0/XI0_57/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_5 XI11_3/net21_10_ xsel_57_ XI11_3/XI0/XI0_57/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_4 XI11_3/net21_11_ xsel_57_ XI11_3/XI0/XI0_57/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_3 XI11_3/net21_12_ xsel_57_ XI11_3/XI0/XI0_57/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_2 XI11_3/net21_13_ xsel_57_ XI11_3/XI0/XI0_57/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_1 XI11_3/net21_14_ xsel_57_ XI11_3/XI0/XI0_57/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_0 XI11_3/net21_15_ xsel_57_ XI11_3/XI0/XI0_57/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_15 XI11_3/XI0/XI0_57/d__15_ xsel_57_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_14 XI11_3/XI0/XI0_57/d__14_ xsel_57_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_13 XI11_3/XI0/XI0_57/d__13_ xsel_57_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_12 XI11_3/XI0/XI0_57/d__12_ xsel_57_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_11 XI11_3/XI0/XI0_57/d__11_ xsel_57_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_10 XI11_3/XI0/XI0_57/d__10_ xsel_57_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_9 XI11_3/XI0/XI0_57/d__9_ xsel_57_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_8 XI11_3/XI0/XI0_57/d__8_ xsel_57_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_7 XI11_3/XI0/XI0_57/d__7_ xsel_57_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_6 XI11_3/XI0/XI0_57/d__6_ xsel_57_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_5 XI11_3/XI0/XI0_57/d__5_ xsel_57_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_4 XI11_3/XI0/XI0_57/d__4_ xsel_57_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_3 XI11_3/XI0/XI0_57/d__3_ xsel_57_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_2 XI11_3/XI0/XI0_57/d__2_ xsel_57_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_1 XI11_3/XI0/XI0_57/d__1_ xsel_57_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_0 XI11_3/XI0/XI0_57/d__0_ xsel_57_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_15 XI11_3/net21_0_ xsel_56_ XI11_3/XI0/XI0_56/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_14 XI11_3/net21_1_ xsel_56_ XI11_3/XI0/XI0_56/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_13 XI11_3/net21_2_ xsel_56_ XI11_3/XI0/XI0_56/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_12 XI11_3/net21_3_ xsel_56_ XI11_3/XI0/XI0_56/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_11 XI11_3/net21_4_ xsel_56_ XI11_3/XI0/XI0_56/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_10 XI11_3/net21_5_ xsel_56_ XI11_3/XI0/XI0_56/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_9 XI11_3/net21_6_ xsel_56_ XI11_3/XI0/XI0_56/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_8 XI11_3/net21_7_ xsel_56_ XI11_3/XI0/XI0_56/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_7 XI11_3/net21_8_ xsel_56_ XI11_3/XI0/XI0_56/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_6 XI11_3/net21_9_ xsel_56_ XI11_3/XI0/XI0_56/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_5 XI11_3/net21_10_ xsel_56_ XI11_3/XI0/XI0_56/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_4 XI11_3/net21_11_ xsel_56_ XI11_3/XI0/XI0_56/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_3 XI11_3/net21_12_ xsel_56_ XI11_3/XI0/XI0_56/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_2 XI11_3/net21_13_ xsel_56_ XI11_3/XI0/XI0_56/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_1 XI11_3/net21_14_ xsel_56_ XI11_3/XI0/XI0_56/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_0 XI11_3/net21_15_ xsel_56_ XI11_3/XI0/XI0_56/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_15 XI11_3/XI0/XI0_56/d__15_ xsel_56_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_14 XI11_3/XI0/XI0_56/d__14_ xsel_56_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_13 XI11_3/XI0/XI0_56/d__13_ xsel_56_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_12 XI11_3/XI0/XI0_56/d__12_ xsel_56_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_11 XI11_3/XI0/XI0_56/d__11_ xsel_56_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_10 XI11_3/XI0/XI0_56/d__10_ xsel_56_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_9 XI11_3/XI0/XI0_56/d__9_ xsel_56_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_8 XI11_3/XI0/XI0_56/d__8_ xsel_56_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_7 XI11_3/XI0/XI0_56/d__7_ xsel_56_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_6 XI11_3/XI0/XI0_56/d__6_ xsel_56_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_5 XI11_3/XI0/XI0_56/d__5_ xsel_56_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_4 XI11_3/XI0/XI0_56/d__4_ xsel_56_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_3 XI11_3/XI0/XI0_56/d__3_ xsel_56_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_2 XI11_3/XI0/XI0_56/d__2_ xsel_56_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_1 XI11_3/XI0/XI0_56/d__1_ xsel_56_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_0 XI11_3/XI0/XI0_56/d__0_ xsel_56_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_15 XI11_3/net21_0_ xsel_55_ XI11_3/XI0/XI0_55/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_14 XI11_3/net21_1_ xsel_55_ XI11_3/XI0/XI0_55/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_13 XI11_3/net21_2_ xsel_55_ XI11_3/XI0/XI0_55/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_12 XI11_3/net21_3_ xsel_55_ XI11_3/XI0/XI0_55/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_11 XI11_3/net21_4_ xsel_55_ XI11_3/XI0/XI0_55/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_10 XI11_3/net21_5_ xsel_55_ XI11_3/XI0/XI0_55/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_9 XI11_3/net21_6_ xsel_55_ XI11_3/XI0/XI0_55/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_8 XI11_3/net21_7_ xsel_55_ XI11_3/XI0/XI0_55/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_7 XI11_3/net21_8_ xsel_55_ XI11_3/XI0/XI0_55/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_6 XI11_3/net21_9_ xsel_55_ XI11_3/XI0/XI0_55/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_5 XI11_3/net21_10_ xsel_55_ XI11_3/XI0/XI0_55/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_4 XI11_3/net21_11_ xsel_55_ XI11_3/XI0/XI0_55/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_3 XI11_3/net21_12_ xsel_55_ XI11_3/XI0/XI0_55/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_2 XI11_3/net21_13_ xsel_55_ XI11_3/XI0/XI0_55/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_1 XI11_3/net21_14_ xsel_55_ XI11_3/XI0/XI0_55/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_0 XI11_3/net21_15_ xsel_55_ XI11_3/XI0/XI0_55/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_15 XI11_3/XI0/XI0_55/d__15_ xsel_55_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_14 XI11_3/XI0/XI0_55/d__14_ xsel_55_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_13 XI11_3/XI0/XI0_55/d__13_ xsel_55_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_12 XI11_3/XI0/XI0_55/d__12_ xsel_55_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_11 XI11_3/XI0/XI0_55/d__11_ xsel_55_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_10 XI11_3/XI0/XI0_55/d__10_ xsel_55_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_9 XI11_3/XI0/XI0_55/d__9_ xsel_55_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_8 XI11_3/XI0/XI0_55/d__8_ xsel_55_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_7 XI11_3/XI0/XI0_55/d__7_ xsel_55_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_6 XI11_3/XI0/XI0_55/d__6_ xsel_55_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_5 XI11_3/XI0/XI0_55/d__5_ xsel_55_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_4 XI11_3/XI0/XI0_55/d__4_ xsel_55_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_3 XI11_3/XI0/XI0_55/d__3_ xsel_55_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_2 XI11_3/XI0/XI0_55/d__2_ xsel_55_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_1 XI11_3/XI0/XI0_55/d__1_ xsel_55_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_0 XI11_3/XI0/XI0_55/d__0_ xsel_55_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_15 XI11_3/net21_0_ xsel_54_ XI11_3/XI0/XI0_54/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_14 XI11_3/net21_1_ xsel_54_ XI11_3/XI0/XI0_54/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_13 XI11_3/net21_2_ xsel_54_ XI11_3/XI0/XI0_54/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_12 XI11_3/net21_3_ xsel_54_ XI11_3/XI0/XI0_54/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_11 XI11_3/net21_4_ xsel_54_ XI11_3/XI0/XI0_54/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_10 XI11_3/net21_5_ xsel_54_ XI11_3/XI0/XI0_54/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_9 XI11_3/net21_6_ xsel_54_ XI11_3/XI0/XI0_54/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_8 XI11_3/net21_7_ xsel_54_ XI11_3/XI0/XI0_54/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_7 XI11_3/net21_8_ xsel_54_ XI11_3/XI0/XI0_54/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_6 XI11_3/net21_9_ xsel_54_ XI11_3/XI0/XI0_54/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_5 XI11_3/net21_10_ xsel_54_ XI11_3/XI0/XI0_54/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_4 XI11_3/net21_11_ xsel_54_ XI11_3/XI0/XI0_54/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_3 XI11_3/net21_12_ xsel_54_ XI11_3/XI0/XI0_54/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_2 XI11_3/net21_13_ xsel_54_ XI11_3/XI0/XI0_54/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_1 XI11_3/net21_14_ xsel_54_ XI11_3/XI0/XI0_54/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_0 XI11_3/net21_15_ xsel_54_ XI11_3/XI0/XI0_54/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_15 XI11_3/XI0/XI0_54/d__15_ xsel_54_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_14 XI11_3/XI0/XI0_54/d__14_ xsel_54_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_13 XI11_3/XI0/XI0_54/d__13_ xsel_54_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_12 XI11_3/XI0/XI0_54/d__12_ xsel_54_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_11 XI11_3/XI0/XI0_54/d__11_ xsel_54_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_10 XI11_3/XI0/XI0_54/d__10_ xsel_54_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_9 XI11_3/XI0/XI0_54/d__9_ xsel_54_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_8 XI11_3/XI0/XI0_54/d__8_ xsel_54_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_7 XI11_3/XI0/XI0_54/d__7_ xsel_54_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_6 XI11_3/XI0/XI0_54/d__6_ xsel_54_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_5 XI11_3/XI0/XI0_54/d__5_ xsel_54_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_4 XI11_3/XI0/XI0_54/d__4_ xsel_54_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_3 XI11_3/XI0/XI0_54/d__3_ xsel_54_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_2 XI11_3/XI0/XI0_54/d__2_ xsel_54_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_1 XI11_3/XI0/XI0_54/d__1_ xsel_54_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_0 XI11_3/XI0/XI0_54/d__0_ xsel_54_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_15 XI11_3/net21_0_ xsel_53_ XI11_3/XI0/XI0_53/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_14 XI11_3/net21_1_ xsel_53_ XI11_3/XI0/XI0_53/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_13 XI11_3/net21_2_ xsel_53_ XI11_3/XI0/XI0_53/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_12 XI11_3/net21_3_ xsel_53_ XI11_3/XI0/XI0_53/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_11 XI11_3/net21_4_ xsel_53_ XI11_3/XI0/XI0_53/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_10 XI11_3/net21_5_ xsel_53_ XI11_3/XI0/XI0_53/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_9 XI11_3/net21_6_ xsel_53_ XI11_3/XI0/XI0_53/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_8 XI11_3/net21_7_ xsel_53_ XI11_3/XI0/XI0_53/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_7 XI11_3/net21_8_ xsel_53_ XI11_3/XI0/XI0_53/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_6 XI11_3/net21_9_ xsel_53_ XI11_3/XI0/XI0_53/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_5 XI11_3/net21_10_ xsel_53_ XI11_3/XI0/XI0_53/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_4 XI11_3/net21_11_ xsel_53_ XI11_3/XI0/XI0_53/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_3 XI11_3/net21_12_ xsel_53_ XI11_3/XI0/XI0_53/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_2 XI11_3/net21_13_ xsel_53_ XI11_3/XI0/XI0_53/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_1 XI11_3/net21_14_ xsel_53_ XI11_3/XI0/XI0_53/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_0 XI11_3/net21_15_ xsel_53_ XI11_3/XI0/XI0_53/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_15 XI11_3/XI0/XI0_53/d__15_ xsel_53_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_14 XI11_3/XI0/XI0_53/d__14_ xsel_53_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_13 XI11_3/XI0/XI0_53/d__13_ xsel_53_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_12 XI11_3/XI0/XI0_53/d__12_ xsel_53_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_11 XI11_3/XI0/XI0_53/d__11_ xsel_53_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_10 XI11_3/XI0/XI0_53/d__10_ xsel_53_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_9 XI11_3/XI0/XI0_53/d__9_ xsel_53_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_8 XI11_3/XI0/XI0_53/d__8_ xsel_53_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_7 XI11_3/XI0/XI0_53/d__7_ xsel_53_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_6 XI11_3/XI0/XI0_53/d__6_ xsel_53_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_5 XI11_3/XI0/XI0_53/d__5_ xsel_53_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_4 XI11_3/XI0/XI0_53/d__4_ xsel_53_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_3 XI11_3/XI0/XI0_53/d__3_ xsel_53_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_2 XI11_3/XI0/XI0_53/d__2_ xsel_53_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_1 XI11_3/XI0/XI0_53/d__1_ xsel_53_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_0 XI11_3/XI0/XI0_53/d__0_ xsel_53_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_15 XI11_3/net21_0_ xsel_52_ XI11_3/XI0/XI0_52/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_14 XI11_3/net21_1_ xsel_52_ XI11_3/XI0/XI0_52/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_13 XI11_3/net21_2_ xsel_52_ XI11_3/XI0/XI0_52/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_12 XI11_3/net21_3_ xsel_52_ XI11_3/XI0/XI0_52/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_11 XI11_3/net21_4_ xsel_52_ XI11_3/XI0/XI0_52/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_10 XI11_3/net21_5_ xsel_52_ XI11_3/XI0/XI0_52/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_9 XI11_3/net21_6_ xsel_52_ XI11_3/XI0/XI0_52/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_8 XI11_3/net21_7_ xsel_52_ XI11_3/XI0/XI0_52/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_7 XI11_3/net21_8_ xsel_52_ XI11_3/XI0/XI0_52/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_6 XI11_3/net21_9_ xsel_52_ XI11_3/XI0/XI0_52/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_5 XI11_3/net21_10_ xsel_52_ XI11_3/XI0/XI0_52/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_4 XI11_3/net21_11_ xsel_52_ XI11_3/XI0/XI0_52/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_3 XI11_3/net21_12_ xsel_52_ XI11_3/XI0/XI0_52/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_2 XI11_3/net21_13_ xsel_52_ XI11_3/XI0/XI0_52/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_1 XI11_3/net21_14_ xsel_52_ XI11_3/XI0/XI0_52/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_0 XI11_3/net21_15_ xsel_52_ XI11_3/XI0/XI0_52/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_15 XI11_3/XI0/XI0_52/d__15_ xsel_52_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_14 XI11_3/XI0/XI0_52/d__14_ xsel_52_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_13 XI11_3/XI0/XI0_52/d__13_ xsel_52_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_12 XI11_3/XI0/XI0_52/d__12_ xsel_52_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_11 XI11_3/XI0/XI0_52/d__11_ xsel_52_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_10 XI11_3/XI0/XI0_52/d__10_ xsel_52_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_9 XI11_3/XI0/XI0_52/d__9_ xsel_52_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_8 XI11_3/XI0/XI0_52/d__8_ xsel_52_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_7 XI11_3/XI0/XI0_52/d__7_ xsel_52_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_6 XI11_3/XI0/XI0_52/d__6_ xsel_52_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_5 XI11_3/XI0/XI0_52/d__5_ xsel_52_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_4 XI11_3/XI0/XI0_52/d__4_ xsel_52_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_3 XI11_3/XI0/XI0_52/d__3_ xsel_52_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_2 XI11_3/XI0/XI0_52/d__2_ xsel_52_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_1 XI11_3/XI0/XI0_52/d__1_ xsel_52_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_0 XI11_3/XI0/XI0_52/d__0_ xsel_52_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_15 XI11_3/net21_0_ xsel_51_ XI11_3/XI0/XI0_51/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_14 XI11_3/net21_1_ xsel_51_ XI11_3/XI0/XI0_51/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_13 XI11_3/net21_2_ xsel_51_ XI11_3/XI0/XI0_51/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_12 XI11_3/net21_3_ xsel_51_ XI11_3/XI0/XI0_51/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_11 XI11_3/net21_4_ xsel_51_ XI11_3/XI0/XI0_51/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_10 XI11_3/net21_5_ xsel_51_ XI11_3/XI0/XI0_51/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_9 XI11_3/net21_6_ xsel_51_ XI11_3/XI0/XI0_51/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_8 XI11_3/net21_7_ xsel_51_ XI11_3/XI0/XI0_51/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_7 XI11_3/net21_8_ xsel_51_ XI11_3/XI0/XI0_51/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_6 XI11_3/net21_9_ xsel_51_ XI11_3/XI0/XI0_51/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_5 XI11_3/net21_10_ xsel_51_ XI11_3/XI0/XI0_51/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_4 XI11_3/net21_11_ xsel_51_ XI11_3/XI0/XI0_51/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_3 XI11_3/net21_12_ xsel_51_ XI11_3/XI0/XI0_51/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_2 XI11_3/net21_13_ xsel_51_ XI11_3/XI0/XI0_51/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_1 XI11_3/net21_14_ xsel_51_ XI11_3/XI0/XI0_51/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_0 XI11_3/net21_15_ xsel_51_ XI11_3/XI0/XI0_51/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_15 XI11_3/XI0/XI0_51/d__15_ xsel_51_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_14 XI11_3/XI0/XI0_51/d__14_ xsel_51_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_13 XI11_3/XI0/XI0_51/d__13_ xsel_51_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_12 XI11_3/XI0/XI0_51/d__12_ xsel_51_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_11 XI11_3/XI0/XI0_51/d__11_ xsel_51_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_10 XI11_3/XI0/XI0_51/d__10_ xsel_51_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_9 XI11_3/XI0/XI0_51/d__9_ xsel_51_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_8 XI11_3/XI0/XI0_51/d__8_ xsel_51_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_7 XI11_3/XI0/XI0_51/d__7_ xsel_51_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_6 XI11_3/XI0/XI0_51/d__6_ xsel_51_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_5 XI11_3/XI0/XI0_51/d__5_ xsel_51_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_4 XI11_3/XI0/XI0_51/d__4_ xsel_51_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_3 XI11_3/XI0/XI0_51/d__3_ xsel_51_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_2 XI11_3/XI0/XI0_51/d__2_ xsel_51_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_1 XI11_3/XI0/XI0_51/d__1_ xsel_51_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_0 XI11_3/XI0/XI0_51/d__0_ xsel_51_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_15 XI11_3/net21_0_ xsel_50_ XI11_3/XI0/XI0_50/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_14 XI11_3/net21_1_ xsel_50_ XI11_3/XI0/XI0_50/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_13 XI11_3/net21_2_ xsel_50_ XI11_3/XI0/XI0_50/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_12 XI11_3/net21_3_ xsel_50_ XI11_3/XI0/XI0_50/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_11 XI11_3/net21_4_ xsel_50_ XI11_3/XI0/XI0_50/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_10 XI11_3/net21_5_ xsel_50_ XI11_3/XI0/XI0_50/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_9 XI11_3/net21_6_ xsel_50_ XI11_3/XI0/XI0_50/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_8 XI11_3/net21_7_ xsel_50_ XI11_3/XI0/XI0_50/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_7 XI11_3/net21_8_ xsel_50_ XI11_3/XI0/XI0_50/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_6 XI11_3/net21_9_ xsel_50_ XI11_3/XI0/XI0_50/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_5 XI11_3/net21_10_ xsel_50_ XI11_3/XI0/XI0_50/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_4 XI11_3/net21_11_ xsel_50_ XI11_3/XI0/XI0_50/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_3 XI11_3/net21_12_ xsel_50_ XI11_3/XI0/XI0_50/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_2 XI11_3/net21_13_ xsel_50_ XI11_3/XI0/XI0_50/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_1 XI11_3/net21_14_ xsel_50_ XI11_3/XI0/XI0_50/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_0 XI11_3/net21_15_ xsel_50_ XI11_3/XI0/XI0_50/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_15 XI11_3/XI0/XI0_50/d__15_ xsel_50_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_14 XI11_3/XI0/XI0_50/d__14_ xsel_50_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_13 XI11_3/XI0/XI0_50/d__13_ xsel_50_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_12 XI11_3/XI0/XI0_50/d__12_ xsel_50_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_11 XI11_3/XI0/XI0_50/d__11_ xsel_50_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_10 XI11_3/XI0/XI0_50/d__10_ xsel_50_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_9 XI11_3/XI0/XI0_50/d__9_ xsel_50_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_8 XI11_3/XI0/XI0_50/d__8_ xsel_50_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_7 XI11_3/XI0/XI0_50/d__7_ xsel_50_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_6 XI11_3/XI0/XI0_50/d__6_ xsel_50_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_5 XI11_3/XI0/XI0_50/d__5_ xsel_50_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_4 XI11_3/XI0/XI0_50/d__4_ xsel_50_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_3 XI11_3/XI0/XI0_50/d__3_ xsel_50_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_2 XI11_3/XI0/XI0_50/d__2_ xsel_50_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_1 XI11_3/XI0/XI0_50/d__1_ xsel_50_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_0 XI11_3/XI0/XI0_50/d__0_ xsel_50_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_15 XI11_3/net21_0_ xsel_49_ XI11_3/XI0/XI0_49/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_14 XI11_3/net21_1_ xsel_49_ XI11_3/XI0/XI0_49/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_13 XI11_3/net21_2_ xsel_49_ XI11_3/XI0/XI0_49/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_12 XI11_3/net21_3_ xsel_49_ XI11_3/XI0/XI0_49/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_11 XI11_3/net21_4_ xsel_49_ XI11_3/XI0/XI0_49/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_10 XI11_3/net21_5_ xsel_49_ XI11_3/XI0/XI0_49/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_9 XI11_3/net21_6_ xsel_49_ XI11_3/XI0/XI0_49/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_8 XI11_3/net21_7_ xsel_49_ XI11_3/XI0/XI0_49/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_7 XI11_3/net21_8_ xsel_49_ XI11_3/XI0/XI0_49/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_6 XI11_3/net21_9_ xsel_49_ XI11_3/XI0/XI0_49/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_5 XI11_3/net21_10_ xsel_49_ XI11_3/XI0/XI0_49/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_4 XI11_3/net21_11_ xsel_49_ XI11_3/XI0/XI0_49/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_3 XI11_3/net21_12_ xsel_49_ XI11_3/XI0/XI0_49/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_2 XI11_3/net21_13_ xsel_49_ XI11_3/XI0/XI0_49/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_1 XI11_3/net21_14_ xsel_49_ XI11_3/XI0/XI0_49/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_0 XI11_3/net21_15_ xsel_49_ XI11_3/XI0/XI0_49/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_15 XI11_3/XI0/XI0_49/d__15_ xsel_49_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_14 XI11_3/XI0/XI0_49/d__14_ xsel_49_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_13 XI11_3/XI0/XI0_49/d__13_ xsel_49_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_12 XI11_3/XI0/XI0_49/d__12_ xsel_49_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_11 XI11_3/XI0/XI0_49/d__11_ xsel_49_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_10 XI11_3/XI0/XI0_49/d__10_ xsel_49_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_9 XI11_3/XI0/XI0_49/d__9_ xsel_49_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_8 XI11_3/XI0/XI0_49/d__8_ xsel_49_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_7 XI11_3/XI0/XI0_49/d__7_ xsel_49_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_6 XI11_3/XI0/XI0_49/d__6_ xsel_49_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_5 XI11_3/XI0/XI0_49/d__5_ xsel_49_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_4 XI11_3/XI0/XI0_49/d__4_ xsel_49_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_3 XI11_3/XI0/XI0_49/d__3_ xsel_49_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_2 XI11_3/XI0/XI0_49/d__2_ xsel_49_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_1 XI11_3/XI0/XI0_49/d__1_ xsel_49_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_0 XI11_3/XI0/XI0_49/d__0_ xsel_49_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_15 XI11_3/net21_0_ xsel_48_ XI11_3/XI0/XI0_48/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_14 XI11_3/net21_1_ xsel_48_ XI11_3/XI0/XI0_48/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_13 XI11_3/net21_2_ xsel_48_ XI11_3/XI0/XI0_48/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_12 XI11_3/net21_3_ xsel_48_ XI11_3/XI0/XI0_48/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_11 XI11_3/net21_4_ xsel_48_ XI11_3/XI0/XI0_48/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_10 XI11_3/net21_5_ xsel_48_ XI11_3/XI0/XI0_48/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_9 XI11_3/net21_6_ xsel_48_ XI11_3/XI0/XI0_48/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_8 XI11_3/net21_7_ xsel_48_ XI11_3/XI0/XI0_48/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_7 XI11_3/net21_8_ xsel_48_ XI11_3/XI0/XI0_48/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_6 XI11_3/net21_9_ xsel_48_ XI11_3/XI0/XI0_48/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_5 XI11_3/net21_10_ xsel_48_ XI11_3/XI0/XI0_48/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_4 XI11_3/net21_11_ xsel_48_ XI11_3/XI0/XI0_48/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_3 XI11_3/net21_12_ xsel_48_ XI11_3/XI0/XI0_48/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_2 XI11_3/net21_13_ xsel_48_ XI11_3/XI0/XI0_48/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_1 XI11_3/net21_14_ xsel_48_ XI11_3/XI0/XI0_48/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_0 XI11_3/net21_15_ xsel_48_ XI11_3/XI0/XI0_48/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_15 XI11_3/XI0/XI0_48/d__15_ xsel_48_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_14 XI11_3/XI0/XI0_48/d__14_ xsel_48_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_13 XI11_3/XI0/XI0_48/d__13_ xsel_48_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_12 XI11_3/XI0/XI0_48/d__12_ xsel_48_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_11 XI11_3/XI0/XI0_48/d__11_ xsel_48_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_10 XI11_3/XI0/XI0_48/d__10_ xsel_48_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_9 XI11_3/XI0/XI0_48/d__9_ xsel_48_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_8 XI11_3/XI0/XI0_48/d__8_ xsel_48_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_7 XI11_3/XI0/XI0_48/d__7_ xsel_48_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_6 XI11_3/XI0/XI0_48/d__6_ xsel_48_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_5 XI11_3/XI0/XI0_48/d__5_ xsel_48_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_4 XI11_3/XI0/XI0_48/d__4_ xsel_48_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_3 XI11_3/XI0/XI0_48/d__3_ xsel_48_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_2 XI11_3/XI0/XI0_48/d__2_ xsel_48_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_1 XI11_3/XI0/XI0_48/d__1_ xsel_48_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_0 XI11_3/XI0/XI0_48/d__0_ xsel_48_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_15 XI11_3/net21_0_ xsel_47_ XI11_3/XI0/XI0_47/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_14 XI11_3/net21_1_ xsel_47_ XI11_3/XI0/XI0_47/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_13 XI11_3/net21_2_ xsel_47_ XI11_3/XI0/XI0_47/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_12 XI11_3/net21_3_ xsel_47_ XI11_3/XI0/XI0_47/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_11 XI11_3/net21_4_ xsel_47_ XI11_3/XI0/XI0_47/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_10 XI11_3/net21_5_ xsel_47_ XI11_3/XI0/XI0_47/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_9 XI11_3/net21_6_ xsel_47_ XI11_3/XI0/XI0_47/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_8 XI11_3/net21_7_ xsel_47_ XI11_3/XI0/XI0_47/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_7 XI11_3/net21_8_ xsel_47_ XI11_3/XI0/XI0_47/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_6 XI11_3/net21_9_ xsel_47_ XI11_3/XI0/XI0_47/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_5 XI11_3/net21_10_ xsel_47_ XI11_3/XI0/XI0_47/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_4 XI11_3/net21_11_ xsel_47_ XI11_3/XI0/XI0_47/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_3 XI11_3/net21_12_ xsel_47_ XI11_3/XI0/XI0_47/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_2 XI11_3/net21_13_ xsel_47_ XI11_3/XI0/XI0_47/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_1 XI11_3/net21_14_ xsel_47_ XI11_3/XI0/XI0_47/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_0 XI11_3/net21_15_ xsel_47_ XI11_3/XI0/XI0_47/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_15 XI11_3/XI0/XI0_47/d__15_ xsel_47_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_14 XI11_3/XI0/XI0_47/d__14_ xsel_47_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_13 XI11_3/XI0/XI0_47/d__13_ xsel_47_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_12 XI11_3/XI0/XI0_47/d__12_ xsel_47_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_11 XI11_3/XI0/XI0_47/d__11_ xsel_47_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_10 XI11_3/XI0/XI0_47/d__10_ xsel_47_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_9 XI11_3/XI0/XI0_47/d__9_ xsel_47_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_8 XI11_3/XI0/XI0_47/d__8_ xsel_47_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_7 XI11_3/XI0/XI0_47/d__7_ xsel_47_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_6 XI11_3/XI0/XI0_47/d__6_ xsel_47_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_5 XI11_3/XI0/XI0_47/d__5_ xsel_47_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_4 XI11_3/XI0/XI0_47/d__4_ xsel_47_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_3 XI11_3/XI0/XI0_47/d__3_ xsel_47_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_2 XI11_3/XI0/XI0_47/d__2_ xsel_47_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_1 XI11_3/XI0/XI0_47/d__1_ xsel_47_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_0 XI11_3/XI0/XI0_47/d__0_ xsel_47_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_15 XI11_3/net21_0_ xsel_46_ XI11_3/XI0/XI0_46/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_14 XI11_3/net21_1_ xsel_46_ XI11_3/XI0/XI0_46/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_13 XI11_3/net21_2_ xsel_46_ XI11_3/XI0/XI0_46/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_12 XI11_3/net21_3_ xsel_46_ XI11_3/XI0/XI0_46/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_11 XI11_3/net21_4_ xsel_46_ XI11_3/XI0/XI0_46/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_10 XI11_3/net21_5_ xsel_46_ XI11_3/XI0/XI0_46/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_9 XI11_3/net21_6_ xsel_46_ XI11_3/XI0/XI0_46/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_8 XI11_3/net21_7_ xsel_46_ XI11_3/XI0/XI0_46/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_7 XI11_3/net21_8_ xsel_46_ XI11_3/XI0/XI0_46/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_6 XI11_3/net21_9_ xsel_46_ XI11_3/XI0/XI0_46/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_5 XI11_3/net21_10_ xsel_46_ XI11_3/XI0/XI0_46/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_4 XI11_3/net21_11_ xsel_46_ XI11_3/XI0/XI0_46/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_3 XI11_3/net21_12_ xsel_46_ XI11_3/XI0/XI0_46/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_2 XI11_3/net21_13_ xsel_46_ XI11_3/XI0/XI0_46/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_1 XI11_3/net21_14_ xsel_46_ XI11_3/XI0/XI0_46/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_0 XI11_3/net21_15_ xsel_46_ XI11_3/XI0/XI0_46/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_15 XI11_3/XI0/XI0_46/d__15_ xsel_46_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_14 XI11_3/XI0/XI0_46/d__14_ xsel_46_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_13 XI11_3/XI0/XI0_46/d__13_ xsel_46_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_12 XI11_3/XI0/XI0_46/d__12_ xsel_46_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_11 XI11_3/XI0/XI0_46/d__11_ xsel_46_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_10 XI11_3/XI0/XI0_46/d__10_ xsel_46_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_9 XI11_3/XI0/XI0_46/d__9_ xsel_46_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_8 XI11_3/XI0/XI0_46/d__8_ xsel_46_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_7 XI11_3/XI0/XI0_46/d__7_ xsel_46_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_6 XI11_3/XI0/XI0_46/d__6_ xsel_46_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_5 XI11_3/XI0/XI0_46/d__5_ xsel_46_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_4 XI11_3/XI0/XI0_46/d__4_ xsel_46_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_3 XI11_3/XI0/XI0_46/d__3_ xsel_46_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_2 XI11_3/XI0/XI0_46/d__2_ xsel_46_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_1 XI11_3/XI0/XI0_46/d__1_ xsel_46_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_0 XI11_3/XI0/XI0_46/d__0_ xsel_46_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_15 XI11_3/net21_0_ xsel_45_ XI11_3/XI0/XI0_45/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_14 XI11_3/net21_1_ xsel_45_ XI11_3/XI0/XI0_45/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_13 XI11_3/net21_2_ xsel_45_ XI11_3/XI0/XI0_45/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_12 XI11_3/net21_3_ xsel_45_ XI11_3/XI0/XI0_45/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_11 XI11_3/net21_4_ xsel_45_ XI11_3/XI0/XI0_45/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_10 XI11_3/net21_5_ xsel_45_ XI11_3/XI0/XI0_45/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_9 XI11_3/net21_6_ xsel_45_ XI11_3/XI0/XI0_45/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_8 XI11_3/net21_7_ xsel_45_ XI11_3/XI0/XI0_45/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_7 XI11_3/net21_8_ xsel_45_ XI11_3/XI0/XI0_45/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_6 XI11_3/net21_9_ xsel_45_ XI11_3/XI0/XI0_45/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_5 XI11_3/net21_10_ xsel_45_ XI11_3/XI0/XI0_45/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_4 XI11_3/net21_11_ xsel_45_ XI11_3/XI0/XI0_45/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_3 XI11_3/net21_12_ xsel_45_ XI11_3/XI0/XI0_45/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_2 XI11_3/net21_13_ xsel_45_ XI11_3/XI0/XI0_45/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_1 XI11_3/net21_14_ xsel_45_ XI11_3/XI0/XI0_45/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_0 XI11_3/net21_15_ xsel_45_ XI11_3/XI0/XI0_45/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_15 XI11_3/XI0/XI0_45/d__15_ xsel_45_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_14 XI11_3/XI0/XI0_45/d__14_ xsel_45_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_13 XI11_3/XI0/XI0_45/d__13_ xsel_45_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_12 XI11_3/XI0/XI0_45/d__12_ xsel_45_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_11 XI11_3/XI0/XI0_45/d__11_ xsel_45_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_10 XI11_3/XI0/XI0_45/d__10_ xsel_45_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_9 XI11_3/XI0/XI0_45/d__9_ xsel_45_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_8 XI11_3/XI0/XI0_45/d__8_ xsel_45_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_7 XI11_3/XI0/XI0_45/d__7_ xsel_45_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_6 XI11_3/XI0/XI0_45/d__6_ xsel_45_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_5 XI11_3/XI0/XI0_45/d__5_ xsel_45_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_4 XI11_3/XI0/XI0_45/d__4_ xsel_45_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_3 XI11_3/XI0/XI0_45/d__3_ xsel_45_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_2 XI11_3/XI0/XI0_45/d__2_ xsel_45_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_1 XI11_3/XI0/XI0_45/d__1_ xsel_45_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_0 XI11_3/XI0/XI0_45/d__0_ xsel_45_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_15 XI11_3/net21_0_ xsel_44_ XI11_3/XI0/XI0_44/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_14 XI11_3/net21_1_ xsel_44_ XI11_3/XI0/XI0_44/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_13 XI11_3/net21_2_ xsel_44_ XI11_3/XI0/XI0_44/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_12 XI11_3/net21_3_ xsel_44_ XI11_3/XI0/XI0_44/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_11 XI11_3/net21_4_ xsel_44_ XI11_3/XI0/XI0_44/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_10 XI11_3/net21_5_ xsel_44_ XI11_3/XI0/XI0_44/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_9 XI11_3/net21_6_ xsel_44_ XI11_3/XI0/XI0_44/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_8 XI11_3/net21_7_ xsel_44_ XI11_3/XI0/XI0_44/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_7 XI11_3/net21_8_ xsel_44_ XI11_3/XI0/XI0_44/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_6 XI11_3/net21_9_ xsel_44_ XI11_3/XI0/XI0_44/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_5 XI11_3/net21_10_ xsel_44_ XI11_3/XI0/XI0_44/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_4 XI11_3/net21_11_ xsel_44_ XI11_3/XI0/XI0_44/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_3 XI11_3/net21_12_ xsel_44_ XI11_3/XI0/XI0_44/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_2 XI11_3/net21_13_ xsel_44_ XI11_3/XI0/XI0_44/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_1 XI11_3/net21_14_ xsel_44_ XI11_3/XI0/XI0_44/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_0 XI11_3/net21_15_ xsel_44_ XI11_3/XI0/XI0_44/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_15 XI11_3/XI0/XI0_44/d__15_ xsel_44_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_14 XI11_3/XI0/XI0_44/d__14_ xsel_44_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_13 XI11_3/XI0/XI0_44/d__13_ xsel_44_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_12 XI11_3/XI0/XI0_44/d__12_ xsel_44_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_11 XI11_3/XI0/XI0_44/d__11_ xsel_44_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_10 XI11_3/XI0/XI0_44/d__10_ xsel_44_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_9 XI11_3/XI0/XI0_44/d__9_ xsel_44_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_8 XI11_3/XI0/XI0_44/d__8_ xsel_44_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_7 XI11_3/XI0/XI0_44/d__7_ xsel_44_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_6 XI11_3/XI0/XI0_44/d__6_ xsel_44_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_5 XI11_3/XI0/XI0_44/d__5_ xsel_44_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_4 XI11_3/XI0/XI0_44/d__4_ xsel_44_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_3 XI11_3/XI0/XI0_44/d__3_ xsel_44_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_2 XI11_3/XI0/XI0_44/d__2_ xsel_44_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_1 XI11_3/XI0/XI0_44/d__1_ xsel_44_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_0 XI11_3/XI0/XI0_44/d__0_ xsel_44_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_15 XI11_3/net21_0_ xsel_43_ XI11_3/XI0/XI0_43/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_14 XI11_3/net21_1_ xsel_43_ XI11_3/XI0/XI0_43/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_13 XI11_3/net21_2_ xsel_43_ XI11_3/XI0/XI0_43/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_12 XI11_3/net21_3_ xsel_43_ XI11_3/XI0/XI0_43/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_11 XI11_3/net21_4_ xsel_43_ XI11_3/XI0/XI0_43/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_10 XI11_3/net21_5_ xsel_43_ XI11_3/XI0/XI0_43/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_9 XI11_3/net21_6_ xsel_43_ XI11_3/XI0/XI0_43/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_8 XI11_3/net21_7_ xsel_43_ XI11_3/XI0/XI0_43/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_7 XI11_3/net21_8_ xsel_43_ XI11_3/XI0/XI0_43/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_6 XI11_3/net21_9_ xsel_43_ XI11_3/XI0/XI0_43/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_5 XI11_3/net21_10_ xsel_43_ XI11_3/XI0/XI0_43/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_4 XI11_3/net21_11_ xsel_43_ XI11_3/XI0/XI0_43/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_3 XI11_3/net21_12_ xsel_43_ XI11_3/XI0/XI0_43/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_2 XI11_3/net21_13_ xsel_43_ XI11_3/XI0/XI0_43/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_1 XI11_3/net21_14_ xsel_43_ XI11_3/XI0/XI0_43/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_0 XI11_3/net21_15_ xsel_43_ XI11_3/XI0/XI0_43/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_15 XI11_3/XI0/XI0_43/d__15_ xsel_43_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_14 XI11_3/XI0/XI0_43/d__14_ xsel_43_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_13 XI11_3/XI0/XI0_43/d__13_ xsel_43_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_12 XI11_3/XI0/XI0_43/d__12_ xsel_43_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_11 XI11_3/XI0/XI0_43/d__11_ xsel_43_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_10 XI11_3/XI0/XI0_43/d__10_ xsel_43_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_9 XI11_3/XI0/XI0_43/d__9_ xsel_43_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_8 XI11_3/XI0/XI0_43/d__8_ xsel_43_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_7 XI11_3/XI0/XI0_43/d__7_ xsel_43_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_6 XI11_3/XI0/XI0_43/d__6_ xsel_43_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_5 XI11_3/XI0/XI0_43/d__5_ xsel_43_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_4 XI11_3/XI0/XI0_43/d__4_ xsel_43_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_3 XI11_3/XI0/XI0_43/d__3_ xsel_43_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_2 XI11_3/XI0/XI0_43/d__2_ xsel_43_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_1 XI11_3/XI0/XI0_43/d__1_ xsel_43_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_0 XI11_3/XI0/XI0_43/d__0_ xsel_43_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_15 XI11_3/net21_0_ xsel_42_ XI11_3/XI0/XI0_42/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_14 XI11_3/net21_1_ xsel_42_ XI11_3/XI0/XI0_42/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_13 XI11_3/net21_2_ xsel_42_ XI11_3/XI0/XI0_42/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_12 XI11_3/net21_3_ xsel_42_ XI11_3/XI0/XI0_42/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_11 XI11_3/net21_4_ xsel_42_ XI11_3/XI0/XI0_42/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_10 XI11_3/net21_5_ xsel_42_ XI11_3/XI0/XI0_42/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_9 XI11_3/net21_6_ xsel_42_ XI11_3/XI0/XI0_42/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_8 XI11_3/net21_7_ xsel_42_ XI11_3/XI0/XI0_42/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_7 XI11_3/net21_8_ xsel_42_ XI11_3/XI0/XI0_42/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_6 XI11_3/net21_9_ xsel_42_ XI11_3/XI0/XI0_42/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_5 XI11_3/net21_10_ xsel_42_ XI11_3/XI0/XI0_42/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_4 XI11_3/net21_11_ xsel_42_ XI11_3/XI0/XI0_42/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_3 XI11_3/net21_12_ xsel_42_ XI11_3/XI0/XI0_42/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_2 XI11_3/net21_13_ xsel_42_ XI11_3/XI0/XI0_42/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_1 XI11_3/net21_14_ xsel_42_ XI11_3/XI0/XI0_42/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_0 XI11_3/net21_15_ xsel_42_ XI11_3/XI0/XI0_42/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_15 XI11_3/XI0/XI0_42/d__15_ xsel_42_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_14 XI11_3/XI0/XI0_42/d__14_ xsel_42_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_13 XI11_3/XI0/XI0_42/d__13_ xsel_42_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_12 XI11_3/XI0/XI0_42/d__12_ xsel_42_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_11 XI11_3/XI0/XI0_42/d__11_ xsel_42_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_10 XI11_3/XI0/XI0_42/d__10_ xsel_42_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_9 XI11_3/XI0/XI0_42/d__9_ xsel_42_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_8 XI11_3/XI0/XI0_42/d__8_ xsel_42_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_7 XI11_3/XI0/XI0_42/d__7_ xsel_42_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_6 XI11_3/XI0/XI0_42/d__6_ xsel_42_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_5 XI11_3/XI0/XI0_42/d__5_ xsel_42_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_4 XI11_3/XI0/XI0_42/d__4_ xsel_42_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_3 XI11_3/XI0/XI0_42/d__3_ xsel_42_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_2 XI11_3/XI0/XI0_42/d__2_ xsel_42_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_1 XI11_3/XI0/XI0_42/d__1_ xsel_42_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_0 XI11_3/XI0/XI0_42/d__0_ xsel_42_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_15 XI11_3/net21_0_ xsel_41_ XI11_3/XI0/XI0_41/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_14 XI11_3/net21_1_ xsel_41_ XI11_3/XI0/XI0_41/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_13 XI11_3/net21_2_ xsel_41_ XI11_3/XI0/XI0_41/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_12 XI11_3/net21_3_ xsel_41_ XI11_3/XI0/XI0_41/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_11 XI11_3/net21_4_ xsel_41_ XI11_3/XI0/XI0_41/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_10 XI11_3/net21_5_ xsel_41_ XI11_3/XI0/XI0_41/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_9 XI11_3/net21_6_ xsel_41_ XI11_3/XI0/XI0_41/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_8 XI11_3/net21_7_ xsel_41_ XI11_3/XI0/XI0_41/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_7 XI11_3/net21_8_ xsel_41_ XI11_3/XI0/XI0_41/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_6 XI11_3/net21_9_ xsel_41_ XI11_3/XI0/XI0_41/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_5 XI11_3/net21_10_ xsel_41_ XI11_3/XI0/XI0_41/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_4 XI11_3/net21_11_ xsel_41_ XI11_3/XI0/XI0_41/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_3 XI11_3/net21_12_ xsel_41_ XI11_3/XI0/XI0_41/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_2 XI11_3/net21_13_ xsel_41_ XI11_3/XI0/XI0_41/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_1 XI11_3/net21_14_ xsel_41_ XI11_3/XI0/XI0_41/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_0 XI11_3/net21_15_ xsel_41_ XI11_3/XI0/XI0_41/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_15 XI11_3/XI0/XI0_41/d__15_ xsel_41_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_14 XI11_3/XI0/XI0_41/d__14_ xsel_41_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_13 XI11_3/XI0/XI0_41/d__13_ xsel_41_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_12 XI11_3/XI0/XI0_41/d__12_ xsel_41_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_11 XI11_3/XI0/XI0_41/d__11_ xsel_41_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_10 XI11_3/XI0/XI0_41/d__10_ xsel_41_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_9 XI11_3/XI0/XI0_41/d__9_ xsel_41_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_8 XI11_3/XI0/XI0_41/d__8_ xsel_41_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_7 XI11_3/XI0/XI0_41/d__7_ xsel_41_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_6 XI11_3/XI0/XI0_41/d__6_ xsel_41_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_5 XI11_3/XI0/XI0_41/d__5_ xsel_41_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_4 XI11_3/XI0/XI0_41/d__4_ xsel_41_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_3 XI11_3/XI0/XI0_41/d__3_ xsel_41_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_2 XI11_3/XI0/XI0_41/d__2_ xsel_41_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_1 XI11_3/XI0/XI0_41/d__1_ xsel_41_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_0 XI11_3/XI0/XI0_41/d__0_ xsel_41_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_15 XI11_3/net21_0_ xsel_40_ XI11_3/XI0/XI0_40/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_14 XI11_3/net21_1_ xsel_40_ XI11_3/XI0/XI0_40/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_13 XI11_3/net21_2_ xsel_40_ XI11_3/XI0/XI0_40/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_12 XI11_3/net21_3_ xsel_40_ XI11_3/XI0/XI0_40/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_11 XI11_3/net21_4_ xsel_40_ XI11_3/XI0/XI0_40/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_10 XI11_3/net21_5_ xsel_40_ XI11_3/XI0/XI0_40/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_9 XI11_3/net21_6_ xsel_40_ XI11_3/XI0/XI0_40/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_8 XI11_3/net21_7_ xsel_40_ XI11_3/XI0/XI0_40/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_7 XI11_3/net21_8_ xsel_40_ XI11_3/XI0/XI0_40/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_6 XI11_3/net21_9_ xsel_40_ XI11_3/XI0/XI0_40/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_5 XI11_3/net21_10_ xsel_40_ XI11_3/XI0/XI0_40/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_4 XI11_3/net21_11_ xsel_40_ XI11_3/XI0/XI0_40/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_3 XI11_3/net21_12_ xsel_40_ XI11_3/XI0/XI0_40/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_2 XI11_3/net21_13_ xsel_40_ XI11_3/XI0/XI0_40/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_1 XI11_3/net21_14_ xsel_40_ XI11_3/XI0/XI0_40/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_0 XI11_3/net21_15_ xsel_40_ XI11_3/XI0/XI0_40/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_15 XI11_3/XI0/XI0_40/d__15_ xsel_40_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_14 XI11_3/XI0/XI0_40/d__14_ xsel_40_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_13 XI11_3/XI0/XI0_40/d__13_ xsel_40_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_12 XI11_3/XI0/XI0_40/d__12_ xsel_40_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_11 XI11_3/XI0/XI0_40/d__11_ xsel_40_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_10 XI11_3/XI0/XI0_40/d__10_ xsel_40_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_9 XI11_3/XI0/XI0_40/d__9_ xsel_40_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_8 XI11_3/XI0/XI0_40/d__8_ xsel_40_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_7 XI11_3/XI0/XI0_40/d__7_ xsel_40_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_6 XI11_3/XI0/XI0_40/d__6_ xsel_40_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_5 XI11_3/XI0/XI0_40/d__5_ xsel_40_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_4 XI11_3/XI0/XI0_40/d__4_ xsel_40_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_3 XI11_3/XI0/XI0_40/d__3_ xsel_40_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_2 XI11_3/XI0/XI0_40/d__2_ xsel_40_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_1 XI11_3/XI0/XI0_40/d__1_ xsel_40_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_0 XI11_3/XI0/XI0_40/d__0_ xsel_40_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_15 XI11_3/net21_0_ xsel_39_ XI11_3/XI0/XI0_39/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_14 XI11_3/net21_1_ xsel_39_ XI11_3/XI0/XI0_39/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_13 XI11_3/net21_2_ xsel_39_ XI11_3/XI0/XI0_39/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_12 XI11_3/net21_3_ xsel_39_ XI11_3/XI0/XI0_39/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_11 XI11_3/net21_4_ xsel_39_ XI11_3/XI0/XI0_39/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_10 XI11_3/net21_5_ xsel_39_ XI11_3/XI0/XI0_39/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_9 XI11_3/net21_6_ xsel_39_ XI11_3/XI0/XI0_39/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_8 XI11_3/net21_7_ xsel_39_ XI11_3/XI0/XI0_39/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_7 XI11_3/net21_8_ xsel_39_ XI11_3/XI0/XI0_39/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_6 XI11_3/net21_9_ xsel_39_ XI11_3/XI0/XI0_39/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_5 XI11_3/net21_10_ xsel_39_ XI11_3/XI0/XI0_39/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_4 XI11_3/net21_11_ xsel_39_ XI11_3/XI0/XI0_39/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_3 XI11_3/net21_12_ xsel_39_ XI11_3/XI0/XI0_39/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_2 XI11_3/net21_13_ xsel_39_ XI11_3/XI0/XI0_39/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_1 XI11_3/net21_14_ xsel_39_ XI11_3/XI0/XI0_39/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_0 XI11_3/net21_15_ xsel_39_ XI11_3/XI0/XI0_39/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_15 XI11_3/XI0/XI0_39/d__15_ xsel_39_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_14 XI11_3/XI0/XI0_39/d__14_ xsel_39_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_13 XI11_3/XI0/XI0_39/d__13_ xsel_39_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_12 XI11_3/XI0/XI0_39/d__12_ xsel_39_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_11 XI11_3/XI0/XI0_39/d__11_ xsel_39_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_10 XI11_3/XI0/XI0_39/d__10_ xsel_39_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_9 XI11_3/XI0/XI0_39/d__9_ xsel_39_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_8 XI11_3/XI0/XI0_39/d__8_ xsel_39_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_7 XI11_3/XI0/XI0_39/d__7_ xsel_39_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_6 XI11_3/XI0/XI0_39/d__6_ xsel_39_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_5 XI11_3/XI0/XI0_39/d__5_ xsel_39_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_4 XI11_3/XI0/XI0_39/d__4_ xsel_39_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_3 XI11_3/XI0/XI0_39/d__3_ xsel_39_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_2 XI11_3/XI0/XI0_39/d__2_ xsel_39_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_1 XI11_3/XI0/XI0_39/d__1_ xsel_39_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_0 XI11_3/XI0/XI0_39/d__0_ xsel_39_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_15 XI11_3/net21_0_ xsel_38_ XI11_3/XI0/XI0_38/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_14 XI11_3/net21_1_ xsel_38_ XI11_3/XI0/XI0_38/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_13 XI11_3/net21_2_ xsel_38_ XI11_3/XI0/XI0_38/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_12 XI11_3/net21_3_ xsel_38_ XI11_3/XI0/XI0_38/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_11 XI11_3/net21_4_ xsel_38_ XI11_3/XI0/XI0_38/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_10 XI11_3/net21_5_ xsel_38_ XI11_3/XI0/XI0_38/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_9 XI11_3/net21_6_ xsel_38_ XI11_3/XI0/XI0_38/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_8 XI11_3/net21_7_ xsel_38_ XI11_3/XI0/XI0_38/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_7 XI11_3/net21_8_ xsel_38_ XI11_3/XI0/XI0_38/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_6 XI11_3/net21_9_ xsel_38_ XI11_3/XI0/XI0_38/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_5 XI11_3/net21_10_ xsel_38_ XI11_3/XI0/XI0_38/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_4 XI11_3/net21_11_ xsel_38_ XI11_3/XI0/XI0_38/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_3 XI11_3/net21_12_ xsel_38_ XI11_3/XI0/XI0_38/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_2 XI11_3/net21_13_ xsel_38_ XI11_3/XI0/XI0_38/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_1 XI11_3/net21_14_ xsel_38_ XI11_3/XI0/XI0_38/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_0 XI11_3/net21_15_ xsel_38_ XI11_3/XI0/XI0_38/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_15 XI11_3/XI0/XI0_38/d__15_ xsel_38_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_14 XI11_3/XI0/XI0_38/d__14_ xsel_38_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_13 XI11_3/XI0/XI0_38/d__13_ xsel_38_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_12 XI11_3/XI0/XI0_38/d__12_ xsel_38_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_11 XI11_3/XI0/XI0_38/d__11_ xsel_38_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_10 XI11_3/XI0/XI0_38/d__10_ xsel_38_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_9 XI11_3/XI0/XI0_38/d__9_ xsel_38_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_8 XI11_3/XI0/XI0_38/d__8_ xsel_38_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_7 XI11_3/XI0/XI0_38/d__7_ xsel_38_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_6 XI11_3/XI0/XI0_38/d__6_ xsel_38_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_5 XI11_3/XI0/XI0_38/d__5_ xsel_38_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_4 XI11_3/XI0/XI0_38/d__4_ xsel_38_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_3 XI11_3/XI0/XI0_38/d__3_ xsel_38_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_2 XI11_3/XI0/XI0_38/d__2_ xsel_38_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_1 XI11_3/XI0/XI0_38/d__1_ xsel_38_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_0 XI11_3/XI0/XI0_38/d__0_ xsel_38_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_15 XI11_3/net21_0_ xsel_37_ XI11_3/XI0/XI0_37/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_14 XI11_3/net21_1_ xsel_37_ XI11_3/XI0/XI0_37/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_13 XI11_3/net21_2_ xsel_37_ XI11_3/XI0/XI0_37/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_12 XI11_3/net21_3_ xsel_37_ XI11_3/XI0/XI0_37/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_11 XI11_3/net21_4_ xsel_37_ XI11_3/XI0/XI0_37/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_10 XI11_3/net21_5_ xsel_37_ XI11_3/XI0/XI0_37/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_9 XI11_3/net21_6_ xsel_37_ XI11_3/XI0/XI0_37/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_8 XI11_3/net21_7_ xsel_37_ XI11_3/XI0/XI0_37/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_7 XI11_3/net21_8_ xsel_37_ XI11_3/XI0/XI0_37/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_6 XI11_3/net21_9_ xsel_37_ XI11_3/XI0/XI0_37/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_5 XI11_3/net21_10_ xsel_37_ XI11_3/XI0/XI0_37/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_4 XI11_3/net21_11_ xsel_37_ XI11_3/XI0/XI0_37/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_3 XI11_3/net21_12_ xsel_37_ XI11_3/XI0/XI0_37/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_2 XI11_3/net21_13_ xsel_37_ XI11_3/XI0/XI0_37/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_1 XI11_3/net21_14_ xsel_37_ XI11_3/XI0/XI0_37/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_0 XI11_3/net21_15_ xsel_37_ XI11_3/XI0/XI0_37/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_15 XI11_3/XI0/XI0_37/d__15_ xsel_37_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_14 XI11_3/XI0/XI0_37/d__14_ xsel_37_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_13 XI11_3/XI0/XI0_37/d__13_ xsel_37_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_12 XI11_3/XI0/XI0_37/d__12_ xsel_37_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_11 XI11_3/XI0/XI0_37/d__11_ xsel_37_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_10 XI11_3/XI0/XI0_37/d__10_ xsel_37_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_9 XI11_3/XI0/XI0_37/d__9_ xsel_37_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_8 XI11_3/XI0/XI0_37/d__8_ xsel_37_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_7 XI11_3/XI0/XI0_37/d__7_ xsel_37_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_6 XI11_3/XI0/XI0_37/d__6_ xsel_37_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_5 XI11_3/XI0/XI0_37/d__5_ xsel_37_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_4 XI11_3/XI0/XI0_37/d__4_ xsel_37_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_3 XI11_3/XI0/XI0_37/d__3_ xsel_37_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_2 XI11_3/XI0/XI0_37/d__2_ xsel_37_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_1 XI11_3/XI0/XI0_37/d__1_ xsel_37_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_0 XI11_3/XI0/XI0_37/d__0_ xsel_37_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_15 XI11_3/net21_0_ xsel_36_ XI11_3/XI0/XI0_36/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_14 XI11_3/net21_1_ xsel_36_ XI11_3/XI0/XI0_36/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_13 XI11_3/net21_2_ xsel_36_ XI11_3/XI0/XI0_36/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_12 XI11_3/net21_3_ xsel_36_ XI11_3/XI0/XI0_36/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_11 XI11_3/net21_4_ xsel_36_ XI11_3/XI0/XI0_36/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_10 XI11_3/net21_5_ xsel_36_ XI11_3/XI0/XI0_36/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_9 XI11_3/net21_6_ xsel_36_ XI11_3/XI0/XI0_36/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_8 XI11_3/net21_7_ xsel_36_ XI11_3/XI0/XI0_36/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_7 XI11_3/net21_8_ xsel_36_ XI11_3/XI0/XI0_36/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_6 XI11_3/net21_9_ xsel_36_ XI11_3/XI0/XI0_36/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_5 XI11_3/net21_10_ xsel_36_ XI11_3/XI0/XI0_36/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_4 XI11_3/net21_11_ xsel_36_ XI11_3/XI0/XI0_36/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_3 XI11_3/net21_12_ xsel_36_ XI11_3/XI0/XI0_36/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_2 XI11_3/net21_13_ xsel_36_ XI11_3/XI0/XI0_36/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_1 XI11_3/net21_14_ xsel_36_ XI11_3/XI0/XI0_36/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_0 XI11_3/net21_15_ xsel_36_ XI11_3/XI0/XI0_36/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_15 XI11_3/XI0/XI0_36/d__15_ xsel_36_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_14 XI11_3/XI0/XI0_36/d__14_ xsel_36_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_13 XI11_3/XI0/XI0_36/d__13_ xsel_36_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_12 XI11_3/XI0/XI0_36/d__12_ xsel_36_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_11 XI11_3/XI0/XI0_36/d__11_ xsel_36_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_10 XI11_3/XI0/XI0_36/d__10_ xsel_36_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_9 XI11_3/XI0/XI0_36/d__9_ xsel_36_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_8 XI11_3/XI0/XI0_36/d__8_ xsel_36_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_7 XI11_3/XI0/XI0_36/d__7_ xsel_36_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_6 XI11_3/XI0/XI0_36/d__6_ xsel_36_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_5 XI11_3/XI0/XI0_36/d__5_ xsel_36_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_4 XI11_3/XI0/XI0_36/d__4_ xsel_36_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_3 XI11_3/XI0/XI0_36/d__3_ xsel_36_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_2 XI11_3/XI0/XI0_36/d__2_ xsel_36_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_1 XI11_3/XI0/XI0_36/d__1_ xsel_36_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_0 XI11_3/XI0/XI0_36/d__0_ xsel_36_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_15 XI11_3/net21_0_ xsel_35_ XI11_3/XI0/XI0_35/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_14 XI11_3/net21_1_ xsel_35_ XI11_3/XI0/XI0_35/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_13 XI11_3/net21_2_ xsel_35_ XI11_3/XI0/XI0_35/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_12 XI11_3/net21_3_ xsel_35_ XI11_3/XI0/XI0_35/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_11 XI11_3/net21_4_ xsel_35_ XI11_3/XI0/XI0_35/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_10 XI11_3/net21_5_ xsel_35_ XI11_3/XI0/XI0_35/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_9 XI11_3/net21_6_ xsel_35_ XI11_3/XI0/XI0_35/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_8 XI11_3/net21_7_ xsel_35_ XI11_3/XI0/XI0_35/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_7 XI11_3/net21_8_ xsel_35_ XI11_3/XI0/XI0_35/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_6 XI11_3/net21_9_ xsel_35_ XI11_3/XI0/XI0_35/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_5 XI11_3/net21_10_ xsel_35_ XI11_3/XI0/XI0_35/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_4 XI11_3/net21_11_ xsel_35_ XI11_3/XI0/XI0_35/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_3 XI11_3/net21_12_ xsel_35_ XI11_3/XI0/XI0_35/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_2 XI11_3/net21_13_ xsel_35_ XI11_3/XI0/XI0_35/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_1 XI11_3/net21_14_ xsel_35_ XI11_3/XI0/XI0_35/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_0 XI11_3/net21_15_ xsel_35_ XI11_3/XI0/XI0_35/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_15 XI11_3/XI0/XI0_35/d__15_ xsel_35_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_14 XI11_3/XI0/XI0_35/d__14_ xsel_35_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_13 XI11_3/XI0/XI0_35/d__13_ xsel_35_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_12 XI11_3/XI0/XI0_35/d__12_ xsel_35_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_11 XI11_3/XI0/XI0_35/d__11_ xsel_35_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_10 XI11_3/XI0/XI0_35/d__10_ xsel_35_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_9 XI11_3/XI0/XI0_35/d__9_ xsel_35_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_8 XI11_3/XI0/XI0_35/d__8_ xsel_35_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_7 XI11_3/XI0/XI0_35/d__7_ xsel_35_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_6 XI11_3/XI0/XI0_35/d__6_ xsel_35_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_5 XI11_3/XI0/XI0_35/d__5_ xsel_35_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_4 XI11_3/XI0/XI0_35/d__4_ xsel_35_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_3 XI11_3/XI0/XI0_35/d__3_ xsel_35_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_2 XI11_3/XI0/XI0_35/d__2_ xsel_35_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_1 XI11_3/XI0/XI0_35/d__1_ xsel_35_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_0 XI11_3/XI0/XI0_35/d__0_ xsel_35_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_15 XI11_3/net21_0_ xsel_34_ XI11_3/XI0/XI0_34/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_14 XI11_3/net21_1_ xsel_34_ XI11_3/XI0/XI0_34/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_13 XI11_3/net21_2_ xsel_34_ XI11_3/XI0/XI0_34/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_12 XI11_3/net21_3_ xsel_34_ XI11_3/XI0/XI0_34/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_11 XI11_3/net21_4_ xsel_34_ XI11_3/XI0/XI0_34/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_10 XI11_3/net21_5_ xsel_34_ XI11_3/XI0/XI0_34/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_9 XI11_3/net21_6_ xsel_34_ XI11_3/XI0/XI0_34/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_8 XI11_3/net21_7_ xsel_34_ XI11_3/XI0/XI0_34/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_7 XI11_3/net21_8_ xsel_34_ XI11_3/XI0/XI0_34/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_6 XI11_3/net21_9_ xsel_34_ XI11_3/XI0/XI0_34/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_5 XI11_3/net21_10_ xsel_34_ XI11_3/XI0/XI0_34/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_4 XI11_3/net21_11_ xsel_34_ XI11_3/XI0/XI0_34/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_3 XI11_3/net21_12_ xsel_34_ XI11_3/XI0/XI0_34/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_2 XI11_3/net21_13_ xsel_34_ XI11_3/XI0/XI0_34/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_1 XI11_3/net21_14_ xsel_34_ XI11_3/XI0/XI0_34/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_0 XI11_3/net21_15_ xsel_34_ XI11_3/XI0/XI0_34/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_15 XI11_3/XI0/XI0_34/d__15_ xsel_34_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_14 XI11_3/XI0/XI0_34/d__14_ xsel_34_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_13 XI11_3/XI0/XI0_34/d__13_ xsel_34_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_12 XI11_3/XI0/XI0_34/d__12_ xsel_34_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_11 XI11_3/XI0/XI0_34/d__11_ xsel_34_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_10 XI11_3/XI0/XI0_34/d__10_ xsel_34_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_9 XI11_3/XI0/XI0_34/d__9_ xsel_34_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_8 XI11_3/XI0/XI0_34/d__8_ xsel_34_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_7 XI11_3/XI0/XI0_34/d__7_ xsel_34_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_6 XI11_3/XI0/XI0_34/d__6_ xsel_34_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_5 XI11_3/XI0/XI0_34/d__5_ xsel_34_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_4 XI11_3/XI0/XI0_34/d__4_ xsel_34_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_3 XI11_3/XI0/XI0_34/d__3_ xsel_34_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_2 XI11_3/XI0/XI0_34/d__2_ xsel_34_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_1 XI11_3/XI0/XI0_34/d__1_ xsel_34_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_0 XI11_3/XI0/XI0_34/d__0_ xsel_34_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_15 XI11_3/net21_0_ xsel_33_ XI11_3/XI0/XI0_33/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_14 XI11_3/net21_1_ xsel_33_ XI11_3/XI0/XI0_33/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_13 XI11_3/net21_2_ xsel_33_ XI11_3/XI0/XI0_33/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_12 XI11_3/net21_3_ xsel_33_ XI11_3/XI0/XI0_33/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_11 XI11_3/net21_4_ xsel_33_ XI11_3/XI0/XI0_33/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_10 XI11_3/net21_5_ xsel_33_ XI11_3/XI0/XI0_33/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_9 XI11_3/net21_6_ xsel_33_ XI11_3/XI0/XI0_33/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_8 XI11_3/net21_7_ xsel_33_ XI11_3/XI0/XI0_33/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_7 XI11_3/net21_8_ xsel_33_ XI11_3/XI0/XI0_33/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_6 XI11_3/net21_9_ xsel_33_ XI11_3/XI0/XI0_33/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_5 XI11_3/net21_10_ xsel_33_ XI11_3/XI0/XI0_33/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_4 XI11_3/net21_11_ xsel_33_ XI11_3/XI0/XI0_33/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_3 XI11_3/net21_12_ xsel_33_ XI11_3/XI0/XI0_33/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_2 XI11_3/net21_13_ xsel_33_ XI11_3/XI0/XI0_33/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_1 XI11_3/net21_14_ xsel_33_ XI11_3/XI0/XI0_33/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_0 XI11_3/net21_15_ xsel_33_ XI11_3/XI0/XI0_33/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_15 XI11_3/XI0/XI0_33/d__15_ xsel_33_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_14 XI11_3/XI0/XI0_33/d__14_ xsel_33_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_13 XI11_3/XI0/XI0_33/d__13_ xsel_33_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_12 XI11_3/XI0/XI0_33/d__12_ xsel_33_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_11 XI11_3/XI0/XI0_33/d__11_ xsel_33_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_10 XI11_3/XI0/XI0_33/d__10_ xsel_33_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_9 XI11_3/XI0/XI0_33/d__9_ xsel_33_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_8 XI11_3/XI0/XI0_33/d__8_ xsel_33_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_7 XI11_3/XI0/XI0_33/d__7_ xsel_33_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_6 XI11_3/XI0/XI0_33/d__6_ xsel_33_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_5 XI11_3/XI0/XI0_33/d__5_ xsel_33_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_4 XI11_3/XI0/XI0_33/d__4_ xsel_33_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_3 XI11_3/XI0/XI0_33/d__3_ xsel_33_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_2 XI11_3/XI0/XI0_33/d__2_ xsel_33_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_1 XI11_3/XI0/XI0_33/d__1_ xsel_33_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_0 XI11_3/XI0/XI0_33/d__0_ xsel_33_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_15 XI11_3/net21_0_ xsel_32_ XI11_3/XI0/XI0_32/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_14 XI11_3/net21_1_ xsel_32_ XI11_3/XI0/XI0_32/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_13 XI11_3/net21_2_ xsel_32_ XI11_3/XI0/XI0_32/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_12 XI11_3/net21_3_ xsel_32_ XI11_3/XI0/XI0_32/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_11 XI11_3/net21_4_ xsel_32_ XI11_3/XI0/XI0_32/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_10 XI11_3/net21_5_ xsel_32_ XI11_3/XI0/XI0_32/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_9 XI11_3/net21_6_ xsel_32_ XI11_3/XI0/XI0_32/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_8 XI11_3/net21_7_ xsel_32_ XI11_3/XI0/XI0_32/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_7 XI11_3/net21_8_ xsel_32_ XI11_3/XI0/XI0_32/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_6 XI11_3/net21_9_ xsel_32_ XI11_3/XI0/XI0_32/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_5 XI11_3/net21_10_ xsel_32_ XI11_3/XI0/XI0_32/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_4 XI11_3/net21_11_ xsel_32_ XI11_3/XI0/XI0_32/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_3 XI11_3/net21_12_ xsel_32_ XI11_3/XI0/XI0_32/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_2 XI11_3/net21_13_ xsel_32_ XI11_3/XI0/XI0_32/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_1 XI11_3/net21_14_ xsel_32_ XI11_3/XI0/XI0_32/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_0 XI11_3/net21_15_ xsel_32_ XI11_3/XI0/XI0_32/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_15 XI11_3/XI0/XI0_32/d__15_ xsel_32_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_14 XI11_3/XI0/XI0_32/d__14_ xsel_32_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_13 XI11_3/XI0/XI0_32/d__13_ xsel_32_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_12 XI11_3/XI0/XI0_32/d__12_ xsel_32_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_11 XI11_3/XI0/XI0_32/d__11_ xsel_32_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_10 XI11_3/XI0/XI0_32/d__10_ xsel_32_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_9 XI11_3/XI0/XI0_32/d__9_ xsel_32_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_8 XI11_3/XI0/XI0_32/d__8_ xsel_32_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_7 XI11_3/XI0/XI0_32/d__7_ xsel_32_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_6 XI11_3/XI0/XI0_32/d__6_ xsel_32_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_5 XI11_3/XI0/XI0_32/d__5_ xsel_32_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_4 XI11_3/XI0/XI0_32/d__4_ xsel_32_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_3 XI11_3/XI0/XI0_32/d__3_ xsel_32_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_2 XI11_3/XI0/XI0_32/d__2_ xsel_32_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_1 XI11_3/XI0/XI0_32/d__1_ xsel_32_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_0 XI11_3/XI0/XI0_32/d__0_ xsel_32_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_15 XI11_3/net21_0_ xsel_31_ XI11_3/XI0/XI0_31/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_14 XI11_3/net21_1_ xsel_31_ XI11_3/XI0/XI0_31/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_13 XI11_3/net21_2_ xsel_31_ XI11_3/XI0/XI0_31/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_12 XI11_3/net21_3_ xsel_31_ XI11_3/XI0/XI0_31/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_11 XI11_3/net21_4_ xsel_31_ XI11_3/XI0/XI0_31/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_10 XI11_3/net21_5_ xsel_31_ XI11_3/XI0/XI0_31/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_9 XI11_3/net21_6_ xsel_31_ XI11_3/XI0/XI0_31/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_8 XI11_3/net21_7_ xsel_31_ XI11_3/XI0/XI0_31/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_7 XI11_3/net21_8_ xsel_31_ XI11_3/XI0/XI0_31/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_6 XI11_3/net21_9_ xsel_31_ XI11_3/XI0/XI0_31/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_5 XI11_3/net21_10_ xsel_31_ XI11_3/XI0/XI0_31/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_4 XI11_3/net21_11_ xsel_31_ XI11_3/XI0/XI0_31/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_3 XI11_3/net21_12_ xsel_31_ XI11_3/XI0/XI0_31/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_2 XI11_3/net21_13_ xsel_31_ XI11_3/XI0/XI0_31/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_1 XI11_3/net21_14_ xsel_31_ XI11_3/XI0/XI0_31/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_0 XI11_3/net21_15_ xsel_31_ XI11_3/XI0/XI0_31/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_15 XI11_3/XI0/XI0_31/d__15_ xsel_31_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_14 XI11_3/XI0/XI0_31/d__14_ xsel_31_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_13 XI11_3/XI0/XI0_31/d__13_ xsel_31_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_12 XI11_3/XI0/XI0_31/d__12_ xsel_31_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_11 XI11_3/XI0/XI0_31/d__11_ xsel_31_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_10 XI11_3/XI0/XI0_31/d__10_ xsel_31_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_9 XI11_3/XI0/XI0_31/d__9_ xsel_31_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_8 XI11_3/XI0/XI0_31/d__8_ xsel_31_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_7 XI11_3/XI0/XI0_31/d__7_ xsel_31_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_6 XI11_3/XI0/XI0_31/d__6_ xsel_31_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_5 XI11_3/XI0/XI0_31/d__5_ xsel_31_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_4 XI11_3/XI0/XI0_31/d__4_ xsel_31_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_3 XI11_3/XI0/XI0_31/d__3_ xsel_31_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_2 XI11_3/XI0/XI0_31/d__2_ xsel_31_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_1 XI11_3/XI0/XI0_31/d__1_ xsel_31_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_0 XI11_3/XI0/XI0_31/d__0_ xsel_31_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_15 XI11_3/net21_0_ xsel_30_ XI11_3/XI0/XI0_30/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_14 XI11_3/net21_1_ xsel_30_ XI11_3/XI0/XI0_30/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_13 XI11_3/net21_2_ xsel_30_ XI11_3/XI0/XI0_30/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_12 XI11_3/net21_3_ xsel_30_ XI11_3/XI0/XI0_30/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_11 XI11_3/net21_4_ xsel_30_ XI11_3/XI0/XI0_30/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_10 XI11_3/net21_5_ xsel_30_ XI11_3/XI0/XI0_30/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_9 XI11_3/net21_6_ xsel_30_ XI11_3/XI0/XI0_30/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_8 XI11_3/net21_7_ xsel_30_ XI11_3/XI0/XI0_30/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_7 XI11_3/net21_8_ xsel_30_ XI11_3/XI0/XI0_30/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_6 XI11_3/net21_9_ xsel_30_ XI11_3/XI0/XI0_30/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_5 XI11_3/net21_10_ xsel_30_ XI11_3/XI0/XI0_30/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_4 XI11_3/net21_11_ xsel_30_ XI11_3/XI0/XI0_30/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_3 XI11_3/net21_12_ xsel_30_ XI11_3/XI0/XI0_30/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_2 XI11_3/net21_13_ xsel_30_ XI11_3/XI0/XI0_30/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_1 XI11_3/net21_14_ xsel_30_ XI11_3/XI0/XI0_30/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_0 XI11_3/net21_15_ xsel_30_ XI11_3/XI0/XI0_30/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_15 XI11_3/XI0/XI0_30/d__15_ xsel_30_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_14 XI11_3/XI0/XI0_30/d__14_ xsel_30_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_13 XI11_3/XI0/XI0_30/d__13_ xsel_30_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_12 XI11_3/XI0/XI0_30/d__12_ xsel_30_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_11 XI11_3/XI0/XI0_30/d__11_ xsel_30_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_10 XI11_3/XI0/XI0_30/d__10_ xsel_30_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_9 XI11_3/XI0/XI0_30/d__9_ xsel_30_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_8 XI11_3/XI0/XI0_30/d__8_ xsel_30_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_7 XI11_3/XI0/XI0_30/d__7_ xsel_30_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_6 XI11_3/XI0/XI0_30/d__6_ xsel_30_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_5 XI11_3/XI0/XI0_30/d__5_ xsel_30_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_4 XI11_3/XI0/XI0_30/d__4_ xsel_30_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_3 XI11_3/XI0/XI0_30/d__3_ xsel_30_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_2 XI11_3/XI0/XI0_30/d__2_ xsel_30_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_1 XI11_3/XI0/XI0_30/d__1_ xsel_30_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_0 XI11_3/XI0/XI0_30/d__0_ xsel_30_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_15 XI11_3/net21_0_ xsel_29_ XI11_3/XI0/XI0_29/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_14 XI11_3/net21_1_ xsel_29_ XI11_3/XI0/XI0_29/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_13 XI11_3/net21_2_ xsel_29_ XI11_3/XI0/XI0_29/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_12 XI11_3/net21_3_ xsel_29_ XI11_3/XI0/XI0_29/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_11 XI11_3/net21_4_ xsel_29_ XI11_3/XI0/XI0_29/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_10 XI11_3/net21_5_ xsel_29_ XI11_3/XI0/XI0_29/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_9 XI11_3/net21_6_ xsel_29_ XI11_3/XI0/XI0_29/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_8 XI11_3/net21_7_ xsel_29_ XI11_3/XI0/XI0_29/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_7 XI11_3/net21_8_ xsel_29_ XI11_3/XI0/XI0_29/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_6 XI11_3/net21_9_ xsel_29_ XI11_3/XI0/XI0_29/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_5 XI11_3/net21_10_ xsel_29_ XI11_3/XI0/XI0_29/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_4 XI11_3/net21_11_ xsel_29_ XI11_3/XI0/XI0_29/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_3 XI11_3/net21_12_ xsel_29_ XI11_3/XI0/XI0_29/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_2 XI11_3/net21_13_ xsel_29_ XI11_3/XI0/XI0_29/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_1 XI11_3/net21_14_ xsel_29_ XI11_3/XI0/XI0_29/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_0 XI11_3/net21_15_ xsel_29_ XI11_3/XI0/XI0_29/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_15 XI11_3/XI0/XI0_29/d__15_ xsel_29_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_14 XI11_3/XI0/XI0_29/d__14_ xsel_29_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_13 XI11_3/XI0/XI0_29/d__13_ xsel_29_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_12 XI11_3/XI0/XI0_29/d__12_ xsel_29_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_11 XI11_3/XI0/XI0_29/d__11_ xsel_29_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_10 XI11_3/XI0/XI0_29/d__10_ xsel_29_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_9 XI11_3/XI0/XI0_29/d__9_ xsel_29_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_8 XI11_3/XI0/XI0_29/d__8_ xsel_29_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_7 XI11_3/XI0/XI0_29/d__7_ xsel_29_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_6 XI11_3/XI0/XI0_29/d__6_ xsel_29_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_5 XI11_3/XI0/XI0_29/d__5_ xsel_29_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_4 XI11_3/XI0/XI0_29/d__4_ xsel_29_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_3 XI11_3/XI0/XI0_29/d__3_ xsel_29_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_2 XI11_3/XI0/XI0_29/d__2_ xsel_29_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_1 XI11_3/XI0/XI0_29/d__1_ xsel_29_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_0 XI11_3/XI0/XI0_29/d__0_ xsel_29_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_15 XI11_3/net21_0_ xsel_28_ XI11_3/XI0/XI0_28/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_14 XI11_3/net21_1_ xsel_28_ XI11_3/XI0/XI0_28/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_13 XI11_3/net21_2_ xsel_28_ XI11_3/XI0/XI0_28/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_12 XI11_3/net21_3_ xsel_28_ XI11_3/XI0/XI0_28/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_11 XI11_3/net21_4_ xsel_28_ XI11_3/XI0/XI0_28/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_10 XI11_3/net21_5_ xsel_28_ XI11_3/XI0/XI0_28/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_9 XI11_3/net21_6_ xsel_28_ XI11_3/XI0/XI0_28/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_8 XI11_3/net21_7_ xsel_28_ XI11_3/XI0/XI0_28/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_7 XI11_3/net21_8_ xsel_28_ XI11_3/XI0/XI0_28/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_6 XI11_3/net21_9_ xsel_28_ XI11_3/XI0/XI0_28/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_5 XI11_3/net21_10_ xsel_28_ XI11_3/XI0/XI0_28/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_4 XI11_3/net21_11_ xsel_28_ XI11_3/XI0/XI0_28/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_3 XI11_3/net21_12_ xsel_28_ XI11_3/XI0/XI0_28/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_2 XI11_3/net21_13_ xsel_28_ XI11_3/XI0/XI0_28/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_1 XI11_3/net21_14_ xsel_28_ XI11_3/XI0/XI0_28/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_0 XI11_3/net21_15_ xsel_28_ XI11_3/XI0/XI0_28/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_15 XI11_3/XI0/XI0_28/d__15_ xsel_28_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_14 XI11_3/XI0/XI0_28/d__14_ xsel_28_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_13 XI11_3/XI0/XI0_28/d__13_ xsel_28_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_12 XI11_3/XI0/XI0_28/d__12_ xsel_28_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_11 XI11_3/XI0/XI0_28/d__11_ xsel_28_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_10 XI11_3/XI0/XI0_28/d__10_ xsel_28_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_9 XI11_3/XI0/XI0_28/d__9_ xsel_28_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_8 XI11_3/XI0/XI0_28/d__8_ xsel_28_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_7 XI11_3/XI0/XI0_28/d__7_ xsel_28_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_6 XI11_3/XI0/XI0_28/d__6_ xsel_28_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_5 XI11_3/XI0/XI0_28/d__5_ xsel_28_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_4 XI11_3/XI0/XI0_28/d__4_ xsel_28_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_3 XI11_3/XI0/XI0_28/d__3_ xsel_28_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_2 XI11_3/XI0/XI0_28/d__2_ xsel_28_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_1 XI11_3/XI0/XI0_28/d__1_ xsel_28_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_0 XI11_3/XI0/XI0_28/d__0_ xsel_28_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_15 XI11_3/net21_0_ xsel_27_ XI11_3/XI0/XI0_27/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_14 XI11_3/net21_1_ xsel_27_ XI11_3/XI0/XI0_27/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_13 XI11_3/net21_2_ xsel_27_ XI11_3/XI0/XI0_27/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_12 XI11_3/net21_3_ xsel_27_ XI11_3/XI0/XI0_27/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_11 XI11_3/net21_4_ xsel_27_ XI11_3/XI0/XI0_27/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_10 XI11_3/net21_5_ xsel_27_ XI11_3/XI0/XI0_27/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_9 XI11_3/net21_6_ xsel_27_ XI11_3/XI0/XI0_27/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_8 XI11_3/net21_7_ xsel_27_ XI11_3/XI0/XI0_27/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_7 XI11_3/net21_8_ xsel_27_ XI11_3/XI0/XI0_27/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_6 XI11_3/net21_9_ xsel_27_ XI11_3/XI0/XI0_27/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_5 XI11_3/net21_10_ xsel_27_ XI11_3/XI0/XI0_27/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_4 XI11_3/net21_11_ xsel_27_ XI11_3/XI0/XI0_27/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_3 XI11_3/net21_12_ xsel_27_ XI11_3/XI0/XI0_27/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_2 XI11_3/net21_13_ xsel_27_ XI11_3/XI0/XI0_27/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_1 XI11_3/net21_14_ xsel_27_ XI11_3/XI0/XI0_27/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_0 XI11_3/net21_15_ xsel_27_ XI11_3/XI0/XI0_27/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_15 XI11_3/XI0/XI0_27/d__15_ xsel_27_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_14 XI11_3/XI0/XI0_27/d__14_ xsel_27_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_13 XI11_3/XI0/XI0_27/d__13_ xsel_27_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_12 XI11_3/XI0/XI0_27/d__12_ xsel_27_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_11 XI11_3/XI0/XI0_27/d__11_ xsel_27_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_10 XI11_3/XI0/XI0_27/d__10_ xsel_27_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_9 XI11_3/XI0/XI0_27/d__9_ xsel_27_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_8 XI11_3/XI0/XI0_27/d__8_ xsel_27_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_7 XI11_3/XI0/XI0_27/d__7_ xsel_27_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_6 XI11_3/XI0/XI0_27/d__6_ xsel_27_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_5 XI11_3/XI0/XI0_27/d__5_ xsel_27_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_4 XI11_3/XI0/XI0_27/d__4_ xsel_27_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_3 XI11_3/XI0/XI0_27/d__3_ xsel_27_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_2 XI11_3/XI0/XI0_27/d__2_ xsel_27_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_1 XI11_3/XI0/XI0_27/d__1_ xsel_27_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_0 XI11_3/XI0/XI0_27/d__0_ xsel_27_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_15 XI11_3/net21_0_ xsel_26_ XI11_3/XI0/XI0_26/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_14 XI11_3/net21_1_ xsel_26_ XI11_3/XI0/XI0_26/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_13 XI11_3/net21_2_ xsel_26_ XI11_3/XI0/XI0_26/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_12 XI11_3/net21_3_ xsel_26_ XI11_3/XI0/XI0_26/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_11 XI11_3/net21_4_ xsel_26_ XI11_3/XI0/XI0_26/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_10 XI11_3/net21_5_ xsel_26_ XI11_3/XI0/XI0_26/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_9 XI11_3/net21_6_ xsel_26_ XI11_3/XI0/XI0_26/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_8 XI11_3/net21_7_ xsel_26_ XI11_3/XI0/XI0_26/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_7 XI11_3/net21_8_ xsel_26_ XI11_3/XI0/XI0_26/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_6 XI11_3/net21_9_ xsel_26_ XI11_3/XI0/XI0_26/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_5 XI11_3/net21_10_ xsel_26_ XI11_3/XI0/XI0_26/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_4 XI11_3/net21_11_ xsel_26_ XI11_3/XI0/XI0_26/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_3 XI11_3/net21_12_ xsel_26_ XI11_3/XI0/XI0_26/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_2 XI11_3/net21_13_ xsel_26_ XI11_3/XI0/XI0_26/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_1 XI11_3/net21_14_ xsel_26_ XI11_3/XI0/XI0_26/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_0 XI11_3/net21_15_ xsel_26_ XI11_3/XI0/XI0_26/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_15 XI11_3/XI0/XI0_26/d__15_ xsel_26_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_14 XI11_3/XI0/XI0_26/d__14_ xsel_26_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_13 XI11_3/XI0/XI0_26/d__13_ xsel_26_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_12 XI11_3/XI0/XI0_26/d__12_ xsel_26_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_11 XI11_3/XI0/XI0_26/d__11_ xsel_26_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_10 XI11_3/XI0/XI0_26/d__10_ xsel_26_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_9 XI11_3/XI0/XI0_26/d__9_ xsel_26_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_8 XI11_3/XI0/XI0_26/d__8_ xsel_26_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_7 XI11_3/XI0/XI0_26/d__7_ xsel_26_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_6 XI11_3/XI0/XI0_26/d__6_ xsel_26_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_5 XI11_3/XI0/XI0_26/d__5_ xsel_26_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_4 XI11_3/XI0/XI0_26/d__4_ xsel_26_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_3 XI11_3/XI0/XI0_26/d__3_ xsel_26_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_2 XI11_3/XI0/XI0_26/d__2_ xsel_26_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_1 XI11_3/XI0/XI0_26/d__1_ xsel_26_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_0 XI11_3/XI0/XI0_26/d__0_ xsel_26_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_15 XI11_3/net21_0_ xsel_25_ XI11_3/XI0/XI0_25/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_14 XI11_3/net21_1_ xsel_25_ XI11_3/XI0/XI0_25/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_13 XI11_3/net21_2_ xsel_25_ XI11_3/XI0/XI0_25/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_12 XI11_3/net21_3_ xsel_25_ XI11_3/XI0/XI0_25/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_11 XI11_3/net21_4_ xsel_25_ XI11_3/XI0/XI0_25/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_10 XI11_3/net21_5_ xsel_25_ XI11_3/XI0/XI0_25/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_9 XI11_3/net21_6_ xsel_25_ XI11_3/XI0/XI0_25/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_8 XI11_3/net21_7_ xsel_25_ XI11_3/XI0/XI0_25/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_7 XI11_3/net21_8_ xsel_25_ XI11_3/XI0/XI0_25/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_6 XI11_3/net21_9_ xsel_25_ XI11_3/XI0/XI0_25/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_5 XI11_3/net21_10_ xsel_25_ XI11_3/XI0/XI0_25/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_4 XI11_3/net21_11_ xsel_25_ XI11_3/XI0/XI0_25/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_3 XI11_3/net21_12_ xsel_25_ XI11_3/XI0/XI0_25/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_2 XI11_3/net21_13_ xsel_25_ XI11_3/XI0/XI0_25/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_1 XI11_3/net21_14_ xsel_25_ XI11_3/XI0/XI0_25/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_0 XI11_3/net21_15_ xsel_25_ XI11_3/XI0/XI0_25/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN1_15 XI11_3/XI0/XI0_25/d__15_ xsel_25_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN1_14 XI11_3/XI0/XI0_25/d__14_ xsel_25_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN1_13 XI11_3/XI0/XI0_25/d__13_ xsel_25_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN1_12 XI11_3/XI0/XI0_25/d__12_ xsel_25_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN1_11 XI11_3/XI0/XI0_25/d__11_ xsel_25_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN1_10 XI11_3/XI0/XI0_25/d__10_ xsel_25_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN1_9 XI11_3/XI0/XI0_25/d__9_ xsel_25_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN1_8 XI11_3/XI0/XI0_25/d__8_ xsel_25_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN1_7 XI11_3/XI0/XI0_25/d__7_ xsel_25_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN1_6 XI11_3/XI0/XI0_25/d__6_ xsel_25_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN1_5 XI11_3/XI0/XI0_25/d__5_ xsel_25_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN1_4 XI11_3/XI0/XI0_25/d__4_ xsel_25_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN1_3 XI11_3/XI0/XI0_25/d__3_ xsel_25_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN1_2 XI11_3/XI0/XI0_25/d__2_ xsel_25_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN1_1 XI11_3/XI0/XI0_25/d__1_ xsel_25_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN1_0 XI11_3/XI0/XI0_25/d__0_ xsel_25_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN0_15 XI11_3/net21_0_ xsel_24_ XI11_3/XI0/XI0_24/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN0_14 XI11_3/net21_1_ xsel_24_ XI11_3/XI0/XI0_24/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN0_13 XI11_3/net21_2_ xsel_24_ XI11_3/XI0/XI0_24/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN0_12 XI11_3/net21_3_ xsel_24_ XI11_3/XI0/XI0_24/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN0_11 XI11_3/net21_4_ xsel_24_ XI11_3/XI0/XI0_24/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN0_10 XI11_3/net21_5_ xsel_24_ XI11_3/XI0/XI0_24/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN0_9 XI11_3/net21_6_ xsel_24_ XI11_3/XI0/XI0_24/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN0_8 XI11_3/net21_7_ xsel_24_ XI11_3/XI0/XI0_24/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN0_7 XI11_3/net21_8_ xsel_24_ XI11_3/XI0/XI0_24/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN0_6 XI11_3/net21_9_ xsel_24_ XI11_3/XI0/XI0_24/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN0_5 XI11_3/net21_10_ xsel_24_ XI11_3/XI0/XI0_24/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN0_4 XI11_3/net21_11_ xsel_24_ XI11_3/XI0/XI0_24/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN0_3 XI11_3/net21_12_ xsel_24_ XI11_3/XI0/XI0_24/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN0_2 XI11_3/net21_13_ xsel_24_ XI11_3/XI0/XI0_24/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN0_1 XI11_3/net21_14_ xsel_24_ XI11_3/XI0/XI0_24/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN0_0 XI11_3/net21_15_ xsel_24_ XI11_3/XI0/XI0_24/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN1_15 XI11_3/XI0/XI0_24/d__15_ xsel_24_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN1_14 XI11_3/XI0/XI0_24/d__14_ xsel_24_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN1_13 XI11_3/XI0/XI0_24/d__13_ xsel_24_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN1_12 XI11_3/XI0/XI0_24/d__12_ xsel_24_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN1_11 XI11_3/XI0/XI0_24/d__11_ xsel_24_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN1_10 XI11_3/XI0/XI0_24/d__10_ xsel_24_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN1_9 XI11_3/XI0/XI0_24/d__9_ xsel_24_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN1_8 XI11_3/XI0/XI0_24/d__8_ xsel_24_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN1_7 XI11_3/XI0/XI0_24/d__7_ xsel_24_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN1_6 XI11_3/XI0/XI0_24/d__6_ xsel_24_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN1_5 XI11_3/XI0/XI0_24/d__5_ xsel_24_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN1_4 XI11_3/XI0/XI0_24/d__4_ xsel_24_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN1_3 XI11_3/XI0/XI0_24/d__3_ xsel_24_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN1_2 XI11_3/XI0/XI0_24/d__2_ xsel_24_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN1_1 XI11_3/XI0/XI0_24/d__1_ xsel_24_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_24/MN1_0 XI11_3/XI0/XI0_24/d__0_ xsel_24_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN0_15 XI11_3/net21_0_ xsel_23_ XI11_3/XI0/XI0_23/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN0_14 XI11_3/net21_1_ xsel_23_ XI11_3/XI0/XI0_23/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN0_13 XI11_3/net21_2_ xsel_23_ XI11_3/XI0/XI0_23/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN0_12 XI11_3/net21_3_ xsel_23_ XI11_3/XI0/XI0_23/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN0_11 XI11_3/net21_4_ xsel_23_ XI11_3/XI0/XI0_23/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN0_10 XI11_3/net21_5_ xsel_23_ XI11_3/XI0/XI0_23/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN0_9 XI11_3/net21_6_ xsel_23_ XI11_3/XI0/XI0_23/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN0_8 XI11_3/net21_7_ xsel_23_ XI11_3/XI0/XI0_23/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN0_7 XI11_3/net21_8_ xsel_23_ XI11_3/XI0/XI0_23/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN0_6 XI11_3/net21_9_ xsel_23_ XI11_3/XI0/XI0_23/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN0_5 XI11_3/net21_10_ xsel_23_ XI11_3/XI0/XI0_23/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN0_4 XI11_3/net21_11_ xsel_23_ XI11_3/XI0/XI0_23/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN0_3 XI11_3/net21_12_ xsel_23_ XI11_3/XI0/XI0_23/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN0_2 XI11_3/net21_13_ xsel_23_ XI11_3/XI0/XI0_23/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN0_1 XI11_3/net21_14_ xsel_23_ XI11_3/XI0/XI0_23/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN0_0 XI11_3/net21_15_ xsel_23_ XI11_3/XI0/XI0_23/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN1_15 XI11_3/XI0/XI0_23/d__15_ xsel_23_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN1_14 XI11_3/XI0/XI0_23/d__14_ xsel_23_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN1_13 XI11_3/XI0/XI0_23/d__13_ xsel_23_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN1_12 XI11_3/XI0/XI0_23/d__12_ xsel_23_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN1_11 XI11_3/XI0/XI0_23/d__11_ xsel_23_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN1_10 XI11_3/XI0/XI0_23/d__10_ xsel_23_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN1_9 XI11_3/XI0/XI0_23/d__9_ xsel_23_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN1_8 XI11_3/XI0/XI0_23/d__8_ xsel_23_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN1_7 XI11_3/XI0/XI0_23/d__7_ xsel_23_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN1_6 XI11_3/XI0/XI0_23/d__6_ xsel_23_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN1_5 XI11_3/XI0/XI0_23/d__5_ xsel_23_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN1_4 XI11_3/XI0/XI0_23/d__4_ xsel_23_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN1_3 XI11_3/XI0/XI0_23/d__3_ xsel_23_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN1_2 XI11_3/XI0/XI0_23/d__2_ xsel_23_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN1_1 XI11_3/XI0/XI0_23/d__1_ xsel_23_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_23/MN1_0 XI11_3/XI0/XI0_23/d__0_ xsel_23_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN0_15 XI11_3/net21_0_ xsel_22_ XI11_3/XI0/XI0_22/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN0_14 XI11_3/net21_1_ xsel_22_ XI11_3/XI0/XI0_22/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN0_13 XI11_3/net21_2_ xsel_22_ XI11_3/XI0/XI0_22/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN0_12 XI11_3/net21_3_ xsel_22_ XI11_3/XI0/XI0_22/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN0_11 XI11_3/net21_4_ xsel_22_ XI11_3/XI0/XI0_22/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN0_10 XI11_3/net21_5_ xsel_22_ XI11_3/XI0/XI0_22/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN0_9 XI11_3/net21_6_ xsel_22_ XI11_3/XI0/XI0_22/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN0_8 XI11_3/net21_7_ xsel_22_ XI11_3/XI0/XI0_22/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN0_7 XI11_3/net21_8_ xsel_22_ XI11_3/XI0/XI0_22/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN0_6 XI11_3/net21_9_ xsel_22_ XI11_3/XI0/XI0_22/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN0_5 XI11_3/net21_10_ xsel_22_ XI11_3/XI0/XI0_22/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN0_4 XI11_3/net21_11_ xsel_22_ XI11_3/XI0/XI0_22/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN0_3 XI11_3/net21_12_ xsel_22_ XI11_3/XI0/XI0_22/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN0_2 XI11_3/net21_13_ xsel_22_ XI11_3/XI0/XI0_22/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN0_1 XI11_3/net21_14_ xsel_22_ XI11_3/XI0/XI0_22/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN0_0 XI11_3/net21_15_ xsel_22_ XI11_3/XI0/XI0_22/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN1_15 XI11_3/XI0/XI0_22/d__15_ xsel_22_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN1_14 XI11_3/XI0/XI0_22/d__14_ xsel_22_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN1_13 XI11_3/XI0/XI0_22/d__13_ xsel_22_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN1_12 XI11_3/XI0/XI0_22/d__12_ xsel_22_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN1_11 XI11_3/XI0/XI0_22/d__11_ xsel_22_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN1_10 XI11_3/XI0/XI0_22/d__10_ xsel_22_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN1_9 XI11_3/XI0/XI0_22/d__9_ xsel_22_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN1_8 XI11_3/XI0/XI0_22/d__8_ xsel_22_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN1_7 XI11_3/XI0/XI0_22/d__7_ xsel_22_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN1_6 XI11_3/XI0/XI0_22/d__6_ xsel_22_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN1_5 XI11_3/XI0/XI0_22/d__5_ xsel_22_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN1_4 XI11_3/XI0/XI0_22/d__4_ xsel_22_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN1_3 XI11_3/XI0/XI0_22/d__3_ xsel_22_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN1_2 XI11_3/XI0/XI0_22/d__2_ xsel_22_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN1_1 XI11_3/XI0/XI0_22/d__1_ xsel_22_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_22/MN1_0 XI11_3/XI0/XI0_22/d__0_ xsel_22_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN0_15 XI11_3/net21_0_ xsel_21_ XI11_3/XI0/XI0_21/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN0_14 XI11_3/net21_1_ xsel_21_ XI11_3/XI0/XI0_21/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN0_13 XI11_3/net21_2_ xsel_21_ XI11_3/XI0/XI0_21/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN0_12 XI11_3/net21_3_ xsel_21_ XI11_3/XI0/XI0_21/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN0_11 XI11_3/net21_4_ xsel_21_ XI11_3/XI0/XI0_21/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN0_10 XI11_3/net21_5_ xsel_21_ XI11_3/XI0/XI0_21/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN0_9 XI11_3/net21_6_ xsel_21_ XI11_3/XI0/XI0_21/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN0_8 XI11_3/net21_7_ xsel_21_ XI11_3/XI0/XI0_21/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN0_7 XI11_3/net21_8_ xsel_21_ XI11_3/XI0/XI0_21/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN0_6 XI11_3/net21_9_ xsel_21_ XI11_3/XI0/XI0_21/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN0_5 XI11_3/net21_10_ xsel_21_ XI11_3/XI0/XI0_21/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN0_4 XI11_3/net21_11_ xsel_21_ XI11_3/XI0/XI0_21/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN0_3 XI11_3/net21_12_ xsel_21_ XI11_3/XI0/XI0_21/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN0_2 XI11_3/net21_13_ xsel_21_ XI11_3/XI0/XI0_21/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN0_1 XI11_3/net21_14_ xsel_21_ XI11_3/XI0/XI0_21/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN0_0 XI11_3/net21_15_ xsel_21_ XI11_3/XI0/XI0_21/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN1_15 XI11_3/XI0/XI0_21/d__15_ xsel_21_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN1_14 XI11_3/XI0/XI0_21/d__14_ xsel_21_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN1_13 XI11_3/XI0/XI0_21/d__13_ xsel_21_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN1_12 XI11_3/XI0/XI0_21/d__12_ xsel_21_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN1_11 XI11_3/XI0/XI0_21/d__11_ xsel_21_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN1_10 XI11_3/XI0/XI0_21/d__10_ xsel_21_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN1_9 XI11_3/XI0/XI0_21/d__9_ xsel_21_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN1_8 XI11_3/XI0/XI0_21/d__8_ xsel_21_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN1_7 XI11_3/XI0/XI0_21/d__7_ xsel_21_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN1_6 XI11_3/XI0/XI0_21/d__6_ xsel_21_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN1_5 XI11_3/XI0/XI0_21/d__5_ xsel_21_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN1_4 XI11_3/XI0/XI0_21/d__4_ xsel_21_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN1_3 XI11_3/XI0/XI0_21/d__3_ xsel_21_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN1_2 XI11_3/XI0/XI0_21/d__2_ xsel_21_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN1_1 XI11_3/XI0/XI0_21/d__1_ xsel_21_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_21/MN1_0 XI11_3/XI0/XI0_21/d__0_ xsel_21_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN0_15 XI11_3/net21_0_ xsel_20_ XI11_3/XI0/XI0_20/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN0_14 XI11_3/net21_1_ xsel_20_ XI11_3/XI0/XI0_20/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN0_13 XI11_3/net21_2_ xsel_20_ XI11_3/XI0/XI0_20/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN0_12 XI11_3/net21_3_ xsel_20_ XI11_3/XI0/XI0_20/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN0_11 XI11_3/net21_4_ xsel_20_ XI11_3/XI0/XI0_20/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN0_10 XI11_3/net21_5_ xsel_20_ XI11_3/XI0/XI0_20/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN0_9 XI11_3/net21_6_ xsel_20_ XI11_3/XI0/XI0_20/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN0_8 XI11_3/net21_7_ xsel_20_ XI11_3/XI0/XI0_20/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN0_7 XI11_3/net21_8_ xsel_20_ XI11_3/XI0/XI0_20/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN0_6 XI11_3/net21_9_ xsel_20_ XI11_3/XI0/XI0_20/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN0_5 XI11_3/net21_10_ xsel_20_ XI11_3/XI0/XI0_20/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN0_4 XI11_3/net21_11_ xsel_20_ XI11_3/XI0/XI0_20/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN0_3 XI11_3/net21_12_ xsel_20_ XI11_3/XI0/XI0_20/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN0_2 XI11_3/net21_13_ xsel_20_ XI11_3/XI0/XI0_20/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN0_1 XI11_3/net21_14_ xsel_20_ XI11_3/XI0/XI0_20/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN0_0 XI11_3/net21_15_ xsel_20_ XI11_3/XI0/XI0_20/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN1_15 XI11_3/XI0/XI0_20/d__15_ xsel_20_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN1_14 XI11_3/XI0/XI0_20/d__14_ xsel_20_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN1_13 XI11_3/XI0/XI0_20/d__13_ xsel_20_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN1_12 XI11_3/XI0/XI0_20/d__12_ xsel_20_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN1_11 XI11_3/XI0/XI0_20/d__11_ xsel_20_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN1_10 XI11_3/XI0/XI0_20/d__10_ xsel_20_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN1_9 XI11_3/XI0/XI0_20/d__9_ xsel_20_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN1_8 XI11_3/XI0/XI0_20/d__8_ xsel_20_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN1_7 XI11_3/XI0/XI0_20/d__7_ xsel_20_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN1_6 XI11_3/XI0/XI0_20/d__6_ xsel_20_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN1_5 XI11_3/XI0/XI0_20/d__5_ xsel_20_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN1_4 XI11_3/XI0/XI0_20/d__4_ xsel_20_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN1_3 XI11_3/XI0/XI0_20/d__3_ xsel_20_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN1_2 XI11_3/XI0/XI0_20/d__2_ xsel_20_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN1_1 XI11_3/XI0/XI0_20/d__1_ xsel_20_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_20/MN1_0 XI11_3/XI0/XI0_20/d__0_ xsel_20_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN0_15 XI11_3/net21_0_ xsel_19_ XI11_3/XI0/XI0_19/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN0_14 XI11_3/net21_1_ xsel_19_ XI11_3/XI0/XI0_19/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN0_13 XI11_3/net21_2_ xsel_19_ XI11_3/XI0/XI0_19/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN0_12 XI11_3/net21_3_ xsel_19_ XI11_3/XI0/XI0_19/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN0_11 XI11_3/net21_4_ xsel_19_ XI11_3/XI0/XI0_19/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN0_10 XI11_3/net21_5_ xsel_19_ XI11_3/XI0/XI0_19/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN0_9 XI11_3/net21_6_ xsel_19_ XI11_3/XI0/XI0_19/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN0_8 XI11_3/net21_7_ xsel_19_ XI11_3/XI0/XI0_19/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN0_7 XI11_3/net21_8_ xsel_19_ XI11_3/XI0/XI0_19/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN0_6 XI11_3/net21_9_ xsel_19_ XI11_3/XI0/XI0_19/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN0_5 XI11_3/net21_10_ xsel_19_ XI11_3/XI0/XI0_19/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN0_4 XI11_3/net21_11_ xsel_19_ XI11_3/XI0/XI0_19/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN0_3 XI11_3/net21_12_ xsel_19_ XI11_3/XI0/XI0_19/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN0_2 XI11_3/net21_13_ xsel_19_ XI11_3/XI0/XI0_19/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN0_1 XI11_3/net21_14_ xsel_19_ XI11_3/XI0/XI0_19/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN0_0 XI11_3/net21_15_ xsel_19_ XI11_3/XI0/XI0_19/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN1_15 XI11_3/XI0/XI0_19/d__15_ xsel_19_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN1_14 XI11_3/XI0/XI0_19/d__14_ xsel_19_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN1_13 XI11_3/XI0/XI0_19/d__13_ xsel_19_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN1_12 XI11_3/XI0/XI0_19/d__12_ xsel_19_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN1_11 XI11_3/XI0/XI0_19/d__11_ xsel_19_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN1_10 XI11_3/XI0/XI0_19/d__10_ xsel_19_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN1_9 XI11_3/XI0/XI0_19/d__9_ xsel_19_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN1_8 XI11_3/XI0/XI0_19/d__8_ xsel_19_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN1_7 XI11_3/XI0/XI0_19/d__7_ xsel_19_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN1_6 XI11_3/XI0/XI0_19/d__6_ xsel_19_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN1_5 XI11_3/XI0/XI0_19/d__5_ xsel_19_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN1_4 XI11_3/XI0/XI0_19/d__4_ xsel_19_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN1_3 XI11_3/XI0/XI0_19/d__3_ xsel_19_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN1_2 XI11_3/XI0/XI0_19/d__2_ xsel_19_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN1_1 XI11_3/XI0/XI0_19/d__1_ xsel_19_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_19/MN1_0 XI11_3/XI0/XI0_19/d__0_ xsel_19_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN0_15 XI11_3/net21_0_ xsel_18_ XI11_3/XI0/XI0_18/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN0_14 XI11_3/net21_1_ xsel_18_ XI11_3/XI0/XI0_18/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN0_13 XI11_3/net21_2_ xsel_18_ XI11_3/XI0/XI0_18/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN0_12 XI11_3/net21_3_ xsel_18_ XI11_3/XI0/XI0_18/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN0_11 XI11_3/net21_4_ xsel_18_ XI11_3/XI0/XI0_18/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN0_10 XI11_3/net21_5_ xsel_18_ XI11_3/XI0/XI0_18/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN0_9 XI11_3/net21_6_ xsel_18_ XI11_3/XI0/XI0_18/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN0_8 XI11_3/net21_7_ xsel_18_ XI11_3/XI0/XI0_18/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN0_7 XI11_3/net21_8_ xsel_18_ XI11_3/XI0/XI0_18/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN0_6 XI11_3/net21_9_ xsel_18_ XI11_3/XI0/XI0_18/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN0_5 XI11_3/net21_10_ xsel_18_ XI11_3/XI0/XI0_18/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN0_4 XI11_3/net21_11_ xsel_18_ XI11_3/XI0/XI0_18/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN0_3 XI11_3/net21_12_ xsel_18_ XI11_3/XI0/XI0_18/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN0_2 XI11_3/net21_13_ xsel_18_ XI11_3/XI0/XI0_18/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN0_1 XI11_3/net21_14_ xsel_18_ XI11_3/XI0/XI0_18/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN0_0 XI11_3/net21_15_ xsel_18_ XI11_3/XI0/XI0_18/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN1_15 XI11_3/XI0/XI0_18/d__15_ xsel_18_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN1_14 XI11_3/XI0/XI0_18/d__14_ xsel_18_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN1_13 XI11_3/XI0/XI0_18/d__13_ xsel_18_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN1_12 XI11_3/XI0/XI0_18/d__12_ xsel_18_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN1_11 XI11_3/XI0/XI0_18/d__11_ xsel_18_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN1_10 XI11_3/XI0/XI0_18/d__10_ xsel_18_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN1_9 XI11_3/XI0/XI0_18/d__9_ xsel_18_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN1_8 XI11_3/XI0/XI0_18/d__8_ xsel_18_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN1_7 XI11_3/XI0/XI0_18/d__7_ xsel_18_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN1_6 XI11_3/XI0/XI0_18/d__6_ xsel_18_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN1_5 XI11_3/XI0/XI0_18/d__5_ xsel_18_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN1_4 XI11_3/XI0/XI0_18/d__4_ xsel_18_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN1_3 XI11_3/XI0/XI0_18/d__3_ xsel_18_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN1_2 XI11_3/XI0/XI0_18/d__2_ xsel_18_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN1_1 XI11_3/XI0/XI0_18/d__1_ xsel_18_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_18/MN1_0 XI11_3/XI0/XI0_18/d__0_ xsel_18_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN0_15 XI11_3/net21_0_ xsel_17_ XI11_3/XI0/XI0_17/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN0_14 XI11_3/net21_1_ xsel_17_ XI11_3/XI0/XI0_17/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN0_13 XI11_3/net21_2_ xsel_17_ XI11_3/XI0/XI0_17/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN0_12 XI11_3/net21_3_ xsel_17_ XI11_3/XI0/XI0_17/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN0_11 XI11_3/net21_4_ xsel_17_ XI11_3/XI0/XI0_17/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN0_10 XI11_3/net21_5_ xsel_17_ XI11_3/XI0/XI0_17/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN0_9 XI11_3/net21_6_ xsel_17_ XI11_3/XI0/XI0_17/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN0_8 XI11_3/net21_7_ xsel_17_ XI11_3/XI0/XI0_17/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN0_7 XI11_3/net21_8_ xsel_17_ XI11_3/XI0/XI0_17/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN0_6 XI11_3/net21_9_ xsel_17_ XI11_3/XI0/XI0_17/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN0_5 XI11_3/net21_10_ xsel_17_ XI11_3/XI0/XI0_17/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN0_4 XI11_3/net21_11_ xsel_17_ XI11_3/XI0/XI0_17/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN0_3 XI11_3/net21_12_ xsel_17_ XI11_3/XI0/XI0_17/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN0_2 XI11_3/net21_13_ xsel_17_ XI11_3/XI0/XI0_17/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN0_1 XI11_3/net21_14_ xsel_17_ XI11_3/XI0/XI0_17/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN0_0 XI11_3/net21_15_ xsel_17_ XI11_3/XI0/XI0_17/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN1_15 XI11_3/XI0/XI0_17/d__15_ xsel_17_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN1_14 XI11_3/XI0/XI0_17/d__14_ xsel_17_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN1_13 XI11_3/XI0/XI0_17/d__13_ xsel_17_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN1_12 XI11_3/XI0/XI0_17/d__12_ xsel_17_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN1_11 XI11_3/XI0/XI0_17/d__11_ xsel_17_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN1_10 XI11_3/XI0/XI0_17/d__10_ xsel_17_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN1_9 XI11_3/XI0/XI0_17/d__9_ xsel_17_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN1_8 XI11_3/XI0/XI0_17/d__8_ xsel_17_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN1_7 XI11_3/XI0/XI0_17/d__7_ xsel_17_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN1_6 XI11_3/XI0/XI0_17/d__6_ xsel_17_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN1_5 XI11_3/XI0/XI0_17/d__5_ xsel_17_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN1_4 XI11_3/XI0/XI0_17/d__4_ xsel_17_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN1_3 XI11_3/XI0/XI0_17/d__3_ xsel_17_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN1_2 XI11_3/XI0/XI0_17/d__2_ xsel_17_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN1_1 XI11_3/XI0/XI0_17/d__1_ xsel_17_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_17/MN1_0 XI11_3/XI0/XI0_17/d__0_ xsel_17_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN0_15 XI11_3/net21_0_ xsel_16_ XI11_3/XI0/XI0_16/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN0_14 XI11_3/net21_1_ xsel_16_ XI11_3/XI0/XI0_16/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN0_13 XI11_3/net21_2_ xsel_16_ XI11_3/XI0/XI0_16/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN0_12 XI11_3/net21_3_ xsel_16_ XI11_3/XI0/XI0_16/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN0_11 XI11_3/net21_4_ xsel_16_ XI11_3/XI0/XI0_16/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN0_10 XI11_3/net21_5_ xsel_16_ XI11_3/XI0/XI0_16/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN0_9 XI11_3/net21_6_ xsel_16_ XI11_3/XI0/XI0_16/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN0_8 XI11_3/net21_7_ xsel_16_ XI11_3/XI0/XI0_16/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN0_7 XI11_3/net21_8_ xsel_16_ XI11_3/XI0/XI0_16/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN0_6 XI11_3/net21_9_ xsel_16_ XI11_3/XI0/XI0_16/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN0_5 XI11_3/net21_10_ xsel_16_ XI11_3/XI0/XI0_16/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN0_4 XI11_3/net21_11_ xsel_16_ XI11_3/XI0/XI0_16/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN0_3 XI11_3/net21_12_ xsel_16_ XI11_3/XI0/XI0_16/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN0_2 XI11_3/net21_13_ xsel_16_ XI11_3/XI0/XI0_16/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN0_1 XI11_3/net21_14_ xsel_16_ XI11_3/XI0/XI0_16/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN0_0 XI11_3/net21_15_ xsel_16_ XI11_3/XI0/XI0_16/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN1_15 XI11_3/XI0/XI0_16/d__15_ xsel_16_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN1_14 XI11_3/XI0/XI0_16/d__14_ xsel_16_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN1_13 XI11_3/XI0/XI0_16/d__13_ xsel_16_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN1_12 XI11_3/XI0/XI0_16/d__12_ xsel_16_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN1_11 XI11_3/XI0/XI0_16/d__11_ xsel_16_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN1_10 XI11_3/XI0/XI0_16/d__10_ xsel_16_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN1_9 XI11_3/XI0/XI0_16/d__9_ xsel_16_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN1_8 XI11_3/XI0/XI0_16/d__8_ xsel_16_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN1_7 XI11_3/XI0/XI0_16/d__7_ xsel_16_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN1_6 XI11_3/XI0/XI0_16/d__6_ xsel_16_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN1_5 XI11_3/XI0/XI0_16/d__5_ xsel_16_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN1_4 XI11_3/XI0/XI0_16/d__4_ xsel_16_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN1_3 XI11_3/XI0/XI0_16/d__3_ xsel_16_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN1_2 XI11_3/XI0/XI0_16/d__2_ xsel_16_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN1_1 XI11_3/XI0/XI0_16/d__1_ xsel_16_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_16/MN1_0 XI11_3/XI0/XI0_16/d__0_ xsel_16_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN0_15 XI11_3/net21_0_ xsel_15_ XI11_3/XI0/XI0_15/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN0_14 XI11_3/net21_1_ xsel_15_ XI11_3/XI0/XI0_15/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN0_13 XI11_3/net21_2_ xsel_15_ XI11_3/XI0/XI0_15/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN0_12 XI11_3/net21_3_ xsel_15_ XI11_3/XI0/XI0_15/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN0_11 XI11_3/net21_4_ xsel_15_ XI11_3/XI0/XI0_15/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN0_10 XI11_3/net21_5_ xsel_15_ XI11_3/XI0/XI0_15/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN0_9 XI11_3/net21_6_ xsel_15_ XI11_3/XI0/XI0_15/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN0_8 XI11_3/net21_7_ xsel_15_ XI11_3/XI0/XI0_15/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN0_7 XI11_3/net21_8_ xsel_15_ XI11_3/XI0/XI0_15/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN0_6 XI11_3/net21_9_ xsel_15_ XI11_3/XI0/XI0_15/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN0_5 XI11_3/net21_10_ xsel_15_ XI11_3/XI0/XI0_15/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN0_4 XI11_3/net21_11_ xsel_15_ XI11_3/XI0/XI0_15/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN0_3 XI11_3/net21_12_ xsel_15_ XI11_3/XI0/XI0_15/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN0_2 XI11_3/net21_13_ xsel_15_ XI11_3/XI0/XI0_15/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN0_1 XI11_3/net21_14_ xsel_15_ XI11_3/XI0/XI0_15/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN0_0 XI11_3/net21_15_ xsel_15_ XI11_3/XI0/XI0_15/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN1_15 XI11_3/XI0/XI0_15/d__15_ xsel_15_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN1_14 XI11_3/XI0/XI0_15/d__14_ xsel_15_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN1_13 XI11_3/XI0/XI0_15/d__13_ xsel_15_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN1_12 XI11_3/XI0/XI0_15/d__12_ xsel_15_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN1_11 XI11_3/XI0/XI0_15/d__11_ xsel_15_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN1_10 XI11_3/XI0/XI0_15/d__10_ xsel_15_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN1_9 XI11_3/XI0/XI0_15/d__9_ xsel_15_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN1_8 XI11_3/XI0/XI0_15/d__8_ xsel_15_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN1_7 XI11_3/XI0/XI0_15/d__7_ xsel_15_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN1_6 XI11_3/XI0/XI0_15/d__6_ xsel_15_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN1_5 XI11_3/XI0/XI0_15/d__5_ xsel_15_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN1_4 XI11_3/XI0/XI0_15/d__4_ xsel_15_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN1_3 XI11_3/XI0/XI0_15/d__3_ xsel_15_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN1_2 XI11_3/XI0/XI0_15/d__2_ xsel_15_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN1_1 XI11_3/XI0/XI0_15/d__1_ xsel_15_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_15/MN1_0 XI11_3/XI0/XI0_15/d__0_ xsel_15_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN0_15 XI11_3/net21_0_ xsel_14_ XI11_3/XI0/XI0_14/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN0_14 XI11_3/net21_1_ xsel_14_ XI11_3/XI0/XI0_14/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN0_13 XI11_3/net21_2_ xsel_14_ XI11_3/XI0/XI0_14/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN0_12 XI11_3/net21_3_ xsel_14_ XI11_3/XI0/XI0_14/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN0_11 XI11_3/net21_4_ xsel_14_ XI11_3/XI0/XI0_14/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN0_10 XI11_3/net21_5_ xsel_14_ XI11_3/XI0/XI0_14/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN0_9 XI11_3/net21_6_ xsel_14_ XI11_3/XI0/XI0_14/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN0_8 XI11_3/net21_7_ xsel_14_ XI11_3/XI0/XI0_14/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN0_7 XI11_3/net21_8_ xsel_14_ XI11_3/XI0/XI0_14/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN0_6 XI11_3/net21_9_ xsel_14_ XI11_3/XI0/XI0_14/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN0_5 XI11_3/net21_10_ xsel_14_ XI11_3/XI0/XI0_14/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN0_4 XI11_3/net21_11_ xsel_14_ XI11_3/XI0/XI0_14/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN0_3 XI11_3/net21_12_ xsel_14_ XI11_3/XI0/XI0_14/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN0_2 XI11_3/net21_13_ xsel_14_ XI11_3/XI0/XI0_14/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN0_1 XI11_3/net21_14_ xsel_14_ XI11_3/XI0/XI0_14/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN0_0 XI11_3/net21_15_ xsel_14_ XI11_3/XI0/XI0_14/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN1_15 XI11_3/XI0/XI0_14/d__15_ xsel_14_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN1_14 XI11_3/XI0/XI0_14/d__14_ xsel_14_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN1_13 XI11_3/XI0/XI0_14/d__13_ xsel_14_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN1_12 XI11_3/XI0/XI0_14/d__12_ xsel_14_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN1_11 XI11_3/XI0/XI0_14/d__11_ xsel_14_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN1_10 XI11_3/XI0/XI0_14/d__10_ xsel_14_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN1_9 XI11_3/XI0/XI0_14/d__9_ xsel_14_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN1_8 XI11_3/XI0/XI0_14/d__8_ xsel_14_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN1_7 XI11_3/XI0/XI0_14/d__7_ xsel_14_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN1_6 XI11_3/XI0/XI0_14/d__6_ xsel_14_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN1_5 XI11_3/XI0/XI0_14/d__5_ xsel_14_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN1_4 XI11_3/XI0/XI0_14/d__4_ xsel_14_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN1_3 XI11_3/XI0/XI0_14/d__3_ xsel_14_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN1_2 XI11_3/XI0/XI0_14/d__2_ xsel_14_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN1_1 XI11_3/XI0/XI0_14/d__1_ xsel_14_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_14/MN1_0 XI11_3/XI0/XI0_14/d__0_ xsel_14_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN0_15 XI11_3/net21_0_ xsel_13_ XI11_3/XI0/XI0_13/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN0_14 XI11_3/net21_1_ xsel_13_ XI11_3/XI0/XI0_13/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN0_13 XI11_3/net21_2_ xsel_13_ XI11_3/XI0/XI0_13/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN0_12 XI11_3/net21_3_ xsel_13_ XI11_3/XI0/XI0_13/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN0_11 XI11_3/net21_4_ xsel_13_ XI11_3/XI0/XI0_13/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN0_10 XI11_3/net21_5_ xsel_13_ XI11_3/XI0/XI0_13/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN0_9 XI11_3/net21_6_ xsel_13_ XI11_3/XI0/XI0_13/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN0_8 XI11_3/net21_7_ xsel_13_ XI11_3/XI0/XI0_13/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN0_7 XI11_3/net21_8_ xsel_13_ XI11_3/XI0/XI0_13/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN0_6 XI11_3/net21_9_ xsel_13_ XI11_3/XI0/XI0_13/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN0_5 XI11_3/net21_10_ xsel_13_ XI11_3/XI0/XI0_13/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN0_4 XI11_3/net21_11_ xsel_13_ XI11_3/XI0/XI0_13/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN0_3 XI11_3/net21_12_ xsel_13_ XI11_3/XI0/XI0_13/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN0_2 XI11_3/net21_13_ xsel_13_ XI11_3/XI0/XI0_13/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN0_1 XI11_3/net21_14_ xsel_13_ XI11_3/XI0/XI0_13/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN0_0 XI11_3/net21_15_ xsel_13_ XI11_3/XI0/XI0_13/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN1_15 XI11_3/XI0/XI0_13/d__15_ xsel_13_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN1_14 XI11_3/XI0/XI0_13/d__14_ xsel_13_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN1_13 XI11_3/XI0/XI0_13/d__13_ xsel_13_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN1_12 XI11_3/XI0/XI0_13/d__12_ xsel_13_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN1_11 XI11_3/XI0/XI0_13/d__11_ xsel_13_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN1_10 XI11_3/XI0/XI0_13/d__10_ xsel_13_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN1_9 XI11_3/XI0/XI0_13/d__9_ xsel_13_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN1_8 XI11_3/XI0/XI0_13/d__8_ xsel_13_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN1_7 XI11_3/XI0/XI0_13/d__7_ xsel_13_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN1_6 XI11_3/XI0/XI0_13/d__6_ xsel_13_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN1_5 XI11_3/XI0/XI0_13/d__5_ xsel_13_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN1_4 XI11_3/XI0/XI0_13/d__4_ xsel_13_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN1_3 XI11_3/XI0/XI0_13/d__3_ xsel_13_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN1_2 XI11_3/XI0/XI0_13/d__2_ xsel_13_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN1_1 XI11_3/XI0/XI0_13/d__1_ xsel_13_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_13/MN1_0 XI11_3/XI0/XI0_13/d__0_ xsel_13_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN0_15 XI11_3/net21_0_ xsel_12_ XI11_3/XI0/XI0_12/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN0_14 XI11_3/net21_1_ xsel_12_ XI11_3/XI0/XI0_12/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN0_13 XI11_3/net21_2_ xsel_12_ XI11_3/XI0/XI0_12/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN0_12 XI11_3/net21_3_ xsel_12_ XI11_3/XI0/XI0_12/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN0_11 XI11_3/net21_4_ xsel_12_ XI11_3/XI0/XI0_12/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN0_10 XI11_3/net21_5_ xsel_12_ XI11_3/XI0/XI0_12/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN0_9 XI11_3/net21_6_ xsel_12_ XI11_3/XI0/XI0_12/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN0_8 XI11_3/net21_7_ xsel_12_ XI11_3/XI0/XI0_12/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN0_7 XI11_3/net21_8_ xsel_12_ XI11_3/XI0/XI0_12/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN0_6 XI11_3/net21_9_ xsel_12_ XI11_3/XI0/XI0_12/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN0_5 XI11_3/net21_10_ xsel_12_ XI11_3/XI0/XI0_12/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN0_4 XI11_3/net21_11_ xsel_12_ XI11_3/XI0/XI0_12/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN0_3 XI11_3/net21_12_ xsel_12_ XI11_3/XI0/XI0_12/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN0_2 XI11_3/net21_13_ xsel_12_ XI11_3/XI0/XI0_12/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN0_1 XI11_3/net21_14_ xsel_12_ XI11_3/XI0/XI0_12/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN0_0 XI11_3/net21_15_ xsel_12_ XI11_3/XI0/XI0_12/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN1_15 XI11_3/XI0/XI0_12/d__15_ xsel_12_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN1_14 XI11_3/XI0/XI0_12/d__14_ xsel_12_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN1_13 XI11_3/XI0/XI0_12/d__13_ xsel_12_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN1_12 XI11_3/XI0/XI0_12/d__12_ xsel_12_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN1_11 XI11_3/XI0/XI0_12/d__11_ xsel_12_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN1_10 XI11_3/XI0/XI0_12/d__10_ xsel_12_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN1_9 XI11_3/XI0/XI0_12/d__9_ xsel_12_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN1_8 XI11_3/XI0/XI0_12/d__8_ xsel_12_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN1_7 XI11_3/XI0/XI0_12/d__7_ xsel_12_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN1_6 XI11_3/XI0/XI0_12/d__6_ xsel_12_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN1_5 XI11_3/XI0/XI0_12/d__5_ xsel_12_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN1_4 XI11_3/XI0/XI0_12/d__4_ xsel_12_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN1_3 XI11_3/XI0/XI0_12/d__3_ xsel_12_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN1_2 XI11_3/XI0/XI0_12/d__2_ xsel_12_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN1_1 XI11_3/XI0/XI0_12/d__1_ xsel_12_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_12/MN1_0 XI11_3/XI0/XI0_12/d__0_ xsel_12_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN0_15 XI11_3/net21_0_ xsel_11_ XI11_3/XI0/XI0_11/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN0_14 XI11_3/net21_1_ xsel_11_ XI11_3/XI0/XI0_11/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN0_13 XI11_3/net21_2_ xsel_11_ XI11_3/XI0/XI0_11/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN0_12 XI11_3/net21_3_ xsel_11_ XI11_3/XI0/XI0_11/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN0_11 XI11_3/net21_4_ xsel_11_ XI11_3/XI0/XI0_11/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN0_10 XI11_3/net21_5_ xsel_11_ XI11_3/XI0/XI0_11/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN0_9 XI11_3/net21_6_ xsel_11_ XI11_3/XI0/XI0_11/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN0_8 XI11_3/net21_7_ xsel_11_ XI11_3/XI0/XI0_11/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN0_7 XI11_3/net21_8_ xsel_11_ XI11_3/XI0/XI0_11/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN0_6 XI11_3/net21_9_ xsel_11_ XI11_3/XI0/XI0_11/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN0_5 XI11_3/net21_10_ xsel_11_ XI11_3/XI0/XI0_11/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN0_4 XI11_3/net21_11_ xsel_11_ XI11_3/XI0/XI0_11/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN0_3 XI11_3/net21_12_ xsel_11_ XI11_3/XI0/XI0_11/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN0_2 XI11_3/net21_13_ xsel_11_ XI11_3/XI0/XI0_11/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN0_1 XI11_3/net21_14_ xsel_11_ XI11_3/XI0/XI0_11/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN0_0 XI11_3/net21_15_ xsel_11_ XI11_3/XI0/XI0_11/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN1_15 XI11_3/XI0/XI0_11/d__15_ xsel_11_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN1_14 XI11_3/XI0/XI0_11/d__14_ xsel_11_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN1_13 XI11_3/XI0/XI0_11/d__13_ xsel_11_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN1_12 XI11_3/XI0/XI0_11/d__12_ xsel_11_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN1_11 XI11_3/XI0/XI0_11/d__11_ xsel_11_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN1_10 XI11_3/XI0/XI0_11/d__10_ xsel_11_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN1_9 XI11_3/XI0/XI0_11/d__9_ xsel_11_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN1_8 XI11_3/XI0/XI0_11/d__8_ xsel_11_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN1_7 XI11_3/XI0/XI0_11/d__7_ xsel_11_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN1_6 XI11_3/XI0/XI0_11/d__6_ xsel_11_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN1_5 XI11_3/XI0/XI0_11/d__5_ xsel_11_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN1_4 XI11_3/XI0/XI0_11/d__4_ xsel_11_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN1_3 XI11_3/XI0/XI0_11/d__3_ xsel_11_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN1_2 XI11_3/XI0/XI0_11/d__2_ xsel_11_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN1_1 XI11_3/XI0/XI0_11/d__1_ xsel_11_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_11/MN1_0 XI11_3/XI0/XI0_11/d__0_ xsel_11_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN0_15 XI11_3/net21_0_ xsel_10_ XI11_3/XI0/XI0_10/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN0_14 XI11_3/net21_1_ xsel_10_ XI11_3/XI0/XI0_10/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN0_13 XI11_3/net21_2_ xsel_10_ XI11_3/XI0/XI0_10/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN0_12 XI11_3/net21_3_ xsel_10_ XI11_3/XI0/XI0_10/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN0_11 XI11_3/net21_4_ xsel_10_ XI11_3/XI0/XI0_10/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN0_10 XI11_3/net21_5_ xsel_10_ XI11_3/XI0/XI0_10/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN0_9 XI11_3/net21_6_ xsel_10_ XI11_3/XI0/XI0_10/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN0_8 XI11_3/net21_7_ xsel_10_ XI11_3/XI0/XI0_10/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN0_7 XI11_3/net21_8_ xsel_10_ XI11_3/XI0/XI0_10/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN0_6 XI11_3/net21_9_ xsel_10_ XI11_3/XI0/XI0_10/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN0_5 XI11_3/net21_10_ xsel_10_ XI11_3/XI0/XI0_10/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN0_4 XI11_3/net21_11_ xsel_10_ XI11_3/XI0/XI0_10/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN0_3 XI11_3/net21_12_ xsel_10_ XI11_3/XI0/XI0_10/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN0_2 XI11_3/net21_13_ xsel_10_ XI11_3/XI0/XI0_10/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN0_1 XI11_3/net21_14_ xsel_10_ XI11_3/XI0/XI0_10/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN0_0 XI11_3/net21_15_ xsel_10_ XI11_3/XI0/XI0_10/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN1_15 XI11_3/XI0/XI0_10/d__15_ xsel_10_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN1_14 XI11_3/XI0/XI0_10/d__14_ xsel_10_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN1_13 XI11_3/XI0/XI0_10/d__13_ xsel_10_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN1_12 XI11_3/XI0/XI0_10/d__12_ xsel_10_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN1_11 XI11_3/XI0/XI0_10/d__11_ xsel_10_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN1_10 XI11_3/XI0/XI0_10/d__10_ xsel_10_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN1_9 XI11_3/XI0/XI0_10/d__9_ xsel_10_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN1_8 XI11_3/XI0/XI0_10/d__8_ xsel_10_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN1_7 XI11_3/XI0/XI0_10/d__7_ xsel_10_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN1_6 XI11_3/XI0/XI0_10/d__6_ xsel_10_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN1_5 XI11_3/XI0/XI0_10/d__5_ xsel_10_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN1_4 XI11_3/XI0/XI0_10/d__4_ xsel_10_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN1_3 XI11_3/XI0/XI0_10/d__3_ xsel_10_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN1_2 XI11_3/XI0/XI0_10/d__2_ xsel_10_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN1_1 XI11_3/XI0/XI0_10/d__1_ xsel_10_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_10/MN1_0 XI11_3/XI0/XI0_10/d__0_ xsel_10_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN0_15 XI11_3/net21_0_ xsel_9_ XI11_3/XI0/XI0_9/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN0_14 XI11_3/net21_1_ xsel_9_ XI11_3/XI0/XI0_9/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN0_13 XI11_3/net21_2_ xsel_9_ XI11_3/XI0/XI0_9/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN0_12 XI11_3/net21_3_ xsel_9_ XI11_3/XI0/XI0_9/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN0_11 XI11_3/net21_4_ xsel_9_ XI11_3/XI0/XI0_9/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN0_10 XI11_3/net21_5_ xsel_9_ XI11_3/XI0/XI0_9/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN0_9 XI11_3/net21_6_ xsel_9_ XI11_3/XI0/XI0_9/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN0_8 XI11_3/net21_7_ xsel_9_ XI11_3/XI0/XI0_9/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN0_7 XI11_3/net21_8_ xsel_9_ XI11_3/XI0/XI0_9/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN0_6 XI11_3/net21_9_ xsel_9_ XI11_3/XI0/XI0_9/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN0_5 XI11_3/net21_10_ xsel_9_ XI11_3/XI0/XI0_9/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN0_4 XI11_3/net21_11_ xsel_9_ XI11_3/XI0/XI0_9/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN0_3 XI11_3/net21_12_ xsel_9_ XI11_3/XI0/XI0_9/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN0_2 XI11_3/net21_13_ xsel_9_ XI11_3/XI0/XI0_9/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN0_1 XI11_3/net21_14_ xsel_9_ XI11_3/XI0/XI0_9/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN0_0 XI11_3/net21_15_ xsel_9_ XI11_3/XI0/XI0_9/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN1_15 XI11_3/XI0/XI0_9/d__15_ xsel_9_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN1_14 XI11_3/XI0/XI0_9/d__14_ xsel_9_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN1_13 XI11_3/XI0/XI0_9/d__13_ xsel_9_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN1_12 XI11_3/XI0/XI0_9/d__12_ xsel_9_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN1_11 XI11_3/XI0/XI0_9/d__11_ xsel_9_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN1_10 XI11_3/XI0/XI0_9/d__10_ xsel_9_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN1_9 XI11_3/XI0/XI0_9/d__9_ xsel_9_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN1_8 XI11_3/XI0/XI0_9/d__8_ xsel_9_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN1_7 XI11_3/XI0/XI0_9/d__7_ xsel_9_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN1_6 XI11_3/XI0/XI0_9/d__6_ xsel_9_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN1_5 XI11_3/XI0/XI0_9/d__5_ xsel_9_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN1_4 XI11_3/XI0/XI0_9/d__4_ xsel_9_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN1_3 XI11_3/XI0/XI0_9/d__3_ xsel_9_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN1_2 XI11_3/XI0/XI0_9/d__2_ xsel_9_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN1_1 XI11_3/XI0/XI0_9/d__1_ xsel_9_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_9/MN1_0 XI11_3/XI0/XI0_9/d__0_ xsel_9_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN0_15 XI11_3/net21_0_ xsel_8_ XI11_3/XI0/XI0_8/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN0_14 XI11_3/net21_1_ xsel_8_ XI11_3/XI0/XI0_8/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN0_13 XI11_3/net21_2_ xsel_8_ XI11_3/XI0/XI0_8/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN0_12 XI11_3/net21_3_ xsel_8_ XI11_3/XI0/XI0_8/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN0_11 XI11_3/net21_4_ xsel_8_ XI11_3/XI0/XI0_8/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN0_10 XI11_3/net21_5_ xsel_8_ XI11_3/XI0/XI0_8/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN0_9 XI11_3/net21_6_ xsel_8_ XI11_3/XI0/XI0_8/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN0_8 XI11_3/net21_7_ xsel_8_ XI11_3/XI0/XI0_8/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN0_7 XI11_3/net21_8_ xsel_8_ XI11_3/XI0/XI0_8/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN0_6 XI11_3/net21_9_ xsel_8_ XI11_3/XI0/XI0_8/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN0_5 XI11_3/net21_10_ xsel_8_ XI11_3/XI0/XI0_8/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN0_4 XI11_3/net21_11_ xsel_8_ XI11_3/XI0/XI0_8/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN0_3 XI11_3/net21_12_ xsel_8_ XI11_3/XI0/XI0_8/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN0_2 XI11_3/net21_13_ xsel_8_ XI11_3/XI0/XI0_8/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN0_1 XI11_3/net21_14_ xsel_8_ XI11_3/XI0/XI0_8/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN0_0 XI11_3/net21_15_ xsel_8_ XI11_3/XI0/XI0_8/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN1_15 XI11_3/XI0/XI0_8/d__15_ xsel_8_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN1_14 XI11_3/XI0/XI0_8/d__14_ xsel_8_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN1_13 XI11_3/XI0/XI0_8/d__13_ xsel_8_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN1_12 XI11_3/XI0/XI0_8/d__12_ xsel_8_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN1_11 XI11_3/XI0/XI0_8/d__11_ xsel_8_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN1_10 XI11_3/XI0/XI0_8/d__10_ xsel_8_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN1_9 XI11_3/XI0/XI0_8/d__9_ xsel_8_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN1_8 XI11_3/XI0/XI0_8/d__8_ xsel_8_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN1_7 XI11_3/XI0/XI0_8/d__7_ xsel_8_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN1_6 XI11_3/XI0/XI0_8/d__6_ xsel_8_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN1_5 XI11_3/XI0/XI0_8/d__5_ xsel_8_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN1_4 XI11_3/XI0/XI0_8/d__4_ xsel_8_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN1_3 XI11_3/XI0/XI0_8/d__3_ xsel_8_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN1_2 XI11_3/XI0/XI0_8/d__2_ xsel_8_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN1_1 XI11_3/XI0/XI0_8/d__1_ xsel_8_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_8/MN1_0 XI11_3/XI0/XI0_8/d__0_ xsel_8_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN0_15 XI11_3/net21_0_ xsel_7_ XI11_3/XI0/XI0_7/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN0_14 XI11_3/net21_1_ xsel_7_ XI11_3/XI0/XI0_7/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN0_13 XI11_3/net21_2_ xsel_7_ XI11_3/XI0/XI0_7/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN0_12 XI11_3/net21_3_ xsel_7_ XI11_3/XI0/XI0_7/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN0_11 XI11_3/net21_4_ xsel_7_ XI11_3/XI0/XI0_7/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN0_10 XI11_3/net21_5_ xsel_7_ XI11_3/XI0/XI0_7/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN0_9 XI11_3/net21_6_ xsel_7_ XI11_3/XI0/XI0_7/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN0_8 XI11_3/net21_7_ xsel_7_ XI11_3/XI0/XI0_7/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN0_7 XI11_3/net21_8_ xsel_7_ XI11_3/XI0/XI0_7/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN0_6 XI11_3/net21_9_ xsel_7_ XI11_3/XI0/XI0_7/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN0_5 XI11_3/net21_10_ xsel_7_ XI11_3/XI0/XI0_7/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN0_4 XI11_3/net21_11_ xsel_7_ XI11_3/XI0/XI0_7/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN0_3 XI11_3/net21_12_ xsel_7_ XI11_3/XI0/XI0_7/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN0_2 XI11_3/net21_13_ xsel_7_ XI11_3/XI0/XI0_7/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN0_1 XI11_3/net21_14_ xsel_7_ XI11_3/XI0/XI0_7/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN0_0 XI11_3/net21_15_ xsel_7_ XI11_3/XI0/XI0_7/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN1_15 XI11_3/XI0/XI0_7/d__15_ xsel_7_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN1_14 XI11_3/XI0/XI0_7/d__14_ xsel_7_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN1_13 XI11_3/XI0/XI0_7/d__13_ xsel_7_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN1_12 XI11_3/XI0/XI0_7/d__12_ xsel_7_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN1_11 XI11_3/XI0/XI0_7/d__11_ xsel_7_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN1_10 XI11_3/XI0/XI0_7/d__10_ xsel_7_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN1_9 XI11_3/XI0/XI0_7/d__9_ xsel_7_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN1_8 XI11_3/XI0/XI0_7/d__8_ xsel_7_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN1_7 XI11_3/XI0/XI0_7/d__7_ xsel_7_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN1_6 XI11_3/XI0/XI0_7/d__6_ xsel_7_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN1_5 XI11_3/XI0/XI0_7/d__5_ xsel_7_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN1_4 XI11_3/XI0/XI0_7/d__4_ xsel_7_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN1_3 XI11_3/XI0/XI0_7/d__3_ xsel_7_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN1_2 XI11_3/XI0/XI0_7/d__2_ xsel_7_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN1_1 XI11_3/XI0/XI0_7/d__1_ xsel_7_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_7/MN1_0 XI11_3/XI0/XI0_7/d__0_ xsel_7_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN0_15 XI11_3/net21_0_ xsel_6_ XI11_3/XI0/XI0_6/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN0_14 XI11_3/net21_1_ xsel_6_ XI11_3/XI0/XI0_6/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN0_13 XI11_3/net21_2_ xsel_6_ XI11_3/XI0/XI0_6/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN0_12 XI11_3/net21_3_ xsel_6_ XI11_3/XI0/XI0_6/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN0_11 XI11_3/net21_4_ xsel_6_ XI11_3/XI0/XI0_6/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN0_10 XI11_3/net21_5_ xsel_6_ XI11_3/XI0/XI0_6/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN0_9 XI11_3/net21_6_ xsel_6_ XI11_3/XI0/XI0_6/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN0_8 XI11_3/net21_7_ xsel_6_ XI11_3/XI0/XI0_6/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN0_7 XI11_3/net21_8_ xsel_6_ XI11_3/XI0/XI0_6/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN0_6 XI11_3/net21_9_ xsel_6_ XI11_3/XI0/XI0_6/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN0_5 XI11_3/net21_10_ xsel_6_ XI11_3/XI0/XI0_6/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN0_4 XI11_3/net21_11_ xsel_6_ XI11_3/XI0/XI0_6/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN0_3 XI11_3/net21_12_ xsel_6_ XI11_3/XI0/XI0_6/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN0_2 XI11_3/net21_13_ xsel_6_ XI11_3/XI0/XI0_6/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN0_1 XI11_3/net21_14_ xsel_6_ XI11_3/XI0/XI0_6/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN0_0 XI11_3/net21_15_ xsel_6_ XI11_3/XI0/XI0_6/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN1_15 XI11_3/XI0/XI0_6/d__15_ xsel_6_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN1_14 XI11_3/XI0/XI0_6/d__14_ xsel_6_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN1_13 XI11_3/XI0/XI0_6/d__13_ xsel_6_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN1_12 XI11_3/XI0/XI0_6/d__12_ xsel_6_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN1_11 XI11_3/XI0/XI0_6/d__11_ xsel_6_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN1_10 XI11_3/XI0/XI0_6/d__10_ xsel_6_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN1_9 XI11_3/XI0/XI0_6/d__9_ xsel_6_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN1_8 XI11_3/XI0/XI0_6/d__8_ xsel_6_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN1_7 XI11_3/XI0/XI0_6/d__7_ xsel_6_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN1_6 XI11_3/XI0/XI0_6/d__6_ xsel_6_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN1_5 XI11_3/XI0/XI0_6/d__5_ xsel_6_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN1_4 XI11_3/XI0/XI0_6/d__4_ xsel_6_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN1_3 XI11_3/XI0/XI0_6/d__3_ xsel_6_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN1_2 XI11_3/XI0/XI0_6/d__2_ xsel_6_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN1_1 XI11_3/XI0/XI0_6/d__1_ xsel_6_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_6/MN1_0 XI11_3/XI0/XI0_6/d__0_ xsel_6_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN0_15 XI11_3/net21_0_ xsel_5_ XI11_3/XI0/XI0_5/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN0_14 XI11_3/net21_1_ xsel_5_ XI11_3/XI0/XI0_5/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN0_13 XI11_3/net21_2_ xsel_5_ XI11_3/XI0/XI0_5/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN0_12 XI11_3/net21_3_ xsel_5_ XI11_3/XI0/XI0_5/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN0_11 XI11_3/net21_4_ xsel_5_ XI11_3/XI0/XI0_5/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN0_10 XI11_3/net21_5_ xsel_5_ XI11_3/XI0/XI0_5/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN0_9 XI11_3/net21_6_ xsel_5_ XI11_3/XI0/XI0_5/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN0_8 XI11_3/net21_7_ xsel_5_ XI11_3/XI0/XI0_5/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN0_7 XI11_3/net21_8_ xsel_5_ XI11_3/XI0/XI0_5/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN0_6 XI11_3/net21_9_ xsel_5_ XI11_3/XI0/XI0_5/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN0_5 XI11_3/net21_10_ xsel_5_ XI11_3/XI0/XI0_5/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN0_4 XI11_3/net21_11_ xsel_5_ XI11_3/XI0/XI0_5/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN0_3 XI11_3/net21_12_ xsel_5_ XI11_3/XI0/XI0_5/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN0_2 XI11_3/net21_13_ xsel_5_ XI11_3/XI0/XI0_5/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN0_1 XI11_3/net21_14_ xsel_5_ XI11_3/XI0/XI0_5/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN0_0 XI11_3/net21_15_ xsel_5_ XI11_3/XI0/XI0_5/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN1_15 XI11_3/XI0/XI0_5/d__15_ xsel_5_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN1_14 XI11_3/XI0/XI0_5/d__14_ xsel_5_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN1_13 XI11_3/XI0/XI0_5/d__13_ xsel_5_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN1_12 XI11_3/XI0/XI0_5/d__12_ xsel_5_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN1_11 XI11_3/XI0/XI0_5/d__11_ xsel_5_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN1_10 XI11_3/XI0/XI0_5/d__10_ xsel_5_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN1_9 XI11_3/XI0/XI0_5/d__9_ xsel_5_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN1_8 XI11_3/XI0/XI0_5/d__8_ xsel_5_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN1_7 XI11_3/XI0/XI0_5/d__7_ xsel_5_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN1_6 XI11_3/XI0/XI0_5/d__6_ xsel_5_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN1_5 XI11_3/XI0/XI0_5/d__5_ xsel_5_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN1_4 XI11_3/XI0/XI0_5/d__4_ xsel_5_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN1_3 XI11_3/XI0/XI0_5/d__3_ xsel_5_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN1_2 XI11_3/XI0/XI0_5/d__2_ xsel_5_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN1_1 XI11_3/XI0/XI0_5/d__1_ xsel_5_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_5/MN1_0 XI11_3/XI0/XI0_5/d__0_ xsel_5_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN0_15 XI11_3/net21_0_ xsel_4_ XI11_3/XI0/XI0_4/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN0_14 XI11_3/net21_1_ xsel_4_ XI11_3/XI0/XI0_4/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN0_13 XI11_3/net21_2_ xsel_4_ XI11_3/XI0/XI0_4/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN0_12 XI11_3/net21_3_ xsel_4_ XI11_3/XI0/XI0_4/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN0_11 XI11_3/net21_4_ xsel_4_ XI11_3/XI0/XI0_4/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN0_10 XI11_3/net21_5_ xsel_4_ XI11_3/XI0/XI0_4/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN0_9 XI11_3/net21_6_ xsel_4_ XI11_3/XI0/XI0_4/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN0_8 XI11_3/net21_7_ xsel_4_ XI11_3/XI0/XI0_4/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN0_7 XI11_3/net21_8_ xsel_4_ XI11_3/XI0/XI0_4/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN0_6 XI11_3/net21_9_ xsel_4_ XI11_3/XI0/XI0_4/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN0_5 XI11_3/net21_10_ xsel_4_ XI11_3/XI0/XI0_4/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN0_4 XI11_3/net21_11_ xsel_4_ XI11_3/XI0/XI0_4/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN0_3 XI11_3/net21_12_ xsel_4_ XI11_3/XI0/XI0_4/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN0_2 XI11_3/net21_13_ xsel_4_ XI11_3/XI0/XI0_4/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN0_1 XI11_3/net21_14_ xsel_4_ XI11_3/XI0/XI0_4/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN0_0 XI11_3/net21_15_ xsel_4_ XI11_3/XI0/XI0_4/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN1_15 XI11_3/XI0/XI0_4/d__15_ xsel_4_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN1_14 XI11_3/XI0/XI0_4/d__14_ xsel_4_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN1_13 XI11_3/XI0/XI0_4/d__13_ xsel_4_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN1_12 XI11_3/XI0/XI0_4/d__12_ xsel_4_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN1_11 XI11_3/XI0/XI0_4/d__11_ xsel_4_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN1_10 XI11_3/XI0/XI0_4/d__10_ xsel_4_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN1_9 XI11_3/XI0/XI0_4/d__9_ xsel_4_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN1_8 XI11_3/XI0/XI0_4/d__8_ xsel_4_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN1_7 XI11_3/XI0/XI0_4/d__7_ xsel_4_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN1_6 XI11_3/XI0/XI0_4/d__6_ xsel_4_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN1_5 XI11_3/XI0/XI0_4/d__5_ xsel_4_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN1_4 XI11_3/XI0/XI0_4/d__4_ xsel_4_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN1_3 XI11_3/XI0/XI0_4/d__3_ xsel_4_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN1_2 XI11_3/XI0/XI0_4/d__2_ xsel_4_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN1_1 XI11_3/XI0/XI0_4/d__1_ xsel_4_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_4/MN1_0 XI11_3/XI0/XI0_4/d__0_ xsel_4_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN0_15 XI11_3/net21_0_ xsel_3_ XI11_3/XI0/XI0_3/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN0_14 XI11_3/net21_1_ xsel_3_ XI11_3/XI0/XI0_3/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN0_13 XI11_3/net21_2_ xsel_3_ XI11_3/XI0/XI0_3/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN0_12 XI11_3/net21_3_ xsel_3_ XI11_3/XI0/XI0_3/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN0_11 XI11_3/net21_4_ xsel_3_ XI11_3/XI0/XI0_3/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN0_10 XI11_3/net21_5_ xsel_3_ XI11_3/XI0/XI0_3/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN0_9 XI11_3/net21_6_ xsel_3_ XI11_3/XI0/XI0_3/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN0_8 XI11_3/net21_7_ xsel_3_ XI11_3/XI0/XI0_3/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN0_7 XI11_3/net21_8_ xsel_3_ XI11_3/XI0/XI0_3/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN0_6 XI11_3/net21_9_ xsel_3_ XI11_3/XI0/XI0_3/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN0_5 XI11_3/net21_10_ xsel_3_ XI11_3/XI0/XI0_3/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN0_4 XI11_3/net21_11_ xsel_3_ XI11_3/XI0/XI0_3/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN0_3 XI11_3/net21_12_ xsel_3_ XI11_3/XI0/XI0_3/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN0_2 XI11_3/net21_13_ xsel_3_ XI11_3/XI0/XI0_3/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN0_1 XI11_3/net21_14_ xsel_3_ XI11_3/XI0/XI0_3/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN0_0 XI11_3/net21_15_ xsel_3_ XI11_3/XI0/XI0_3/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN1_15 XI11_3/XI0/XI0_3/d__15_ xsel_3_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN1_14 XI11_3/XI0/XI0_3/d__14_ xsel_3_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN1_13 XI11_3/XI0/XI0_3/d__13_ xsel_3_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN1_12 XI11_3/XI0/XI0_3/d__12_ xsel_3_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN1_11 XI11_3/XI0/XI0_3/d__11_ xsel_3_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN1_10 XI11_3/XI0/XI0_3/d__10_ xsel_3_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN1_9 XI11_3/XI0/XI0_3/d__9_ xsel_3_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN1_8 XI11_3/XI0/XI0_3/d__8_ xsel_3_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN1_7 XI11_3/XI0/XI0_3/d__7_ xsel_3_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN1_6 XI11_3/XI0/XI0_3/d__6_ xsel_3_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN1_5 XI11_3/XI0/XI0_3/d__5_ xsel_3_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN1_4 XI11_3/XI0/XI0_3/d__4_ xsel_3_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN1_3 XI11_3/XI0/XI0_3/d__3_ xsel_3_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN1_2 XI11_3/XI0/XI0_3/d__2_ xsel_3_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN1_1 XI11_3/XI0/XI0_3/d__1_ xsel_3_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_3/MN1_0 XI11_3/XI0/XI0_3/d__0_ xsel_3_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN0_15 XI11_3/net21_0_ xsel_2_ XI11_3/XI0/XI0_2/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN0_14 XI11_3/net21_1_ xsel_2_ XI11_3/XI0/XI0_2/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN0_13 XI11_3/net21_2_ xsel_2_ XI11_3/XI0/XI0_2/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN0_12 XI11_3/net21_3_ xsel_2_ XI11_3/XI0/XI0_2/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN0_11 XI11_3/net21_4_ xsel_2_ XI11_3/XI0/XI0_2/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN0_10 XI11_3/net21_5_ xsel_2_ XI11_3/XI0/XI0_2/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN0_9 XI11_3/net21_6_ xsel_2_ XI11_3/XI0/XI0_2/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN0_8 XI11_3/net21_7_ xsel_2_ XI11_3/XI0/XI0_2/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN0_7 XI11_3/net21_8_ xsel_2_ XI11_3/XI0/XI0_2/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN0_6 XI11_3/net21_9_ xsel_2_ XI11_3/XI0/XI0_2/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN0_5 XI11_3/net21_10_ xsel_2_ XI11_3/XI0/XI0_2/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN0_4 XI11_3/net21_11_ xsel_2_ XI11_3/XI0/XI0_2/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN0_3 XI11_3/net21_12_ xsel_2_ XI11_3/XI0/XI0_2/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN0_2 XI11_3/net21_13_ xsel_2_ XI11_3/XI0/XI0_2/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN0_1 XI11_3/net21_14_ xsel_2_ XI11_3/XI0/XI0_2/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN0_0 XI11_3/net21_15_ xsel_2_ XI11_3/XI0/XI0_2/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN1_15 XI11_3/XI0/XI0_2/d__15_ xsel_2_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN1_14 XI11_3/XI0/XI0_2/d__14_ xsel_2_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN1_13 XI11_3/XI0/XI0_2/d__13_ xsel_2_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN1_12 XI11_3/XI0/XI0_2/d__12_ xsel_2_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN1_11 XI11_3/XI0/XI0_2/d__11_ xsel_2_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN1_10 XI11_3/XI0/XI0_2/d__10_ xsel_2_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN1_9 XI11_3/XI0/XI0_2/d__9_ xsel_2_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN1_8 XI11_3/XI0/XI0_2/d__8_ xsel_2_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN1_7 XI11_3/XI0/XI0_2/d__7_ xsel_2_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN1_6 XI11_3/XI0/XI0_2/d__6_ xsel_2_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN1_5 XI11_3/XI0/XI0_2/d__5_ xsel_2_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN1_4 XI11_3/XI0/XI0_2/d__4_ xsel_2_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN1_3 XI11_3/XI0/XI0_2/d__3_ xsel_2_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN1_2 XI11_3/XI0/XI0_2/d__2_ xsel_2_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN1_1 XI11_3/XI0/XI0_2/d__1_ xsel_2_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_2/MN1_0 XI11_3/XI0/XI0_2/d__0_ xsel_2_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN0_15 XI11_3/net21_0_ xsel_1_ XI11_3/XI0/XI0_1/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN0_14 XI11_3/net21_1_ xsel_1_ XI11_3/XI0/XI0_1/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN0_13 XI11_3/net21_2_ xsel_1_ XI11_3/XI0/XI0_1/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN0_12 XI11_3/net21_3_ xsel_1_ XI11_3/XI0/XI0_1/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN0_11 XI11_3/net21_4_ xsel_1_ XI11_3/XI0/XI0_1/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN0_10 XI11_3/net21_5_ xsel_1_ XI11_3/XI0/XI0_1/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN0_9 XI11_3/net21_6_ xsel_1_ XI11_3/XI0/XI0_1/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN0_8 XI11_3/net21_7_ xsel_1_ XI11_3/XI0/XI0_1/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN0_7 XI11_3/net21_8_ xsel_1_ XI11_3/XI0/XI0_1/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN0_6 XI11_3/net21_9_ xsel_1_ XI11_3/XI0/XI0_1/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN0_5 XI11_3/net21_10_ xsel_1_ XI11_3/XI0/XI0_1/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN0_4 XI11_3/net21_11_ xsel_1_ XI11_3/XI0/XI0_1/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN0_3 XI11_3/net21_12_ xsel_1_ XI11_3/XI0/XI0_1/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN0_2 XI11_3/net21_13_ xsel_1_ XI11_3/XI0/XI0_1/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN0_1 XI11_3/net21_14_ xsel_1_ XI11_3/XI0/XI0_1/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN0_0 XI11_3/net21_15_ xsel_1_ XI11_3/XI0/XI0_1/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN1_15 XI11_3/XI0/XI0_1/d__15_ xsel_1_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN1_14 XI11_3/XI0/XI0_1/d__14_ xsel_1_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN1_13 XI11_3/XI0/XI0_1/d__13_ xsel_1_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN1_12 XI11_3/XI0/XI0_1/d__12_ xsel_1_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN1_11 XI11_3/XI0/XI0_1/d__11_ xsel_1_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN1_10 XI11_3/XI0/XI0_1/d__10_ xsel_1_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN1_9 XI11_3/XI0/XI0_1/d__9_ xsel_1_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN1_8 XI11_3/XI0/XI0_1/d__8_ xsel_1_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN1_7 XI11_3/XI0/XI0_1/d__7_ xsel_1_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN1_6 XI11_3/XI0/XI0_1/d__6_ xsel_1_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN1_5 XI11_3/XI0/XI0_1/d__5_ xsel_1_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN1_4 XI11_3/XI0/XI0_1/d__4_ xsel_1_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN1_3 XI11_3/XI0/XI0_1/d__3_ xsel_1_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN1_2 XI11_3/XI0/XI0_1/d__2_ xsel_1_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN1_1 XI11_3/XI0/XI0_1/d__1_ xsel_1_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_1/MN1_0 XI11_3/XI0/XI0_1/d__0_ xsel_1_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN0_15 XI11_3/net21_0_ xsel_0_ XI11_3/XI0/XI0_0/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN0_14 XI11_3/net21_1_ xsel_0_ XI11_3/XI0/XI0_0/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN0_13 XI11_3/net21_2_ xsel_0_ XI11_3/XI0/XI0_0/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN0_12 XI11_3/net21_3_ xsel_0_ XI11_3/XI0/XI0_0/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN0_11 XI11_3/net21_4_ xsel_0_ XI11_3/XI0/XI0_0/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN0_10 XI11_3/net21_5_ xsel_0_ XI11_3/XI0/XI0_0/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN0_9 XI11_3/net21_6_ xsel_0_ XI11_3/XI0/XI0_0/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN0_8 XI11_3/net21_7_ xsel_0_ XI11_3/XI0/XI0_0/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN0_7 XI11_3/net21_8_ xsel_0_ XI11_3/XI0/XI0_0/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN0_6 XI11_3/net21_9_ xsel_0_ XI11_3/XI0/XI0_0/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN0_5 XI11_3/net21_10_ xsel_0_ XI11_3/XI0/XI0_0/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN0_4 XI11_3/net21_11_ xsel_0_ XI11_3/XI0/XI0_0/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN0_3 XI11_3/net21_12_ xsel_0_ XI11_3/XI0/XI0_0/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN0_2 XI11_3/net21_13_ xsel_0_ XI11_3/XI0/XI0_0/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN0_1 XI11_3/net21_14_ xsel_0_ XI11_3/XI0/XI0_0/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN0_0 XI11_3/net21_15_ xsel_0_ XI11_3/XI0/XI0_0/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN1_15 XI11_3/XI0/XI0_0/d__15_ xsel_0_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN1_14 XI11_3/XI0/XI0_0/d__14_ xsel_0_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN1_13 XI11_3/XI0/XI0_0/d__13_ xsel_0_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN1_12 XI11_3/XI0/XI0_0/d__12_ xsel_0_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN1_11 XI11_3/XI0/XI0_0/d__11_ xsel_0_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN1_10 XI11_3/XI0/XI0_0/d__10_ xsel_0_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN1_9 XI11_3/XI0/XI0_0/d__9_ xsel_0_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN1_8 XI11_3/XI0/XI0_0/d__8_ xsel_0_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN1_7 XI11_3/XI0/XI0_0/d__7_ xsel_0_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN1_6 XI11_3/XI0/XI0_0/d__6_ xsel_0_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN1_5 XI11_3/XI0/XI0_0/d__5_ xsel_0_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN1_4 XI11_3/XI0/XI0_0/d__4_ xsel_0_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN1_3 XI11_3/XI0/XI0_0/d__3_ xsel_0_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN1_2 XI11_3/XI0/XI0_0/d__2_ xsel_0_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN1_1 XI11_3/XI0/XI0_0/d__1_ xsel_0_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_0/MN1_0 XI11_3/XI0/XI0_0/d__0_ xsel_0_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI2/MN0_15 XI11_2/net21_0_ ysel_15_ XI11_2/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN0_14 XI11_2/net21_1_ ysel_14_ XI11_2/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN0_13 XI11_2/net21_2_ ysel_13_ XI11_2/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN0_12 XI11_2/net21_3_ ysel_12_ XI11_2/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN0_11 XI11_2/net21_4_ ysel_11_ XI11_2/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN0_10 XI11_2/net21_5_ ysel_10_ XI11_2/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN0_9 XI11_2/net21_6_ ysel_9_ XI11_2/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN0_8 XI11_2/net21_7_ ysel_8_ XI11_2/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN0_7 XI11_2/net21_8_ ysel_7_ XI11_2/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN0_6 XI11_2/net21_9_ ysel_6_ XI11_2/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN0_5 XI11_2/net21_10_ ysel_5_ XI11_2/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN0_4 XI11_2/net21_11_ ysel_4_ XI11_2/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN0_3 XI11_2/net21_12_ ysel_3_ XI11_2/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN0_2 XI11_2/net21_13_ ysel_2_ XI11_2/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN0_1 XI11_2/net21_14_ ysel_1_ XI11_2/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN0_0 XI11_2/net21_15_ ysel_0_ XI11_2/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN1_15 XI11_2/net20_0_ ysel_15_ XI11_2/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN1_14 XI11_2/net20_1_ ysel_14_ XI11_2/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN1_13 XI11_2/net20_2_ ysel_13_ XI11_2/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN1_12 XI11_2/net20_3_ ysel_12_ XI11_2/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN1_11 XI11_2/net20_4_ ysel_11_ XI11_2/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN1_10 XI11_2/net20_5_ ysel_10_ XI11_2/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN1_9 XI11_2/net20_6_ ysel_9_ XI11_2/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN1_8 XI11_2/net20_7_ ysel_8_ XI11_2/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN1_7 XI11_2/net20_8_ ysel_7_ XI11_2/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN1_6 XI11_2/net20_9_ ysel_6_ XI11_2/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN1_5 XI11_2/net20_10_ ysel_5_ XI11_2/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN1_4 XI11_2/net20_11_ ysel_4_ XI11_2/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN1_3 XI11_2/net20_12_ ysel_3_ XI11_2/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN1_2 XI11_2/net20_13_ ysel_2_ XI11_2/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN1_1 XI11_2/net20_14_ ysel_1_ XI11_2/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI2/MN1_0 XI11_2/net20_15_ ysel_0_ XI11_2/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_2/XI4/MN8 vdd XI11_2/XI4/net8 XI11_2/net12 vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_2/XI4/MP0 XI11_2/net9 XI11_2/XI4/net23 vdd vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_2/XI4/MP4 XI11_2/net12 XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI4/MP1 XI11_2/net9 XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI4/MP5 XI11_2/net12 XI11_2/preck XI11_2/net9 vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI4/MN7 vdd XI11_2/XI4/net090 DOUT_2_ vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_2/XI4/MP3 gnd XI11_2/XI4/net089 XI11_2/net12 gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_2/XI4/MN5 XI11_2/net9 XI11_2/XI4/net0103 gnd gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_2/XI4/MN4 XI11_2/XI4/data_out_ XI11_2/XI4/net32 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_2/XI4/MN0 XI11_2/XI4/data_out XI11_2/XI4/net52 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_2/XI4/MN9 gnd XI11_2/XI4/net0112 DOUT_2_ gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_2/XI1_15/MP2 XI11_2/net20_0_ XI11_2/preck XI11_2/net21_0_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI1_15/MP1 XI11_2/net20_0_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_15/MP0 XI11_2/net21_0_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_14/MP2 XI11_2/net20_1_ XI11_2/preck XI11_2/net21_1_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI1_14/MP1 XI11_2/net20_1_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_14/MP0 XI11_2/net21_1_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_13/MP2 XI11_2/net20_2_ XI11_2/preck XI11_2/net21_2_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI1_13/MP1 XI11_2/net20_2_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_13/MP0 XI11_2/net21_2_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_12/MP2 XI11_2/net20_3_ XI11_2/preck XI11_2/net21_3_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI1_12/MP1 XI11_2/net20_3_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_12/MP0 XI11_2/net21_3_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_11/MP2 XI11_2/net20_4_ XI11_2/preck XI11_2/net21_4_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI1_11/MP1 XI11_2/net20_4_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_11/MP0 XI11_2/net21_4_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_10/MP2 XI11_2/net20_5_ XI11_2/preck XI11_2/net21_5_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI1_10/MP1 XI11_2/net20_5_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_10/MP0 XI11_2/net21_5_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_9/MP2 XI11_2/net20_6_ XI11_2/preck XI11_2/net21_6_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI1_9/MP1 XI11_2/net20_6_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_9/MP0 XI11_2/net21_6_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_8/MP2 XI11_2/net20_7_ XI11_2/preck XI11_2/net21_7_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI1_8/MP1 XI11_2/net20_7_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_8/MP0 XI11_2/net21_7_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_7/MP2 XI11_2/net20_8_ XI11_2/preck XI11_2/net21_8_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI1_7/MP1 XI11_2/net20_8_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_7/MP0 XI11_2/net21_8_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_6/MP2 XI11_2/net20_9_ XI11_2/preck XI11_2/net21_9_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI1_6/MP1 XI11_2/net20_9_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_6/MP0 XI11_2/net21_9_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_5/MP2 XI11_2/net20_10_ XI11_2/preck XI11_2/net21_10_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI1_5/MP1 XI11_2/net20_10_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_5/MP0 XI11_2/net21_10_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_4/MP2 XI11_2/net20_11_ XI11_2/preck XI11_2/net21_11_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI1_4/MP1 XI11_2/net20_11_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_4/MP0 XI11_2/net21_11_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_3/MP2 XI11_2/net20_12_ XI11_2/preck XI11_2/net21_12_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI1_3/MP1 XI11_2/net20_12_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_3/MP0 XI11_2/net21_12_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_2/MP2 XI11_2/net20_13_ XI11_2/preck XI11_2/net21_13_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI1_2/MP1 XI11_2/net20_13_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_2/MP0 XI11_2/net21_13_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_1/MP2 XI11_2/net20_14_ XI11_2/preck XI11_2/net21_14_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI1_1/MP1 XI11_2/net20_14_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_1/MP0 XI11_2/net21_14_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_0/MP2 XI11_2/net20_15_ XI11_2/preck XI11_2/net21_15_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_2/XI1_0/MP1 XI11_2/net20_15_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI1_0/MP0 XI11_2/net21_15_ XI11_2/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_2/XI0/MN0_15 gnd gnd XI11_2/net21_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN0_14 gnd gnd XI11_2/net21_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN0_13 gnd gnd XI11_2/net21_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN0_12 gnd gnd XI11_2/net21_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN0_11 gnd gnd XI11_2/net21_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN0_10 gnd gnd XI11_2/net21_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN0_9 gnd gnd XI11_2/net21_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN0_8 gnd gnd XI11_2/net21_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN0_7 gnd gnd XI11_2/net21_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN0_6 gnd gnd XI11_2/net21_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN0_5 gnd gnd XI11_2/net21_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN0_4 gnd gnd XI11_2/net21_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN0_3 gnd gnd XI11_2/net21_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN0_2 gnd gnd XI11_2/net21_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN0_1 gnd gnd XI11_2/net21_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN0_0 gnd gnd XI11_2/net21_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN1_15 gnd gnd XI11_2/net20_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN1_14 gnd gnd XI11_2/net20_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN1_13 gnd gnd XI11_2/net20_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN1_12 gnd gnd XI11_2/net20_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN1_11 gnd gnd XI11_2/net20_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN1_10 gnd gnd XI11_2/net20_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN1_9 gnd gnd XI11_2/net20_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN1_8 gnd gnd XI11_2/net20_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN1_7 gnd gnd XI11_2/net20_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN1_6 gnd gnd XI11_2/net20_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN1_5 gnd gnd XI11_2/net20_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN1_4 gnd gnd XI11_2/net20_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN1_3 gnd gnd XI11_2/net20_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN1_2 gnd gnd XI11_2/net20_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN1_1 gnd gnd XI11_2/net20_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/MN1_0 gnd gnd XI11_2/net20_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN0_15 XI11_2/net21_0_ xsel_63_ XI11_2/XI0/XI0_63/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN0_14 XI11_2/net21_1_ xsel_63_ XI11_2/XI0/XI0_63/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN0_13 XI11_2/net21_2_ xsel_63_ XI11_2/XI0/XI0_63/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN0_12 XI11_2/net21_3_ xsel_63_ XI11_2/XI0/XI0_63/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN0_11 XI11_2/net21_4_ xsel_63_ XI11_2/XI0/XI0_63/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN0_10 XI11_2/net21_5_ xsel_63_ XI11_2/XI0/XI0_63/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN0_9 XI11_2/net21_6_ xsel_63_ XI11_2/XI0/XI0_63/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN0_8 XI11_2/net21_7_ xsel_63_ XI11_2/XI0/XI0_63/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN0_7 XI11_2/net21_8_ xsel_63_ XI11_2/XI0/XI0_63/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN0_6 XI11_2/net21_9_ xsel_63_ XI11_2/XI0/XI0_63/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN0_5 XI11_2/net21_10_ xsel_63_ XI11_2/XI0/XI0_63/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN0_4 XI11_2/net21_11_ xsel_63_ XI11_2/XI0/XI0_63/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN0_3 XI11_2/net21_12_ xsel_63_ XI11_2/XI0/XI0_63/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN0_2 XI11_2/net21_13_ xsel_63_ XI11_2/XI0/XI0_63/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN0_1 XI11_2/net21_14_ xsel_63_ XI11_2/XI0/XI0_63/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN0_0 XI11_2/net21_15_ xsel_63_ XI11_2/XI0/XI0_63/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN1_15 XI11_2/XI0/XI0_63/d__15_ xsel_63_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN1_14 XI11_2/XI0/XI0_63/d__14_ xsel_63_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN1_13 XI11_2/XI0/XI0_63/d__13_ xsel_63_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN1_12 XI11_2/XI0/XI0_63/d__12_ xsel_63_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN1_11 XI11_2/XI0/XI0_63/d__11_ xsel_63_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN1_10 XI11_2/XI0/XI0_63/d__10_ xsel_63_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN1_9 XI11_2/XI0/XI0_63/d__9_ xsel_63_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN1_8 XI11_2/XI0/XI0_63/d__8_ xsel_63_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN1_7 XI11_2/XI0/XI0_63/d__7_ xsel_63_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN1_6 XI11_2/XI0/XI0_63/d__6_ xsel_63_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN1_5 XI11_2/XI0/XI0_63/d__5_ xsel_63_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN1_4 XI11_2/XI0/XI0_63/d__4_ xsel_63_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN1_3 XI11_2/XI0/XI0_63/d__3_ xsel_63_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN1_2 XI11_2/XI0/XI0_63/d__2_ xsel_63_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN1_1 XI11_2/XI0/XI0_63/d__1_ xsel_63_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_63/MN1_0 XI11_2/XI0/XI0_63/d__0_ xsel_63_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN0_15 XI11_2/net21_0_ xsel_62_ XI11_2/XI0/XI0_62/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN0_14 XI11_2/net21_1_ xsel_62_ XI11_2/XI0/XI0_62/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN0_13 XI11_2/net21_2_ xsel_62_ XI11_2/XI0/XI0_62/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN0_12 XI11_2/net21_3_ xsel_62_ XI11_2/XI0/XI0_62/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN0_11 XI11_2/net21_4_ xsel_62_ XI11_2/XI0/XI0_62/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN0_10 XI11_2/net21_5_ xsel_62_ XI11_2/XI0/XI0_62/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN0_9 XI11_2/net21_6_ xsel_62_ XI11_2/XI0/XI0_62/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN0_8 XI11_2/net21_7_ xsel_62_ XI11_2/XI0/XI0_62/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN0_7 XI11_2/net21_8_ xsel_62_ XI11_2/XI0/XI0_62/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN0_6 XI11_2/net21_9_ xsel_62_ XI11_2/XI0/XI0_62/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN0_5 XI11_2/net21_10_ xsel_62_ XI11_2/XI0/XI0_62/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN0_4 XI11_2/net21_11_ xsel_62_ XI11_2/XI0/XI0_62/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN0_3 XI11_2/net21_12_ xsel_62_ XI11_2/XI0/XI0_62/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN0_2 XI11_2/net21_13_ xsel_62_ XI11_2/XI0/XI0_62/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN0_1 XI11_2/net21_14_ xsel_62_ XI11_2/XI0/XI0_62/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN0_0 XI11_2/net21_15_ xsel_62_ XI11_2/XI0/XI0_62/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN1_15 XI11_2/XI0/XI0_62/d__15_ xsel_62_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN1_14 XI11_2/XI0/XI0_62/d__14_ xsel_62_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN1_13 XI11_2/XI0/XI0_62/d__13_ xsel_62_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN1_12 XI11_2/XI0/XI0_62/d__12_ xsel_62_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN1_11 XI11_2/XI0/XI0_62/d__11_ xsel_62_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN1_10 XI11_2/XI0/XI0_62/d__10_ xsel_62_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN1_9 XI11_2/XI0/XI0_62/d__9_ xsel_62_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN1_8 XI11_2/XI0/XI0_62/d__8_ xsel_62_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN1_7 XI11_2/XI0/XI0_62/d__7_ xsel_62_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN1_6 XI11_2/XI0/XI0_62/d__6_ xsel_62_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN1_5 XI11_2/XI0/XI0_62/d__5_ xsel_62_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN1_4 XI11_2/XI0/XI0_62/d__4_ xsel_62_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN1_3 XI11_2/XI0/XI0_62/d__3_ xsel_62_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN1_2 XI11_2/XI0/XI0_62/d__2_ xsel_62_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN1_1 XI11_2/XI0/XI0_62/d__1_ xsel_62_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_62/MN1_0 XI11_2/XI0/XI0_62/d__0_ xsel_62_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN0_15 XI11_2/net21_0_ xsel_61_ XI11_2/XI0/XI0_61/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN0_14 XI11_2/net21_1_ xsel_61_ XI11_2/XI0/XI0_61/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN0_13 XI11_2/net21_2_ xsel_61_ XI11_2/XI0/XI0_61/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN0_12 XI11_2/net21_3_ xsel_61_ XI11_2/XI0/XI0_61/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN0_11 XI11_2/net21_4_ xsel_61_ XI11_2/XI0/XI0_61/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN0_10 XI11_2/net21_5_ xsel_61_ XI11_2/XI0/XI0_61/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN0_9 XI11_2/net21_6_ xsel_61_ XI11_2/XI0/XI0_61/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN0_8 XI11_2/net21_7_ xsel_61_ XI11_2/XI0/XI0_61/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN0_7 XI11_2/net21_8_ xsel_61_ XI11_2/XI0/XI0_61/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN0_6 XI11_2/net21_9_ xsel_61_ XI11_2/XI0/XI0_61/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN0_5 XI11_2/net21_10_ xsel_61_ XI11_2/XI0/XI0_61/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN0_4 XI11_2/net21_11_ xsel_61_ XI11_2/XI0/XI0_61/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN0_3 XI11_2/net21_12_ xsel_61_ XI11_2/XI0/XI0_61/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN0_2 XI11_2/net21_13_ xsel_61_ XI11_2/XI0/XI0_61/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN0_1 XI11_2/net21_14_ xsel_61_ XI11_2/XI0/XI0_61/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN0_0 XI11_2/net21_15_ xsel_61_ XI11_2/XI0/XI0_61/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN1_15 XI11_2/XI0/XI0_61/d__15_ xsel_61_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN1_14 XI11_2/XI0/XI0_61/d__14_ xsel_61_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN1_13 XI11_2/XI0/XI0_61/d__13_ xsel_61_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN1_12 XI11_2/XI0/XI0_61/d__12_ xsel_61_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN1_11 XI11_2/XI0/XI0_61/d__11_ xsel_61_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN1_10 XI11_2/XI0/XI0_61/d__10_ xsel_61_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN1_9 XI11_2/XI0/XI0_61/d__9_ xsel_61_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN1_8 XI11_2/XI0/XI0_61/d__8_ xsel_61_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN1_7 XI11_2/XI0/XI0_61/d__7_ xsel_61_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN1_6 XI11_2/XI0/XI0_61/d__6_ xsel_61_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN1_5 XI11_2/XI0/XI0_61/d__5_ xsel_61_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN1_4 XI11_2/XI0/XI0_61/d__4_ xsel_61_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN1_3 XI11_2/XI0/XI0_61/d__3_ xsel_61_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN1_2 XI11_2/XI0/XI0_61/d__2_ xsel_61_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN1_1 XI11_2/XI0/XI0_61/d__1_ xsel_61_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_61/MN1_0 XI11_2/XI0/XI0_61/d__0_ xsel_61_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN0_15 XI11_2/net21_0_ xsel_60_ XI11_2/XI0/XI0_60/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN0_14 XI11_2/net21_1_ xsel_60_ XI11_2/XI0/XI0_60/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN0_13 XI11_2/net21_2_ xsel_60_ XI11_2/XI0/XI0_60/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN0_12 XI11_2/net21_3_ xsel_60_ XI11_2/XI0/XI0_60/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN0_11 XI11_2/net21_4_ xsel_60_ XI11_2/XI0/XI0_60/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN0_10 XI11_2/net21_5_ xsel_60_ XI11_2/XI0/XI0_60/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN0_9 XI11_2/net21_6_ xsel_60_ XI11_2/XI0/XI0_60/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN0_8 XI11_2/net21_7_ xsel_60_ XI11_2/XI0/XI0_60/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN0_7 XI11_2/net21_8_ xsel_60_ XI11_2/XI0/XI0_60/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN0_6 XI11_2/net21_9_ xsel_60_ XI11_2/XI0/XI0_60/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN0_5 XI11_2/net21_10_ xsel_60_ XI11_2/XI0/XI0_60/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN0_4 XI11_2/net21_11_ xsel_60_ XI11_2/XI0/XI0_60/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN0_3 XI11_2/net21_12_ xsel_60_ XI11_2/XI0/XI0_60/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN0_2 XI11_2/net21_13_ xsel_60_ XI11_2/XI0/XI0_60/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN0_1 XI11_2/net21_14_ xsel_60_ XI11_2/XI0/XI0_60/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN0_0 XI11_2/net21_15_ xsel_60_ XI11_2/XI0/XI0_60/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN1_15 XI11_2/XI0/XI0_60/d__15_ xsel_60_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN1_14 XI11_2/XI0/XI0_60/d__14_ xsel_60_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN1_13 XI11_2/XI0/XI0_60/d__13_ xsel_60_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN1_12 XI11_2/XI0/XI0_60/d__12_ xsel_60_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN1_11 XI11_2/XI0/XI0_60/d__11_ xsel_60_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN1_10 XI11_2/XI0/XI0_60/d__10_ xsel_60_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN1_9 XI11_2/XI0/XI0_60/d__9_ xsel_60_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN1_8 XI11_2/XI0/XI0_60/d__8_ xsel_60_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN1_7 XI11_2/XI0/XI0_60/d__7_ xsel_60_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN1_6 XI11_2/XI0/XI0_60/d__6_ xsel_60_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN1_5 XI11_2/XI0/XI0_60/d__5_ xsel_60_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN1_4 XI11_2/XI0/XI0_60/d__4_ xsel_60_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN1_3 XI11_2/XI0/XI0_60/d__3_ xsel_60_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN1_2 XI11_2/XI0/XI0_60/d__2_ xsel_60_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN1_1 XI11_2/XI0/XI0_60/d__1_ xsel_60_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_60/MN1_0 XI11_2/XI0/XI0_60/d__0_ xsel_60_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN0_15 XI11_2/net21_0_ xsel_59_ XI11_2/XI0/XI0_59/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN0_14 XI11_2/net21_1_ xsel_59_ XI11_2/XI0/XI0_59/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN0_13 XI11_2/net21_2_ xsel_59_ XI11_2/XI0/XI0_59/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN0_12 XI11_2/net21_3_ xsel_59_ XI11_2/XI0/XI0_59/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN0_11 XI11_2/net21_4_ xsel_59_ XI11_2/XI0/XI0_59/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN0_10 XI11_2/net21_5_ xsel_59_ XI11_2/XI0/XI0_59/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN0_9 XI11_2/net21_6_ xsel_59_ XI11_2/XI0/XI0_59/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN0_8 XI11_2/net21_7_ xsel_59_ XI11_2/XI0/XI0_59/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN0_7 XI11_2/net21_8_ xsel_59_ XI11_2/XI0/XI0_59/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN0_6 XI11_2/net21_9_ xsel_59_ XI11_2/XI0/XI0_59/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN0_5 XI11_2/net21_10_ xsel_59_ XI11_2/XI0/XI0_59/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN0_4 XI11_2/net21_11_ xsel_59_ XI11_2/XI0/XI0_59/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN0_3 XI11_2/net21_12_ xsel_59_ XI11_2/XI0/XI0_59/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN0_2 XI11_2/net21_13_ xsel_59_ XI11_2/XI0/XI0_59/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN0_1 XI11_2/net21_14_ xsel_59_ XI11_2/XI0/XI0_59/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN0_0 XI11_2/net21_15_ xsel_59_ XI11_2/XI0/XI0_59/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN1_15 XI11_2/XI0/XI0_59/d__15_ xsel_59_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN1_14 XI11_2/XI0/XI0_59/d__14_ xsel_59_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN1_13 XI11_2/XI0/XI0_59/d__13_ xsel_59_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN1_12 XI11_2/XI0/XI0_59/d__12_ xsel_59_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN1_11 XI11_2/XI0/XI0_59/d__11_ xsel_59_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN1_10 XI11_2/XI0/XI0_59/d__10_ xsel_59_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN1_9 XI11_2/XI0/XI0_59/d__9_ xsel_59_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN1_8 XI11_2/XI0/XI0_59/d__8_ xsel_59_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN1_7 XI11_2/XI0/XI0_59/d__7_ xsel_59_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN1_6 XI11_2/XI0/XI0_59/d__6_ xsel_59_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN1_5 XI11_2/XI0/XI0_59/d__5_ xsel_59_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN1_4 XI11_2/XI0/XI0_59/d__4_ xsel_59_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN1_3 XI11_2/XI0/XI0_59/d__3_ xsel_59_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN1_2 XI11_2/XI0/XI0_59/d__2_ xsel_59_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN1_1 XI11_2/XI0/XI0_59/d__1_ xsel_59_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_59/MN1_0 XI11_2/XI0/XI0_59/d__0_ xsel_59_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN0_15 XI11_2/net21_0_ xsel_58_ XI11_2/XI0/XI0_58/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN0_14 XI11_2/net21_1_ xsel_58_ XI11_2/XI0/XI0_58/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN0_13 XI11_2/net21_2_ xsel_58_ XI11_2/XI0/XI0_58/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN0_12 XI11_2/net21_3_ xsel_58_ XI11_2/XI0/XI0_58/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN0_11 XI11_2/net21_4_ xsel_58_ XI11_2/XI0/XI0_58/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN0_10 XI11_2/net21_5_ xsel_58_ XI11_2/XI0/XI0_58/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN0_9 XI11_2/net21_6_ xsel_58_ XI11_2/XI0/XI0_58/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN0_8 XI11_2/net21_7_ xsel_58_ XI11_2/XI0/XI0_58/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN0_7 XI11_2/net21_8_ xsel_58_ XI11_2/XI0/XI0_58/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN0_6 XI11_2/net21_9_ xsel_58_ XI11_2/XI0/XI0_58/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN0_5 XI11_2/net21_10_ xsel_58_ XI11_2/XI0/XI0_58/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN0_4 XI11_2/net21_11_ xsel_58_ XI11_2/XI0/XI0_58/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN0_3 XI11_2/net21_12_ xsel_58_ XI11_2/XI0/XI0_58/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN0_2 XI11_2/net21_13_ xsel_58_ XI11_2/XI0/XI0_58/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN0_1 XI11_2/net21_14_ xsel_58_ XI11_2/XI0/XI0_58/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN0_0 XI11_2/net21_15_ xsel_58_ XI11_2/XI0/XI0_58/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN1_15 XI11_2/XI0/XI0_58/d__15_ xsel_58_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN1_14 XI11_2/XI0/XI0_58/d__14_ xsel_58_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN1_13 XI11_2/XI0/XI0_58/d__13_ xsel_58_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN1_12 XI11_2/XI0/XI0_58/d__12_ xsel_58_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN1_11 XI11_2/XI0/XI0_58/d__11_ xsel_58_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN1_10 XI11_2/XI0/XI0_58/d__10_ xsel_58_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN1_9 XI11_2/XI0/XI0_58/d__9_ xsel_58_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN1_8 XI11_2/XI0/XI0_58/d__8_ xsel_58_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN1_7 XI11_2/XI0/XI0_58/d__7_ xsel_58_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN1_6 XI11_2/XI0/XI0_58/d__6_ xsel_58_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN1_5 XI11_2/XI0/XI0_58/d__5_ xsel_58_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN1_4 XI11_2/XI0/XI0_58/d__4_ xsel_58_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN1_3 XI11_2/XI0/XI0_58/d__3_ xsel_58_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN1_2 XI11_2/XI0/XI0_58/d__2_ xsel_58_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN1_1 XI11_2/XI0/XI0_58/d__1_ xsel_58_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_58/MN1_0 XI11_2/XI0/XI0_58/d__0_ xsel_58_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN0_15 XI11_2/net21_0_ xsel_57_ XI11_2/XI0/XI0_57/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN0_14 XI11_2/net21_1_ xsel_57_ XI11_2/XI0/XI0_57/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN0_13 XI11_2/net21_2_ xsel_57_ XI11_2/XI0/XI0_57/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN0_12 XI11_2/net21_3_ xsel_57_ XI11_2/XI0/XI0_57/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN0_11 XI11_2/net21_4_ xsel_57_ XI11_2/XI0/XI0_57/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN0_10 XI11_2/net21_5_ xsel_57_ XI11_2/XI0/XI0_57/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN0_9 XI11_2/net21_6_ xsel_57_ XI11_2/XI0/XI0_57/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN0_8 XI11_2/net21_7_ xsel_57_ XI11_2/XI0/XI0_57/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN0_7 XI11_2/net21_8_ xsel_57_ XI11_2/XI0/XI0_57/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN0_6 XI11_2/net21_9_ xsel_57_ XI11_2/XI0/XI0_57/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN0_5 XI11_2/net21_10_ xsel_57_ XI11_2/XI0/XI0_57/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN0_4 XI11_2/net21_11_ xsel_57_ XI11_2/XI0/XI0_57/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN0_3 XI11_2/net21_12_ xsel_57_ XI11_2/XI0/XI0_57/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN0_2 XI11_2/net21_13_ xsel_57_ XI11_2/XI0/XI0_57/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN0_1 XI11_2/net21_14_ xsel_57_ XI11_2/XI0/XI0_57/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN0_0 XI11_2/net21_15_ xsel_57_ XI11_2/XI0/XI0_57/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN1_15 XI11_2/XI0/XI0_57/d__15_ xsel_57_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN1_14 XI11_2/XI0/XI0_57/d__14_ xsel_57_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN1_13 XI11_2/XI0/XI0_57/d__13_ xsel_57_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN1_12 XI11_2/XI0/XI0_57/d__12_ xsel_57_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN1_11 XI11_2/XI0/XI0_57/d__11_ xsel_57_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN1_10 XI11_2/XI0/XI0_57/d__10_ xsel_57_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN1_9 XI11_2/XI0/XI0_57/d__9_ xsel_57_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN1_8 XI11_2/XI0/XI0_57/d__8_ xsel_57_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN1_7 XI11_2/XI0/XI0_57/d__7_ xsel_57_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN1_6 XI11_2/XI0/XI0_57/d__6_ xsel_57_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN1_5 XI11_2/XI0/XI0_57/d__5_ xsel_57_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN1_4 XI11_2/XI0/XI0_57/d__4_ xsel_57_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN1_3 XI11_2/XI0/XI0_57/d__3_ xsel_57_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN1_2 XI11_2/XI0/XI0_57/d__2_ xsel_57_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN1_1 XI11_2/XI0/XI0_57/d__1_ xsel_57_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_57/MN1_0 XI11_2/XI0/XI0_57/d__0_ xsel_57_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN0_15 XI11_2/net21_0_ xsel_56_ XI11_2/XI0/XI0_56/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN0_14 XI11_2/net21_1_ xsel_56_ XI11_2/XI0/XI0_56/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN0_13 XI11_2/net21_2_ xsel_56_ XI11_2/XI0/XI0_56/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN0_12 XI11_2/net21_3_ xsel_56_ XI11_2/XI0/XI0_56/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN0_11 XI11_2/net21_4_ xsel_56_ XI11_2/XI0/XI0_56/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN0_10 XI11_2/net21_5_ xsel_56_ XI11_2/XI0/XI0_56/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN0_9 XI11_2/net21_6_ xsel_56_ XI11_2/XI0/XI0_56/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN0_8 XI11_2/net21_7_ xsel_56_ XI11_2/XI0/XI0_56/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN0_7 XI11_2/net21_8_ xsel_56_ XI11_2/XI0/XI0_56/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN0_6 XI11_2/net21_9_ xsel_56_ XI11_2/XI0/XI0_56/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN0_5 XI11_2/net21_10_ xsel_56_ XI11_2/XI0/XI0_56/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN0_4 XI11_2/net21_11_ xsel_56_ XI11_2/XI0/XI0_56/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN0_3 XI11_2/net21_12_ xsel_56_ XI11_2/XI0/XI0_56/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN0_2 XI11_2/net21_13_ xsel_56_ XI11_2/XI0/XI0_56/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN0_1 XI11_2/net21_14_ xsel_56_ XI11_2/XI0/XI0_56/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN0_0 XI11_2/net21_15_ xsel_56_ XI11_2/XI0/XI0_56/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN1_15 XI11_2/XI0/XI0_56/d__15_ xsel_56_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN1_14 XI11_2/XI0/XI0_56/d__14_ xsel_56_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN1_13 XI11_2/XI0/XI0_56/d__13_ xsel_56_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN1_12 XI11_2/XI0/XI0_56/d__12_ xsel_56_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN1_11 XI11_2/XI0/XI0_56/d__11_ xsel_56_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN1_10 XI11_2/XI0/XI0_56/d__10_ xsel_56_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN1_9 XI11_2/XI0/XI0_56/d__9_ xsel_56_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN1_8 XI11_2/XI0/XI0_56/d__8_ xsel_56_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN1_7 XI11_2/XI0/XI0_56/d__7_ xsel_56_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN1_6 XI11_2/XI0/XI0_56/d__6_ xsel_56_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN1_5 XI11_2/XI0/XI0_56/d__5_ xsel_56_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN1_4 XI11_2/XI0/XI0_56/d__4_ xsel_56_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN1_3 XI11_2/XI0/XI0_56/d__3_ xsel_56_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN1_2 XI11_2/XI0/XI0_56/d__2_ xsel_56_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN1_1 XI11_2/XI0/XI0_56/d__1_ xsel_56_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_56/MN1_0 XI11_2/XI0/XI0_56/d__0_ xsel_56_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN0_15 XI11_2/net21_0_ xsel_55_ XI11_2/XI0/XI0_55/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN0_14 XI11_2/net21_1_ xsel_55_ XI11_2/XI0/XI0_55/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN0_13 XI11_2/net21_2_ xsel_55_ XI11_2/XI0/XI0_55/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN0_12 XI11_2/net21_3_ xsel_55_ XI11_2/XI0/XI0_55/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN0_11 XI11_2/net21_4_ xsel_55_ XI11_2/XI0/XI0_55/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN0_10 XI11_2/net21_5_ xsel_55_ XI11_2/XI0/XI0_55/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN0_9 XI11_2/net21_6_ xsel_55_ XI11_2/XI0/XI0_55/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN0_8 XI11_2/net21_7_ xsel_55_ XI11_2/XI0/XI0_55/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN0_7 XI11_2/net21_8_ xsel_55_ XI11_2/XI0/XI0_55/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN0_6 XI11_2/net21_9_ xsel_55_ XI11_2/XI0/XI0_55/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN0_5 XI11_2/net21_10_ xsel_55_ XI11_2/XI0/XI0_55/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN0_4 XI11_2/net21_11_ xsel_55_ XI11_2/XI0/XI0_55/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN0_3 XI11_2/net21_12_ xsel_55_ XI11_2/XI0/XI0_55/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN0_2 XI11_2/net21_13_ xsel_55_ XI11_2/XI0/XI0_55/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN0_1 XI11_2/net21_14_ xsel_55_ XI11_2/XI0/XI0_55/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN0_0 XI11_2/net21_15_ xsel_55_ XI11_2/XI0/XI0_55/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN1_15 XI11_2/XI0/XI0_55/d__15_ xsel_55_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN1_14 XI11_2/XI0/XI0_55/d__14_ xsel_55_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN1_13 XI11_2/XI0/XI0_55/d__13_ xsel_55_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN1_12 XI11_2/XI0/XI0_55/d__12_ xsel_55_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN1_11 XI11_2/XI0/XI0_55/d__11_ xsel_55_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN1_10 XI11_2/XI0/XI0_55/d__10_ xsel_55_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN1_9 XI11_2/XI0/XI0_55/d__9_ xsel_55_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN1_8 XI11_2/XI0/XI0_55/d__8_ xsel_55_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN1_7 XI11_2/XI0/XI0_55/d__7_ xsel_55_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN1_6 XI11_2/XI0/XI0_55/d__6_ xsel_55_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN1_5 XI11_2/XI0/XI0_55/d__5_ xsel_55_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN1_4 XI11_2/XI0/XI0_55/d__4_ xsel_55_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN1_3 XI11_2/XI0/XI0_55/d__3_ xsel_55_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN1_2 XI11_2/XI0/XI0_55/d__2_ xsel_55_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN1_1 XI11_2/XI0/XI0_55/d__1_ xsel_55_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_55/MN1_0 XI11_2/XI0/XI0_55/d__0_ xsel_55_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN0_15 XI11_2/net21_0_ xsel_54_ XI11_2/XI0/XI0_54/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN0_14 XI11_2/net21_1_ xsel_54_ XI11_2/XI0/XI0_54/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN0_13 XI11_2/net21_2_ xsel_54_ XI11_2/XI0/XI0_54/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN0_12 XI11_2/net21_3_ xsel_54_ XI11_2/XI0/XI0_54/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN0_11 XI11_2/net21_4_ xsel_54_ XI11_2/XI0/XI0_54/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN0_10 XI11_2/net21_5_ xsel_54_ XI11_2/XI0/XI0_54/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN0_9 XI11_2/net21_6_ xsel_54_ XI11_2/XI0/XI0_54/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN0_8 XI11_2/net21_7_ xsel_54_ XI11_2/XI0/XI0_54/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN0_7 XI11_2/net21_8_ xsel_54_ XI11_2/XI0/XI0_54/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN0_6 XI11_2/net21_9_ xsel_54_ XI11_2/XI0/XI0_54/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN0_5 XI11_2/net21_10_ xsel_54_ XI11_2/XI0/XI0_54/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN0_4 XI11_2/net21_11_ xsel_54_ XI11_2/XI0/XI0_54/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN0_3 XI11_2/net21_12_ xsel_54_ XI11_2/XI0/XI0_54/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN0_2 XI11_2/net21_13_ xsel_54_ XI11_2/XI0/XI0_54/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN0_1 XI11_2/net21_14_ xsel_54_ XI11_2/XI0/XI0_54/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN0_0 XI11_2/net21_15_ xsel_54_ XI11_2/XI0/XI0_54/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN1_15 XI11_2/XI0/XI0_54/d__15_ xsel_54_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN1_14 XI11_2/XI0/XI0_54/d__14_ xsel_54_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN1_13 XI11_2/XI0/XI0_54/d__13_ xsel_54_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN1_12 XI11_2/XI0/XI0_54/d__12_ xsel_54_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN1_11 XI11_2/XI0/XI0_54/d__11_ xsel_54_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN1_10 XI11_2/XI0/XI0_54/d__10_ xsel_54_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN1_9 XI11_2/XI0/XI0_54/d__9_ xsel_54_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN1_8 XI11_2/XI0/XI0_54/d__8_ xsel_54_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN1_7 XI11_2/XI0/XI0_54/d__7_ xsel_54_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN1_6 XI11_2/XI0/XI0_54/d__6_ xsel_54_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN1_5 XI11_2/XI0/XI0_54/d__5_ xsel_54_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN1_4 XI11_2/XI0/XI0_54/d__4_ xsel_54_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN1_3 XI11_2/XI0/XI0_54/d__3_ xsel_54_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN1_2 XI11_2/XI0/XI0_54/d__2_ xsel_54_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN1_1 XI11_2/XI0/XI0_54/d__1_ xsel_54_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_54/MN1_0 XI11_2/XI0/XI0_54/d__0_ xsel_54_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN0_15 XI11_2/net21_0_ xsel_53_ XI11_2/XI0/XI0_53/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN0_14 XI11_2/net21_1_ xsel_53_ XI11_2/XI0/XI0_53/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN0_13 XI11_2/net21_2_ xsel_53_ XI11_2/XI0/XI0_53/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN0_12 XI11_2/net21_3_ xsel_53_ XI11_2/XI0/XI0_53/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN0_11 XI11_2/net21_4_ xsel_53_ XI11_2/XI0/XI0_53/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN0_10 XI11_2/net21_5_ xsel_53_ XI11_2/XI0/XI0_53/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN0_9 XI11_2/net21_6_ xsel_53_ XI11_2/XI0/XI0_53/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN0_8 XI11_2/net21_7_ xsel_53_ XI11_2/XI0/XI0_53/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN0_7 XI11_2/net21_8_ xsel_53_ XI11_2/XI0/XI0_53/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN0_6 XI11_2/net21_9_ xsel_53_ XI11_2/XI0/XI0_53/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN0_5 XI11_2/net21_10_ xsel_53_ XI11_2/XI0/XI0_53/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN0_4 XI11_2/net21_11_ xsel_53_ XI11_2/XI0/XI0_53/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN0_3 XI11_2/net21_12_ xsel_53_ XI11_2/XI0/XI0_53/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN0_2 XI11_2/net21_13_ xsel_53_ XI11_2/XI0/XI0_53/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN0_1 XI11_2/net21_14_ xsel_53_ XI11_2/XI0/XI0_53/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN0_0 XI11_2/net21_15_ xsel_53_ XI11_2/XI0/XI0_53/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN1_15 XI11_2/XI0/XI0_53/d__15_ xsel_53_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN1_14 XI11_2/XI0/XI0_53/d__14_ xsel_53_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN1_13 XI11_2/XI0/XI0_53/d__13_ xsel_53_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN1_12 XI11_2/XI0/XI0_53/d__12_ xsel_53_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN1_11 XI11_2/XI0/XI0_53/d__11_ xsel_53_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN1_10 XI11_2/XI0/XI0_53/d__10_ xsel_53_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN1_9 XI11_2/XI0/XI0_53/d__9_ xsel_53_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN1_8 XI11_2/XI0/XI0_53/d__8_ xsel_53_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN1_7 XI11_2/XI0/XI0_53/d__7_ xsel_53_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN1_6 XI11_2/XI0/XI0_53/d__6_ xsel_53_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN1_5 XI11_2/XI0/XI0_53/d__5_ xsel_53_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN1_4 XI11_2/XI0/XI0_53/d__4_ xsel_53_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN1_3 XI11_2/XI0/XI0_53/d__3_ xsel_53_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN1_2 XI11_2/XI0/XI0_53/d__2_ xsel_53_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN1_1 XI11_2/XI0/XI0_53/d__1_ xsel_53_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_53/MN1_0 XI11_2/XI0/XI0_53/d__0_ xsel_53_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN0_15 XI11_2/net21_0_ xsel_52_ XI11_2/XI0/XI0_52/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN0_14 XI11_2/net21_1_ xsel_52_ XI11_2/XI0/XI0_52/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN0_13 XI11_2/net21_2_ xsel_52_ XI11_2/XI0/XI0_52/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN0_12 XI11_2/net21_3_ xsel_52_ XI11_2/XI0/XI0_52/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN0_11 XI11_2/net21_4_ xsel_52_ XI11_2/XI0/XI0_52/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN0_10 XI11_2/net21_5_ xsel_52_ XI11_2/XI0/XI0_52/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN0_9 XI11_2/net21_6_ xsel_52_ XI11_2/XI0/XI0_52/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN0_8 XI11_2/net21_7_ xsel_52_ XI11_2/XI0/XI0_52/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN0_7 XI11_2/net21_8_ xsel_52_ XI11_2/XI0/XI0_52/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN0_6 XI11_2/net21_9_ xsel_52_ XI11_2/XI0/XI0_52/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN0_5 XI11_2/net21_10_ xsel_52_ XI11_2/XI0/XI0_52/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN0_4 XI11_2/net21_11_ xsel_52_ XI11_2/XI0/XI0_52/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN0_3 XI11_2/net21_12_ xsel_52_ XI11_2/XI0/XI0_52/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN0_2 XI11_2/net21_13_ xsel_52_ XI11_2/XI0/XI0_52/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN0_1 XI11_2/net21_14_ xsel_52_ XI11_2/XI0/XI0_52/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN0_0 XI11_2/net21_15_ xsel_52_ XI11_2/XI0/XI0_52/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN1_15 XI11_2/XI0/XI0_52/d__15_ xsel_52_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN1_14 XI11_2/XI0/XI0_52/d__14_ xsel_52_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN1_13 XI11_2/XI0/XI0_52/d__13_ xsel_52_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN1_12 XI11_2/XI0/XI0_52/d__12_ xsel_52_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN1_11 XI11_2/XI0/XI0_52/d__11_ xsel_52_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN1_10 XI11_2/XI0/XI0_52/d__10_ xsel_52_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN1_9 XI11_2/XI0/XI0_52/d__9_ xsel_52_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN1_8 XI11_2/XI0/XI0_52/d__8_ xsel_52_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN1_7 XI11_2/XI0/XI0_52/d__7_ xsel_52_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN1_6 XI11_2/XI0/XI0_52/d__6_ xsel_52_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN1_5 XI11_2/XI0/XI0_52/d__5_ xsel_52_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN1_4 XI11_2/XI0/XI0_52/d__4_ xsel_52_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN1_3 XI11_2/XI0/XI0_52/d__3_ xsel_52_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN1_2 XI11_2/XI0/XI0_52/d__2_ xsel_52_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN1_1 XI11_2/XI0/XI0_52/d__1_ xsel_52_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_52/MN1_0 XI11_2/XI0/XI0_52/d__0_ xsel_52_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN0_15 XI11_2/net21_0_ xsel_51_ XI11_2/XI0/XI0_51/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN0_14 XI11_2/net21_1_ xsel_51_ XI11_2/XI0/XI0_51/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN0_13 XI11_2/net21_2_ xsel_51_ XI11_2/XI0/XI0_51/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN0_12 XI11_2/net21_3_ xsel_51_ XI11_2/XI0/XI0_51/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN0_11 XI11_2/net21_4_ xsel_51_ XI11_2/XI0/XI0_51/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN0_10 XI11_2/net21_5_ xsel_51_ XI11_2/XI0/XI0_51/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN0_9 XI11_2/net21_6_ xsel_51_ XI11_2/XI0/XI0_51/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN0_8 XI11_2/net21_7_ xsel_51_ XI11_2/XI0/XI0_51/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN0_7 XI11_2/net21_8_ xsel_51_ XI11_2/XI0/XI0_51/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN0_6 XI11_2/net21_9_ xsel_51_ XI11_2/XI0/XI0_51/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN0_5 XI11_2/net21_10_ xsel_51_ XI11_2/XI0/XI0_51/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN0_4 XI11_2/net21_11_ xsel_51_ XI11_2/XI0/XI0_51/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN0_3 XI11_2/net21_12_ xsel_51_ XI11_2/XI0/XI0_51/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN0_2 XI11_2/net21_13_ xsel_51_ XI11_2/XI0/XI0_51/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN0_1 XI11_2/net21_14_ xsel_51_ XI11_2/XI0/XI0_51/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN0_0 XI11_2/net21_15_ xsel_51_ XI11_2/XI0/XI0_51/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN1_15 XI11_2/XI0/XI0_51/d__15_ xsel_51_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN1_14 XI11_2/XI0/XI0_51/d__14_ xsel_51_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN1_13 XI11_2/XI0/XI0_51/d__13_ xsel_51_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN1_12 XI11_2/XI0/XI0_51/d__12_ xsel_51_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN1_11 XI11_2/XI0/XI0_51/d__11_ xsel_51_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN1_10 XI11_2/XI0/XI0_51/d__10_ xsel_51_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN1_9 XI11_2/XI0/XI0_51/d__9_ xsel_51_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN1_8 XI11_2/XI0/XI0_51/d__8_ xsel_51_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN1_7 XI11_2/XI0/XI0_51/d__7_ xsel_51_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN1_6 XI11_2/XI0/XI0_51/d__6_ xsel_51_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN1_5 XI11_2/XI0/XI0_51/d__5_ xsel_51_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN1_4 XI11_2/XI0/XI0_51/d__4_ xsel_51_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN1_3 XI11_2/XI0/XI0_51/d__3_ xsel_51_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN1_2 XI11_2/XI0/XI0_51/d__2_ xsel_51_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN1_1 XI11_2/XI0/XI0_51/d__1_ xsel_51_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_51/MN1_0 XI11_2/XI0/XI0_51/d__0_ xsel_51_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN0_15 XI11_2/net21_0_ xsel_50_ XI11_2/XI0/XI0_50/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN0_14 XI11_2/net21_1_ xsel_50_ XI11_2/XI0/XI0_50/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN0_13 XI11_2/net21_2_ xsel_50_ XI11_2/XI0/XI0_50/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN0_12 XI11_2/net21_3_ xsel_50_ XI11_2/XI0/XI0_50/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN0_11 XI11_2/net21_4_ xsel_50_ XI11_2/XI0/XI0_50/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN0_10 XI11_2/net21_5_ xsel_50_ XI11_2/XI0/XI0_50/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN0_9 XI11_2/net21_6_ xsel_50_ XI11_2/XI0/XI0_50/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN0_8 XI11_2/net21_7_ xsel_50_ XI11_2/XI0/XI0_50/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN0_7 XI11_2/net21_8_ xsel_50_ XI11_2/XI0/XI0_50/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN0_6 XI11_2/net21_9_ xsel_50_ XI11_2/XI0/XI0_50/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN0_5 XI11_2/net21_10_ xsel_50_ XI11_2/XI0/XI0_50/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN0_4 XI11_2/net21_11_ xsel_50_ XI11_2/XI0/XI0_50/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN0_3 XI11_2/net21_12_ xsel_50_ XI11_2/XI0/XI0_50/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN0_2 XI11_2/net21_13_ xsel_50_ XI11_2/XI0/XI0_50/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN0_1 XI11_2/net21_14_ xsel_50_ XI11_2/XI0/XI0_50/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN0_0 XI11_2/net21_15_ xsel_50_ XI11_2/XI0/XI0_50/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN1_15 XI11_2/XI0/XI0_50/d__15_ xsel_50_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN1_14 XI11_2/XI0/XI0_50/d__14_ xsel_50_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN1_13 XI11_2/XI0/XI0_50/d__13_ xsel_50_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN1_12 XI11_2/XI0/XI0_50/d__12_ xsel_50_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN1_11 XI11_2/XI0/XI0_50/d__11_ xsel_50_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN1_10 XI11_2/XI0/XI0_50/d__10_ xsel_50_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN1_9 XI11_2/XI0/XI0_50/d__9_ xsel_50_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN1_8 XI11_2/XI0/XI0_50/d__8_ xsel_50_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN1_7 XI11_2/XI0/XI0_50/d__7_ xsel_50_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN1_6 XI11_2/XI0/XI0_50/d__6_ xsel_50_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN1_5 XI11_2/XI0/XI0_50/d__5_ xsel_50_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN1_4 XI11_2/XI0/XI0_50/d__4_ xsel_50_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN1_3 XI11_2/XI0/XI0_50/d__3_ xsel_50_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN1_2 XI11_2/XI0/XI0_50/d__2_ xsel_50_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN1_1 XI11_2/XI0/XI0_50/d__1_ xsel_50_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_50/MN1_0 XI11_2/XI0/XI0_50/d__0_ xsel_50_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN0_15 XI11_2/net21_0_ xsel_49_ XI11_2/XI0/XI0_49/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN0_14 XI11_2/net21_1_ xsel_49_ XI11_2/XI0/XI0_49/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN0_13 XI11_2/net21_2_ xsel_49_ XI11_2/XI0/XI0_49/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN0_12 XI11_2/net21_3_ xsel_49_ XI11_2/XI0/XI0_49/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN0_11 XI11_2/net21_4_ xsel_49_ XI11_2/XI0/XI0_49/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN0_10 XI11_2/net21_5_ xsel_49_ XI11_2/XI0/XI0_49/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN0_9 XI11_2/net21_6_ xsel_49_ XI11_2/XI0/XI0_49/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN0_8 XI11_2/net21_7_ xsel_49_ XI11_2/XI0/XI0_49/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN0_7 XI11_2/net21_8_ xsel_49_ XI11_2/XI0/XI0_49/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN0_6 XI11_2/net21_9_ xsel_49_ XI11_2/XI0/XI0_49/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN0_5 XI11_2/net21_10_ xsel_49_ XI11_2/XI0/XI0_49/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN0_4 XI11_2/net21_11_ xsel_49_ XI11_2/XI0/XI0_49/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN0_3 XI11_2/net21_12_ xsel_49_ XI11_2/XI0/XI0_49/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN0_2 XI11_2/net21_13_ xsel_49_ XI11_2/XI0/XI0_49/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN0_1 XI11_2/net21_14_ xsel_49_ XI11_2/XI0/XI0_49/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN0_0 XI11_2/net21_15_ xsel_49_ XI11_2/XI0/XI0_49/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN1_15 XI11_2/XI0/XI0_49/d__15_ xsel_49_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN1_14 XI11_2/XI0/XI0_49/d__14_ xsel_49_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN1_13 XI11_2/XI0/XI0_49/d__13_ xsel_49_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN1_12 XI11_2/XI0/XI0_49/d__12_ xsel_49_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN1_11 XI11_2/XI0/XI0_49/d__11_ xsel_49_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN1_10 XI11_2/XI0/XI0_49/d__10_ xsel_49_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN1_9 XI11_2/XI0/XI0_49/d__9_ xsel_49_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN1_8 XI11_2/XI0/XI0_49/d__8_ xsel_49_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN1_7 XI11_2/XI0/XI0_49/d__7_ xsel_49_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN1_6 XI11_2/XI0/XI0_49/d__6_ xsel_49_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN1_5 XI11_2/XI0/XI0_49/d__5_ xsel_49_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN1_4 XI11_2/XI0/XI0_49/d__4_ xsel_49_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN1_3 XI11_2/XI0/XI0_49/d__3_ xsel_49_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN1_2 XI11_2/XI0/XI0_49/d__2_ xsel_49_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN1_1 XI11_2/XI0/XI0_49/d__1_ xsel_49_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_49/MN1_0 XI11_2/XI0/XI0_49/d__0_ xsel_49_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN0_15 XI11_2/net21_0_ xsel_48_ XI11_2/XI0/XI0_48/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN0_14 XI11_2/net21_1_ xsel_48_ XI11_2/XI0/XI0_48/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN0_13 XI11_2/net21_2_ xsel_48_ XI11_2/XI0/XI0_48/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN0_12 XI11_2/net21_3_ xsel_48_ XI11_2/XI0/XI0_48/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN0_11 XI11_2/net21_4_ xsel_48_ XI11_2/XI0/XI0_48/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN0_10 XI11_2/net21_5_ xsel_48_ XI11_2/XI0/XI0_48/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN0_9 XI11_2/net21_6_ xsel_48_ XI11_2/XI0/XI0_48/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN0_8 XI11_2/net21_7_ xsel_48_ XI11_2/XI0/XI0_48/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN0_7 XI11_2/net21_8_ xsel_48_ XI11_2/XI0/XI0_48/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN0_6 XI11_2/net21_9_ xsel_48_ XI11_2/XI0/XI0_48/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN0_5 XI11_2/net21_10_ xsel_48_ XI11_2/XI0/XI0_48/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN0_4 XI11_2/net21_11_ xsel_48_ XI11_2/XI0/XI0_48/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN0_3 XI11_2/net21_12_ xsel_48_ XI11_2/XI0/XI0_48/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN0_2 XI11_2/net21_13_ xsel_48_ XI11_2/XI0/XI0_48/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN0_1 XI11_2/net21_14_ xsel_48_ XI11_2/XI0/XI0_48/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN0_0 XI11_2/net21_15_ xsel_48_ XI11_2/XI0/XI0_48/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN1_15 XI11_2/XI0/XI0_48/d__15_ xsel_48_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN1_14 XI11_2/XI0/XI0_48/d__14_ xsel_48_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN1_13 XI11_2/XI0/XI0_48/d__13_ xsel_48_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN1_12 XI11_2/XI0/XI0_48/d__12_ xsel_48_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN1_11 XI11_2/XI0/XI0_48/d__11_ xsel_48_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN1_10 XI11_2/XI0/XI0_48/d__10_ xsel_48_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN1_9 XI11_2/XI0/XI0_48/d__9_ xsel_48_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN1_8 XI11_2/XI0/XI0_48/d__8_ xsel_48_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN1_7 XI11_2/XI0/XI0_48/d__7_ xsel_48_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN1_6 XI11_2/XI0/XI0_48/d__6_ xsel_48_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN1_5 XI11_2/XI0/XI0_48/d__5_ xsel_48_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN1_4 XI11_2/XI0/XI0_48/d__4_ xsel_48_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN1_3 XI11_2/XI0/XI0_48/d__3_ xsel_48_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN1_2 XI11_2/XI0/XI0_48/d__2_ xsel_48_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN1_1 XI11_2/XI0/XI0_48/d__1_ xsel_48_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_48/MN1_0 XI11_2/XI0/XI0_48/d__0_ xsel_48_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN0_15 XI11_2/net21_0_ xsel_47_ XI11_2/XI0/XI0_47/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN0_14 XI11_2/net21_1_ xsel_47_ XI11_2/XI0/XI0_47/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN0_13 XI11_2/net21_2_ xsel_47_ XI11_2/XI0/XI0_47/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN0_12 XI11_2/net21_3_ xsel_47_ XI11_2/XI0/XI0_47/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN0_11 XI11_2/net21_4_ xsel_47_ XI11_2/XI0/XI0_47/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN0_10 XI11_2/net21_5_ xsel_47_ XI11_2/XI0/XI0_47/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN0_9 XI11_2/net21_6_ xsel_47_ XI11_2/XI0/XI0_47/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN0_8 XI11_2/net21_7_ xsel_47_ XI11_2/XI0/XI0_47/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN0_7 XI11_2/net21_8_ xsel_47_ XI11_2/XI0/XI0_47/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN0_6 XI11_2/net21_9_ xsel_47_ XI11_2/XI0/XI0_47/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN0_5 XI11_2/net21_10_ xsel_47_ XI11_2/XI0/XI0_47/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN0_4 XI11_2/net21_11_ xsel_47_ XI11_2/XI0/XI0_47/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN0_3 XI11_2/net21_12_ xsel_47_ XI11_2/XI0/XI0_47/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN0_2 XI11_2/net21_13_ xsel_47_ XI11_2/XI0/XI0_47/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN0_1 XI11_2/net21_14_ xsel_47_ XI11_2/XI0/XI0_47/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN0_0 XI11_2/net21_15_ xsel_47_ XI11_2/XI0/XI0_47/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN1_15 XI11_2/XI0/XI0_47/d__15_ xsel_47_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN1_14 XI11_2/XI0/XI0_47/d__14_ xsel_47_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN1_13 XI11_2/XI0/XI0_47/d__13_ xsel_47_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN1_12 XI11_2/XI0/XI0_47/d__12_ xsel_47_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN1_11 XI11_2/XI0/XI0_47/d__11_ xsel_47_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN1_10 XI11_2/XI0/XI0_47/d__10_ xsel_47_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN1_9 XI11_2/XI0/XI0_47/d__9_ xsel_47_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN1_8 XI11_2/XI0/XI0_47/d__8_ xsel_47_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN1_7 XI11_2/XI0/XI0_47/d__7_ xsel_47_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN1_6 XI11_2/XI0/XI0_47/d__6_ xsel_47_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN1_5 XI11_2/XI0/XI0_47/d__5_ xsel_47_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN1_4 XI11_2/XI0/XI0_47/d__4_ xsel_47_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN1_3 XI11_2/XI0/XI0_47/d__3_ xsel_47_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN1_2 XI11_2/XI0/XI0_47/d__2_ xsel_47_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN1_1 XI11_2/XI0/XI0_47/d__1_ xsel_47_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_47/MN1_0 XI11_2/XI0/XI0_47/d__0_ xsel_47_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN0_15 XI11_2/net21_0_ xsel_46_ XI11_2/XI0/XI0_46/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN0_14 XI11_2/net21_1_ xsel_46_ XI11_2/XI0/XI0_46/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN0_13 XI11_2/net21_2_ xsel_46_ XI11_2/XI0/XI0_46/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN0_12 XI11_2/net21_3_ xsel_46_ XI11_2/XI0/XI0_46/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN0_11 XI11_2/net21_4_ xsel_46_ XI11_2/XI0/XI0_46/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN0_10 XI11_2/net21_5_ xsel_46_ XI11_2/XI0/XI0_46/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN0_9 XI11_2/net21_6_ xsel_46_ XI11_2/XI0/XI0_46/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN0_8 XI11_2/net21_7_ xsel_46_ XI11_2/XI0/XI0_46/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN0_7 XI11_2/net21_8_ xsel_46_ XI11_2/XI0/XI0_46/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN0_6 XI11_2/net21_9_ xsel_46_ XI11_2/XI0/XI0_46/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN0_5 XI11_2/net21_10_ xsel_46_ XI11_2/XI0/XI0_46/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN0_4 XI11_2/net21_11_ xsel_46_ XI11_2/XI0/XI0_46/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN0_3 XI11_2/net21_12_ xsel_46_ XI11_2/XI0/XI0_46/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN0_2 XI11_2/net21_13_ xsel_46_ XI11_2/XI0/XI0_46/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN0_1 XI11_2/net21_14_ xsel_46_ XI11_2/XI0/XI0_46/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN0_0 XI11_2/net21_15_ xsel_46_ XI11_2/XI0/XI0_46/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN1_15 XI11_2/XI0/XI0_46/d__15_ xsel_46_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN1_14 XI11_2/XI0/XI0_46/d__14_ xsel_46_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN1_13 XI11_2/XI0/XI0_46/d__13_ xsel_46_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN1_12 XI11_2/XI0/XI0_46/d__12_ xsel_46_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN1_11 XI11_2/XI0/XI0_46/d__11_ xsel_46_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN1_10 XI11_2/XI0/XI0_46/d__10_ xsel_46_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN1_9 XI11_2/XI0/XI0_46/d__9_ xsel_46_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN1_8 XI11_2/XI0/XI0_46/d__8_ xsel_46_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN1_7 XI11_2/XI0/XI0_46/d__7_ xsel_46_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN1_6 XI11_2/XI0/XI0_46/d__6_ xsel_46_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN1_5 XI11_2/XI0/XI0_46/d__5_ xsel_46_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN1_4 XI11_2/XI0/XI0_46/d__4_ xsel_46_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN1_3 XI11_2/XI0/XI0_46/d__3_ xsel_46_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN1_2 XI11_2/XI0/XI0_46/d__2_ xsel_46_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN1_1 XI11_2/XI0/XI0_46/d__1_ xsel_46_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_46/MN1_0 XI11_2/XI0/XI0_46/d__0_ xsel_46_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN0_15 XI11_2/net21_0_ xsel_45_ XI11_2/XI0/XI0_45/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN0_14 XI11_2/net21_1_ xsel_45_ XI11_2/XI0/XI0_45/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN0_13 XI11_2/net21_2_ xsel_45_ XI11_2/XI0/XI0_45/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN0_12 XI11_2/net21_3_ xsel_45_ XI11_2/XI0/XI0_45/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN0_11 XI11_2/net21_4_ xsel_45_ XI11_2/XI0/XI0_45/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN0_10 XI11_2/net21_5_ xsel_45_ XI11_2/XI0/XI0_45/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN0_9 XI11_2/net21_6_ xsel_45_ XI11_2/XI0/XI0_45/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN0_8 XI11_2/net21_7_ xsel_45_ XI11_2/XI0/XI0_45/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN0_7 XI11_2/net21_8_ xsel_45_ XI11_2/XI0/XI0_45/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN0_6 XI11_2/net21_9_ xsel_45_ XI11_2/XI0/XI0_45/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN0_5 XI11_2/net21_10_ xsel_45_ XI11_2/XI0/XI0_45/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN0_4 XI11_2/net21_11_ xsel_45_ XI11_2/XI0/XI0_45/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN0_3 XI11_2/net21_12_ xsel_45_ XI11_2/XI0/XI0_45/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN0_2 XI11_2/net21_13_ xsel_45_ XI11_2/XI0/XI0_45/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN0_1 XI11_2/net21_14_ xsel_45_ XI11_2/XI0/XI0_45/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN0_0 XI11_2/net21_15_ xsel_45_ XI11_2/XI0/XI0_45/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN1_15 XI11_2/XI0/XI0_45/d__15_ xsel_45_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN1_14 XI11_2/XI0/XI0_45/d__14_ xsel_45_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN1_13 XI11_2/XI0/XI0_45/d__13_ xsel_45_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN1_12 XI11_2/XI0/XI0_45/d__12_ xsel_45_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN1_11 XI11_2/XI0/XI0_45/d__11_ xsel_45_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN1_10 XI11_2/XI0/XI0_45/d__10_ xsel_45_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN1_9 XI11_2/XI0/XI0_45/d__9_ xsel_45_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN1_8 XI11_2/XI0/XI0_45/d__8_ xsel_45_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN1_7 XI11_2/XI0/XI0_45/d__7_ xsel_45_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN1_6 XI11_2/XI0/XI0_45/d__6_ xsel_45_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN1_5 XI11_2/XI0/XI0_45/d__5_ xsel_45_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN1_4 XI11_2/XI0/XI0_45/d__4_ xsel_45_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN1_3 XI11_2/XI0/XI0_45/d__3_ xsel_45_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN1_2 XI11_2/XI0/XI0_45/d__2_ xsel_45_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN1_1 XI11_2/XI0/XI0_45/d__1_ xsel_45_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_45/MN1_0 XI11_2/XI0/XI0_45/d__0_ xsel_45_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN0_15 XI11_2/net21_0_ xsel_44_ XI11_2/XI0/XI0_44/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN0_14 XI11_2/net21_1_ xsel_44_ XI11_2/XI0/XI0_44/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN0_13 XI11_2/net21_2_ xsel_44_ XI11_2/XI0/XI0_44/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN0_12 XI11_2/net21_3_ xsel_44_ XI11_2/XI0/XI0_44/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN0_11 XI11_2/net21_4_ xsel_44_ XI11_2/XI0/XI0_44/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN0_10 XI11_2/net21_5_ xsel_44_ XI11_2/XI0/XI0_44/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN0_9 XI11_2/net21_6_ xsel_44_ XI11_2/XI0/XI0_44/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN0_8 XI11_2/net21_7_ xsel_44_ XI11_2/XI0/XI0_44/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN0_7 XI11_2/net21_8_ xsel_44_ XI11_2/XI0/XI0_44/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN0_6 XI11_2/net21_9_ xsel_44_ XI11_2/XI0/XI0_44/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN0_5 XI11_2/net21_10_ xsel_44_ XI11_2/XI0/XI0_44/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN0_4 XI11_2/net21_11_ xsel_44_ XI11_2/XI0/XI0_44/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN0_3 XI11_2/net21_12_ xsel_44_ XI11_2/XI0/XI0_44/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN0_2 XI11_2/net21_13_ xsel_44_ XI11_2/XI0/XI0_44/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN0_1 XI11_2/net21_14_ xsel_44_ XI11_2/XI0/XI0_44/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN0_0 XI11_2/net21_15_ xsel_44_ XI11_2/XI0/XI0_44/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN1_15 XI11_2/XI0/XI0_44/d__15_ xsel_44_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN1_14 XI11_2/XI0/XI0_44/d__14_ xsel_44_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN1_13 XI11_2/XI0/XI0_44/d__13_ xsel_44_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN1_12 XI11_2/XI0/XI0_44/d__12_ xsel_44_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN1_11 XI11_2/XI0/XI0_44/d__11_ xsel_44_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN1_10 XI11_2/XI0/XI0_44/d__10_ xsel_44_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN1_9 XI11_2/XI0/XI0_44/d__9_ xsel_44_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN1_8 XI11_2/XI0/XI0_44/d__8_ xsel_44_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN1_7 XI11_2/XI0/XI0_44/d__7_ xsel_44_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN1_6 XI11_2/XI0/XI0_44/d__6_ xsel_44_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN1_5 XI11_2/XI0/XI0_44/d__5_ xsel_44_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN1_4 XI11_2/XI0/XI0_44/d__4_ xsel_44_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN1_3 XI11_2/XI0/XI0_44/d__3_ xsel_44_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN1_2 XI11_2/XI0/XI0_44/d__2_ xsel_44_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN1_1 XI11_2/XI0/XI0_44/d__1_ xsel_44_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_44/MN1_0 XI11_2/XI0/XI0_44/d__0_ xsel_44_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN0_15 XI11_2/net21_0_ xsel_43_ XI11_2/XI0/XI0_43/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN0_14 XI11_2/net21_1_ xsel_43_ XI11_2/XI0/XI0_43/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN0_13 XI11_2/net21_2_ xsel_43_ XI11_2/XI0/XI0_43/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN0_12 XI11_2/net21_3_ xsel_43_ XI11_2/XI0/XI0_43/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN0_11 XI11_2/net21_4_ xsel_43_ XI11_2/XI0/XI0_43/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN0_10 XI11_2/net21_5_ xsel_43_ XI11_2/XI0/XI0_43/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN0_9 XI11_2/net21_6_ xsel_43_ XI11_2/XI0/XI0_43/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN0_8 XI11_2/net21_7_ xsel_43_ XI11_2/XI0/XI0_43/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN0_7 XI11_2/net21_8_ xsel_43_ XI11_2/XI0/XI0_43/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN0_6 XI11_2/net21_9_ xsel_43_ XI11_2/XI0/XI0_43/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN0_5 XI11_2/net21_10_ xsel_43_ XI11_2/XI0/XI0_43/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN0_4 XI11_2/net21_11_ xsel_43_ XI11_2/XI0/XI0_43/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN0_3 XI11_2/net21_12_ xsel_43_ XI11_2/XI0/XI0_43/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN0_2 XI11_2/net21_13_ xsel_43_ XI11_2/XI0/XI0_43/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN0_1 XI11_2/net21_14_ xsel_43_ XI11_2/XI0/XI0_43/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN0_0 XI11_2/net21_15_ xsel_43_ XI11_2/XI0/XI0_43/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN1_15 XI11_2/XI0/XI0_43/d__15_ xsel_43_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN1_14 XI11_2/XI0/XI0_43/d__14_ xsel_43_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN1_13 XI11_2/XI0/XI0_43/d__13_ xsel_43_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN1_12 XI11_2/XI0/XI0_43/d__12_ xsel_43_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN1_11 XI11_2/XI0/XI0_43/d__11_ xsel_43_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN1_10 XI11_2/XI0/XI0_43/d__10_ xsel_43_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN1_9 XI11_2/XI0/XI0_43/d__9_ xsel_43_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN1_8 XI11_2/XI0/XI0_43/d__8_ xsel_43_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN1_7 XI11_2/XI0/XI0_43/d__7_ xsel_43_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN1_6 XI11_2/XI0/XI0_43/d__6_ xsel_43_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN1_5 XI11_2/XI0/XI0_43/d__5_ xsel_43_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN1_4 XI11_2/XI0/XI0_43/d__4_ xsel_43_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN1_3 XI11_2/XI0/XI0_43/d__3_ xsel_43_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN1_2 XI11_2/XI0/XI0_43/d__2_ xsel_43_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN1_1 XI11_2/XI0/XI0_43/d__1_ xsel_43_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_43/MN1_0 XI11_2/XI0/XI0_43/d__0_ xsel_43_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN0_15 XI11_2/net21_0_ xsel_42_ XI11_2/XI0/XI0_42/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN0_14 XI11_2/net21_1_ xsel_42_ XI11_2/XI0/XI0_42/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN0_13 XI11_2/net21_2_ xsel_42_ XI11_2/XI0/XI0_42/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN0_12 XI11_2/net21_3_ xsel_42_ XI11_2/XI0/XI0_42/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN0_11 XI11_2/net21_4_ xsel_42_ XI11_2/XI0/XI0_42/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN0_10 XI11_2/net21_5_ xsel_42_ XI11_2/XI0/XI0_42/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN0_9 XI11_2/net21_6_ xsel_42_ XI11_2/XI0/XI0_42/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN0_8 XI11_2/net21_7_ xsel_42_ XI11_2/XI0/XI0_42/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN0_7 XI11_2/net21_8_ xsel_42_ XI11_2/XI0/XI0_42/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN0_6 XI11_2/net21_9_ xsel_42_ XI11_2/XI0/XI0_42/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN0_5 XI11_2/net21_10_ xsel_42_ XI11_2/XI0/XI0_42/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN0_4 XI11_2/net21_11_ xsel_42_ XI11_2/XI0/XI0_42/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN0_3 XI11_2/net21_12_ xsel_42_ XI11_2/XI0/XI0_42/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN0_2 XI11_2/net21_13_ xsel_42_ XI11_2/XI0/XI0_42/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN0_1 XI11_2/net21_14_ xsel_42_ XI11_2/XI0/XI0_42/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN0_0 XI11_2/net21_15_ xsel_42_ XI11_2/XI0/XI0_42/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN1_15 XI11_2/XI0/XI0_42/d__15_ xsel_42_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN1_14 XI11_2/XI0/XI0_42/d__14_ xsel_42_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN1_13 XI11_2/XI0/XI0_42/d__13_ xsel_42_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN1_12 XI11_2/XI0/XI0_42/d__12_ xsel_42_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN1_11 XI11_2/XI0/XI0_42/d__11_ xsel_42_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN1_10 XI11_2/XI0/XI0_42/d__10_ xsel_42_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN1_9 XI11_2/XI0/XI0_42/d__9_ xsel_42_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN1_8 XI11_2/XI0/XI0_42/d__8_ xsel_42_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN1_7 XI11_2/XI0/XI0_42/d__7_ xsel_42_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN1_6 XI11_2/XI0/XI0_42/d__6_ xsel_42_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN1_5 XI11_2/XI0/XI0_42/d__5_ xsel_42_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN1_4 XI11_2/XI0/XI0_42/d__4_ xsel_42_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN1_3 XI11_2/XI0/XI0_42/d__3_ xsel_42_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN1_2 XI11_2/XI0/XI0_42/d__2_ xsel_42_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN1_1 XI11_2/XI0/XI0_42/d__1_ xsel_42_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_42/MN1_0 XI11_2/XI0/XI0_42/d__0_ xsel_42_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN0_15 XI11_2/net21_0_ xsel_41_ XI11_2/XI0/XI0_41/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN0_14 XI11_2/net21_1_ xsel_41_ XI11_2/XI0/XI0_41/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN0_13 XI11_2/net21_2_ xsel_41_ XI11_2/XI0/XI0_41/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN0_12 XI11_2/net21_3_ xsel_41_ XI11_2/XI0/XI0_41/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN0_11 XI11_2/net21_4_ xsel_41_ XI11_2/XI0/XI0_41/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN0_10 XI11_2/net21_5_ xsel_41_ XI11_2/XI0/XI0_41/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN0_9 XI11_2/net21_6_ xsel_41_ XI11_2/XI0/XI0_41/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN0_8 XI11_2/net21_7_ xsel_41_ XI11_2/XI0/XI0_41/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN0_7 XI11_2/net21_8_ xsel_41_ XI11_2/XI0/XI0_41/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN0_6 XI11_2/net21_9_ xsel_41_ XI11_2/XI0/XI0_41/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN0_5 XI11_2/net21_10_ xsel_41_ XI11_2/XI0/XI0_41/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN0_4 XI11_2/net21_11_ xsel_41_ XI11_2/XI0/XI0_41/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN0_3 XI11_2/net21_12_ xsel_41_ XI11_2/XI0/XI0_41/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN0_2 XI11_2/net21_13_ xsel_41_ XI11_2/XI0/XI0_41/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN0_1 XI11_2/net21_14_ xsel_41_ XI11_2/XI0/XI0_41/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN0_0 XI11_2/net21_15_ xsel_41_ XI11_2/XI0/XI0_41/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN1_15 XI11_2/XI0/XI0_41/d__15_ xsel_41_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN1_14 XI11_2/XI0/XI0_41/d__14_ xsel_41_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN1_13 XI11_2/XI0/XI0_41/d__13_ xsel_41_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN1_12 XI11_2/XI0/XI0_41/d__12_ xsel_41_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN1_11 XI11_2/XI0/XI0_41/d__11_ xsel_41_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN1_10 XI11_2/XI0/XI0_41/d__10_ xsel_41_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN1_9 XI11_2/XI0/XI0_41/d__9_ xsel_41_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN1_8 XI11_2/XI0/XI0_41/d__8_ xsel_41_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN1_7 XI11_2/XI0/XI0_41/d__7_ xsel_41_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN1_6 XI11_2/XI0/XI0_41/d__6_ xsel_41_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN1_5 XI11_2/XI0/XI0_41/d__5_ xsel_41_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN1_4 XI11_2/XI0/XI0_41/d__4_ xsel_41_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN1_3 XI11_2/XI0/XI0_41/d__3_ xsel_41_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN1_2 XI11_2/XI0/XI0_41/d__2_ xsel_41_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN1_1 XI11_2/XI0/XI0_41/d__1_ xsel_41_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_41/MN1_0 XI11_2/XI0/XI0_41/d__0_ xsel_41_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN0_15 XI11_2/net21_0_ xsel_40_ XI11_2/XI0/XI0_40/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN0_14 XI11_2/net21_1_ xsel_40_ XI11_2/XI0/XI0_40/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN0_13 XI11_2/net21_2_ xsel_40_ XI11_2/XI0/XI0_40/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN0_12 XI11_2/net21_3_ xsel_40_ XI11_2/XI0/XI0_40/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN0_11 XI11_2/net21_4_ xsel_40_ XI11_2/XI0/XI0_40/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN0_10 XI11_2/net21_5_ xsel_40_ XI11_2/XI0/XI0_40/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN0_9 XI11_2/net21_6_ xsel_40_ XI11_2/XI0/XI0_40/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN0_8 XI11_2/net21_7_ xsel_40_ XI11_2/XI0/XI0_40/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN0_7 XI11_2/net21_8_ xsel_40_ XI11_2/XI0/XI0_40/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN0_6 XI11_2/net21_9_ xsel_40_ XI11_2/XI0/XI0_40/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN0_5 XI11_2/net21_10_ xsel_40_ XI11_2/XI0/XI0_40/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN0_4 XI11_2/net21_11_ xsel_40_ XI11_2/XI0/XI0_40/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN0_3 XI11_2/net21_12_ xsel_40_ XI11_2/XI0/XI0_40/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN0_2 XI11_2/net21_13_ xsel_40_ XI11_2/XI0/XI0_40/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN0_1 XI11_2/net21_14_ xsel_40_ XI11_2/XI0/XI0_40/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN0_0 XI11_2/net21_15_ xsel_40_ XI11_2/XI0/XI0_40/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN1_15 XI11_2/XI0/XI0_40/d__15_ xsel_40_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN1_14 XI11_2/XI0/XI0_40/d__14_ xsel_40_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN1_13 XI11_2/XI0/XI0_40/d__13_ xsel_40_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN1_12 XI11_2/XI0/XI0_40/d__12_ xsel_40_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN1_11 XI11_2/XI0/XI0_40/d__11_ xsel_40_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN1_10 XI11_2/XI0/XI0_40/d__10_ xsel_40_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN1_9 XI11_2/XI0/XI0_40/d__9_ xsel_40_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN1_8 XI11_2/XI0/XI0_40/d__8_ xsel_40_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN1_7 XI11_2/XI0/XI0_40/d__7_ xsel_40_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN1_6 XI11_2/XI0/XI0_40/d__6_ xsel_40_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN1_5 XI11_2/XI0/XI0_40/d__5_ xsel_40_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN1_4 XI11_2/XI0/XI0_40/d__4_ xsel_40_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN1_3 XI11_2/XI0/XI0_40/d__3_ xsel_40_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN1_2 XI11_2/XI0/XI0_40/d__2_ xsel_40_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN1_1 XI11_2/XI0/XI0_40/d__1_ xsel_40_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_40/MN1_0 XI11_2/XI0/XI0_40/d__0_ xsel_40_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN0_15 XI11_2/net21_0_ xsel_39_ XI11_2/XI0/XI0_39/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN0_14 XI11_2/net21_1_ xsel_39_ XI11_2/XI0/XI0_39/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN0_13 XI11_2/net21_2_ xsel_39_ XI11_2/XI0/XI0_39/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN0_12 XI11_2/net21_3_ xsel_39_ XI11_2/XI0/XI0_39/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN0_11 XI11_2/net21_4_ xsel_39_ XI11_2/XI0/XI0_39/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN0_10 XI11_2/net21_5_ xsel_39_ XI11_2/XI0/XI0_39/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN0_9 XI11_2/net21_6_ xsel_39_ XI11_2/XI0/XI0_39/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN0_8 XI11_2/net21_7_ xsel_39_ XI11_2/XI0/XI0_39/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN0_7 XI11_2/net21_8_ xsel_39_ XI11_2/XI0/XI0_39/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN0_6 XI11_2/net21_9_ xsel_39_ XI11_2/XI0/XI0_39/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN0_5 XI11_2/net21_10_ xsel_39_ XI11_2/XI0/XI0_39/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN0_4 XI11_2/net21_11_ xsel_39_ XI11_2/XI0/XI0_39/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN0_3 XI11_2/net21_12_ xsel_39_ XI11_2/XI0/XI0_39/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN0_2 XI11_2/net21_13_ xsel_39_ XI11_2/XI0/XI0_39/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN0_1 XI11_2/net21_14_ xsel_39_ XI11_2/XI0/XI0_39/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN0_0 XI11_2/net21_15_ xsel_39_ XI11_2/XI0/XI0_39/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN1_15 XI11_2/XI0/XI0_39/d__15_ xsel_39_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN1_14 XI11_2/XI0/XI0_39/d__14_ xsel_39_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN1_13 XI11_2/XI0/XI0_39/d__13_ xsel_39_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN1_12 XI11_2/XI0/XI0_39/d__12_ xsel_39_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN1_11 XI11_2/XI0/XI0_39/d__11_ xsel_39_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN1_10 XI11_2/XI0/XI0_39/d__10_ xsel_39_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN1_9 XI11_2/XI0/XI0_39/d__9_ xsel_39_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN1_8 XI11_2/XI0/XI0_39/d__8_ xsel_39_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN1_7 XI11_2/XI0/XI0_39/d__7_ xsel_39_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN1_6 XI11_2/XI0/XI0_39/d__6_ xsel_39_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN1_5 XI11_2/XI0/XI0_39/d__5_ xsel_39_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN1_4 XI11_2/XI0/XI0_39/d__4_ xsel_39_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN1_3 XI11_2/XI0/XI0_39/d__3_ xsel_39_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN1_2 XI11_2/XI0/XI0_39/d__2_ xsel_39_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN1_1 XI11_2/XI0/XI0_39/d__1_ xsel_39_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_39/MN1_0 XI11_2/XI0/XI0_39/d__0_ xsel_39_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN0_15 XI11_2/net21_0_ xsel_38_ XI11_2/XI0/XI0_38/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN0_14 XI11_2/net21_1_ xsel_38_ XI11_2/XI0/XI0_38/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN0_13 XI11_2/net21_2_ xsel_38_ XI11_2/XI0/XI0_38/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN0_12 XI11_2/net21_3_ xsel_38_ XI11_2/XI0/XI0_38/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN0_11 XI11_2/net21_4_ xsel_38_ XI11_2/XI0/XI0_38/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN0_10 XI11_2/net21_5_ xsel_38_ XI11_2/XI0/XI0_38/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN0_9 XI11_2/net21_6_ xsel_38_ XI11_2/XI0/XI0_38/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN0_8 XI11_2/net21_7_ xsel_38_ XI11_2/XI0/XI0_38/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN0_7 XI11_2/net21_8_ xsel_38_ XI11_2/XI0/XI0_38/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN0_6 XI11_2/net21_9_ xsel_38_ XI11_2/XI0/XI0_38/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN0_5 XI11_2/net21_10_ xsel_38_ XI11_2/XI0/XI0_38/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN0_4 XI11_2/net21_11_ xsel_38_ XI11_2/XI0/XI0_38/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN0_3 XI11_2/net21_12_ xsel_38_ XI11_2/XI0/XI0_38/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN0_2 XI11_2/net21_13_ xsel_38_ XI11_2/XI0/XI0_38/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN0_1 XI11_2/net21_14_ xsel_38_ XI11_2/XI0/XI0_38/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN0_0 XI11_2/net21_15_ xsel_38_ XI11_2/XI0/XI0_38/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN1_15 XI11_2/XI0/XI0_38/d__15_ xsel_38_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN1_14 XI11_2/XI0/XI0_38/d__14_ xsel_38_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN1_13 XI11_2/XI0/XI0_38/d__13_ xsel_38_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN1_12 XI11_2/XI0/XI0_38/d__12_ xsel_38_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN1_11 XI11_2/XI0/XI0_38/d__11_ xsel_38_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN1_10 XI11_2/XI0/XI0_38/d__10_ xsel_38_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN1_9 XI11_2/XI0/XI0_38/d__9_ xsel_38_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN1_8 XI11_2/XI0/XI0_38/d__8_ xsel_38_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN1_7 XI11_2/XI0/XI0_38/d__7_ xsel_38_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN1_6 XI11_2/XI0/XI0_38/d__6_ xsel_38_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN1_5 XI11_2/XI0/XI0_38/d__5_ xsel_38_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN1_4 XI11_2/XI0/XI0_38/d__4_ xsel_38_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN1_3 XI11_2/XI0/XI0_38/d__3_ xsel_38_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN1_2 XI11_2/XI0/XI0_38/d__2_ xsel_38_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN1_1 XI11_2/XI0/XI0_38/d__1_ xsel_38_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_38/MN1_0 XI11_2/XI0/XI0_38/d__0_ xsel_38_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN0_15 XI11_2/net21_0_ xsel_37_ XI11_2/XI0/XI0_37/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN0_14 XI11_2/net21_1_ xsel_37_ XI11_2/XI0/XI0_37/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN0_13 XI11_2/net21_2_ xsel_37_ XI11_2/XI0/XI0_37/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN0_12 XI11_2/net21_3_ xsel_37_ XI11_2/XI0/XI0_37/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN0_11 XI11_2/net21_4_ xsel_37_ XI11_2/XI0/XI0_37/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN0_10 XI11_2/net21_5_ xsel_37_ XI11_2/XI0/XI0_37/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN0_9 XI11_2/net21_6_ xsel_37_ XI11_2/XI0/XI0_37/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN0_8 XI11_2/net21_7_ xsel_37_ XI11_2/XI0/XI0_37/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN0_7 XI11_2/net21_8_ xsel_37_ XI11_2/XI0/XI0_37/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN0_6 XI11_2/net21_9_ xsel_37_ XI11_2/XI0/XI0_37/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN0_5 XI11_2/net21_10_ xsel_37_ XI11_2/XI0/XI0_37/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN0_4 XI11_2/net21_11_ xsel_37_ XI11_2/XI0/XI0_37/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN0_3 XI11_2/net21_12_ xsel_37_ XI11_2/XI0/XI0_37/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN0_2 XI11_2/net21_13_ xsel_37_ XI11_2/XI0/XI0_37/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN0_1 XI11_2/net21_14_ xsel_37_ XI11_2/XI0/XI0_37/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN0_0 XI11_2/net21_15_ xsel_37_ XI11_2/XI0/XI0_37/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN1_15 XI11_2/XI0/XI0_37/d__15_ xsel_37_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN1_14 XI11_2/XI0/XI0_37/d__14_ xsel_37_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN1_13 XI11_2/XI0/XI0_37/d__13_ xsel_37_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN1_12 XI11_2/XI0/XI0_37/d__12_ xsel_37_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN1_11 XI11_2/XI0/XI0_37/d__11_ xsel_37_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN1_10 XI11_2/XI0/XI0_37/d__10_ xsel_37_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN1_9 XI11_2/XI0/XI0_37/d__9_ xsel_37_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN1_8 XI11_2/XI0/XI0_37/d__8_ xsel_37_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN1_7 XI11_2/XI0/XI0_37/d__7_ xsel_37_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN1_6 XI11_2/XI0/XI0_37/d__6_ xsel_37_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN1_5 XI11_2/XI0/XI0_37/d__5_ xsel_37_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN1_4 XI11_2/XI0/XI0_37/d__4_ xsel_37_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN1_3 XI11_2/XI0/XI0_37/d__3_ xsel_37_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN1_2 XI11_2/XI0/XI0_37/d__2_ xsel_37_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN1_1 XI11_2/XI0/XI0_37/d__1_ xsel_37_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_37/MN1_0 XI11_2/XI0/XI0_37/d__0_ xsel_37_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN0_15 XI11_2/net21_0_ xsel_36_ XI11_2/XI0/XI0_36/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN0_14 XI11_2/net21_1_ xsel_36_ XI11_2/XI0/XI0_36/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN0_13 XI11_2/net21_2_ xsel_36_ XI11_2/XI0/XI0_36/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN0_12 XI11_2/net21_3_ xsel_36_ XI11_2/XI0/XI0_36/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN0_11 XI11_2/net21_4_ xsel_36_ XI11_2/XI0/XI0_36/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN0_10 XI11_2/net21_5_ xsel_36_ XI11_2/XI0/XI0_36/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN0_9 XI11_2/net21_6_ xsel_36_ XI11_2/XI0/XI0_36/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN0_8 XI11_2/net21_7_ xsel_36_ XI11_2/XI0/XI0_36/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN0_7 XI11_2/net21_8_ xsel_36_ XI11_2/XI0/XI0_36/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN0_6 XI11_2/net21_9_ xsel_36_ XI11_2/XI0/XI0_36/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN0_5 XI11_2/net21_10_ xsel_36_ XI11_2/XI0/XI0_36/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN0_4 XI11_2/net21_11_ xsel_36_ XI11_2/XI0/XI0_36/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN0_3 XI11_2/net21_12_ xsel_36_ XI11_2/XI0/XI0_36/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN0_2 XI11_2/net21_13_ xsel_36_ XI11_2/XI0/XI0_36/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN0_1 XI11_2/net21_14_ xsel_36_ XI11_2/XI0/XI0_36/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN0_0 XI11_2/net21_15_ xsel_36_ XI11_2/XI0/XI0_36/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN1_15 XI11_2/XI0/XI0_36/d__15_ xsel_36_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN1_14 XI11_2/XI0/XI0_36/d__14_ xsel_36_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN1_13 XI11_2/XI0/XI0_36/d__13_ xsel_36_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN1_12 XI11_2/XI0/XI0_36/d__12_ xsel_36_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN1_11 XI11_2/XI0/XI0_36/d__11_ xsel_36_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN1_10 XI11_2/XI0/XI0_36/d__10_ xsel_36_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN1_9 XI11_2/XI0/XI0_36/d__9_ xsel_36_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN1_8 XI11_2/XI0/XI0_36/d__8_ xsel_36_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN1_7 XI11_2/XI0/XI0_36/d__7_ xsel_36_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN1_6 XI11_2/XI0/XI0_36/d__6_ xsel_36_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN1_5 XI11_2/XI0/XI0_36/d__5_ xsel_36_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN1_4 XI11_2/XI0/XI0_36/d__4_ xsel_36_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN1_3 XI11_2/XI0/XI0_36/d__3_ xsel_36_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN1_2 XI11_2/XI0/XI0_36/d__2_ xsel_36_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN1_1 XI11_2/XI0/XI0_36/d__1_ xsel_36_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_36/MN1_0 XI11_2/XI0/XI0_36/d__0_ xsel_36_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN0_15 XI11_2/net21_0_ xsel_35_ XI11_2/XI0/XI0_35/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN0_14 XI11_2/net21_1_ xsel_35_ XI11_2/XI0/XI0_35/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN0_13 XI11_2/net21_2_ xsel_35_ XI11_2/XI0/XI0_35/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN0_12 XI11_2/net21_3_ xsel_35_ XI11_2/XI0/XI0_35/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN0_11 XI11_2/net21_4_ xsel_35_ XI11_2/XI0/XI0_35/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN0_10 XI11_2/net21_5_ xsel_35_ XI11_2/XI0/XI0_35/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN0_9 XI11_2/net21_6_ xsel_35_ XI11_2/XI0/XI0_35/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN0_8 XI11_2/net21_7_ xsel_35_ XI11_2/XI0/XI0_35/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN0_7 XI11_2/net21_8_ xsel_35_ XI11_2/XI0/XI0_35/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN0_6 XI11_2/net21_9_ xsel_35_ XI11_2/XI0/XI0_35/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN0_5 XI11_2/net21_10_ xsel_35_ XI11_2/XI0/XI0_35/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN0_4 XI11_2/net21_11_ xsel_35_ XI11_2/XI0/XI0_35/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN0_3 XI11_2/net21_12_ xsel_35_ XI11_2/XI0/XI0_35/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN0_2 XI11_2/net21_13_ xsel_35_ XI11_2/XI0/XI0_35/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN0_1 XI11_2/net21_14_ xsel_35_ XI11_2/XI0/XI0_35/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN0_0 XI11_2/net21_15_ xsel_35_ XI11_2/XI0/XI0_35/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN1_15 XI11_2/XI0/XI0_35/d__15_ xsel_35_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN1_14 XI11_2/XI0/XI0_35/d__14_ xsel_35_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN1_13 XI11_2/XI0/XI0_35/d__13_ xsel_35_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN1_12 XI11_2/XI0/XI0_35/d__12_ xsel_35_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN1_11 XI11_2/XI0/XI0_35/d__11_ xsel_35_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN1_10 XI11_2/XI0/XI0_35/d__10_ xsel_35_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN1_9 XI11_2/XI0/XI0_35/d__9_ xsel_35_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN1_8 XI11_2/XI0/XI0_35/d__8_ xsel_35_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN1_7 XI11_2/XI0/XI0_35/d__7_ xsel_35_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN1_6 XI11_2/XI0/XI0_35/d__6_ xsel_35_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN1_5 XI11_2/XI0/XI0_35/d__5_ xsel_35_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN1_4 XI11_2/XI0/XI0_35/d__4_ xsel_35_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN1_3 XI11_2/XI0/XI0_35/d__3_ xsel_35_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN1_2 XI11_2/XI0/XI0_35/d__2_ xsel_35_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN1_1 XI11_2/XI0/XI0_35/d__1_ xsel_35_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_35/MN1_0 XI11_2/XI0/XI0_35/d__0_ xsel_35_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN0_15 XI11_2/net21_0_ xsel_34_ XI11_2/XI0/XI0_34/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN0_14 XI11_2/net21_1_ xsel_34_ XI11_2/XI0/XI0_34/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN0_13 XI11_2/net21_2_ xsel_34_ XI11_2/XI0/XI0_34/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN0_12 XI11_2/net21_3_ xsel_34_ XI11_2/XI0/XI0_34/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN0_11 XI11_2/net21_4_ xsel_34_ XI11_2/XI0/XI0_34/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN0_10 XI11_2/net21_5_ xsel_34_ XI11_2/XI0/XI0_34/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN0_9 XI11_2/net21_6_ xsel_34_ XI11_2/XI0/XI0_34/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN0_8 XI11_2/net21_7_ xsel_34_ XI11_2/XI0/XI0_34/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN0_7 XI11_2/net21_8_ xsel_34_ XI11_2/XI0/XI0_34/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN0_6 XI11_2/net21_9_ xsel_34_ XI11_2/XI0/XI0_34/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN0_5 XI11_2/net21_10_ xsel_34_ XI11_2/XI0/XI0_34/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN0_4 XI11_2/net21_11_ xsel_34_ XI11_2/XI0/XI0_34/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN0_3 XI11_2/net21_12_ xsel_34_ XI11_2/XI0/XI0_34/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN0_2 XI11_2/net21_13_ xsel_34_ XI11_2/XI0/XI0_34/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN0_1 XI11_2/net21_14_ xsel_34_ XI11_2/XI0/XI0_34/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN0_0 XI11_2/net21_15_ xsel_34_ XI11_2/XI0/XI0_34/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN1_15 XI11_2/XI0/XI0_34/d__15_ xsel_34_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN1_14 XI11_2/XI0/XI0_34/d__14_ xsel_34_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN1_13 XI11_2/XI0/XI0_34/d__13_ xsel_34_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN1_12 XI11_2/XI0/XI0_34/d__12_ xsel_34_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN1_11 XI11_2/XI0/XI0_34/d__11_ xsel_34_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN1_10 XI11_2/XI0/XI0_34/d__10_ xsel_34_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN1_9 XI11_2/XI0/XI0_34/d__9_ xsel_34_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN1_8 XI11_2/XI0/XI0_34/d__8_ xsel_34_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN1_7 XI11_2/XI0/XI0_34/d__7_ xsel_34_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN1_6 XI11_2/XI0/XI0_34/d__6_ xsel_34_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN1_5 XI11_2/XI0/XI0_34/d__5_ xsel_34_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN1_4 XI11_2/XI0/XI0_34/d__4_ xsel_34_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN1_3 XI11_2/XI0/XI0_34/d__3_ xsel_34_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN1_2 XI11_2/XI0/XI0_34/d__2_ xsel_34_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN1_1 XI11_2/XI0/XI0_34/d__1_ xsel_34_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_34/MN1_0 XI11_2/XI0/XI0_34/d__0_ xsel_34_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN0_15 XI11_2/net21_0_ xsel_33_ XI11_2/XI0/XI0_33/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN0_14 XI11_2/net21_1_ xsel_33_ XI11_2/XI0/XI0_33/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN0_13 XI11_2/net21_2_ xsel_33_ XI11_2/XI0/XI0_33/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN0_12 XI11_2/net21_3_ xsel_33_ XI11_2/XI0/XI0_33/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN0_11 XI11_2/net21_4_ xsel_33_ XI11_2/XI0/XI0_33/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN0_10 XI11_2/net21_5_ xsel_33_ XI11_2/XI0/XI0_33/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN0_9 XI11_2/net21_6_ xsel_33_ XI11_2/XI0/XI0_33/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN0_8 XI11_2/net21_7_ xsel_33_ XI11_2/XI0/XI0_33/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN0_7 XI11_2/net21_8_ xsel_33_ XI11_2/XI0/XI0_33/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN0_6 XI11_2/net21_9_ xsel_33_ XI11_2/XI0/XI0_33/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN0_5 XI11_2/net21_10_ xsel_33_ XI11_2/XI0/XI0_33/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN0_4 XI11_2/net21_11_ xsel_33_ XI11_2/XI0/XI0_33/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN0_3 XI11_2/net21_12_ xsel_33_ XI11_2/XI0/XI0_33/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN0_2 XI11_2/net21_13_ xsel_33_ XI11_2/XI0/XI0_33/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN0_1 XI11_2/net21_14_ xsel_33_ XI11_2/XI0/XI0_33/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN0_0 XI11_2/net21_15_ xsel_33_ XI11_2/XI0/XI0_33/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN1_15 XI11_2/XI0/XI0_33/d__15_ xsel_33_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN1_14 XI11_2/XI0/XI0_33/d__14_ xsel_33_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN1_13 XI11_2/XI0/XI0_33/d__13_ xsel_33_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN1_12 XI11_2/XI0/XI0_33/d__12_ xsel_33_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN1_11 XI11_2/XI0/XI0_33/d__11_ xsel_33_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN1_10 XI11_2/XI0/XI0_33/d__10_ xsel_33_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN1_9 XI11_2/XI0/XI0_33/d__9_ xsel_33_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN1_8 XI11_2/XI0/XI0_33/d__8_ xsel_33_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN1_7 XI11_2/XI0/XI0_33/d__7_ xsel_33_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN1_6 XI11_2/XI0/XI0_33/d__6_ xsel_33_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN1_5 XI11_2/XI0/XI0_33/d__5_ xsel_33_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN1_4 XI11_2/XI0/XI0_33/d__4_ xsel_33_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN1_3 XI11_2/XI0/XI0_33/d__3_ xsel_33_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN1_2 XI11_2/XI0/XI0_33/d__2_ xsel_33_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN1_1 XI11_2/XI0/XI0_33/d__1_ xsel_33_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_33/MN1_0 XI11_2/XI0/XI0_33/d__0_ xsel_33_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN0_15 XI11_2/net21_0_ xsel_32_ XI11_2/XI0/XI0_32/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN0_14 XI11_2/net21_1_ xsel_32_ XI11_2/XI0/XI0_32/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN0_13 XI11_2/net21_2_ xsel_32_ XI11_2/XI0/XI0_32/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN0_12 XI11_2/net21_3_ xsel_32_ XI11_2/XI0/XI0_32/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN0_11 XI11_2/net21_4_ xsel_32_ XI11_2/XI0/XI0_32/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN0_10 XI11_2/net21_5_ xsel_32_ XI11_2/XI0/XI0_32/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN0_9 XI11_2/net21_6_ xsel_32_ XI11_2/XI0/XI0_32/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN0_8 XI11_2/net21_7_ xsel_32_ XI11_2/XI0/XI0_32/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN0_7 XI11_2/net21_8_ xsel_32_ XI11_2/XI0/XI0_32/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN0_6 XI11_2/net21_9_ xsel_32_ XI11_2/XI0/XI0_32/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN0_5 XI11_2/net21_10_ xsel_32_ XI11_2/XI0/XI0_32/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN0_4 XI11_2/net21_11_ xsel_32_ XI11_2/XI0/XI0_32/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN0_3 XI11_2/net21_12_ xsel_32_ XI11_2/XI0/XI0_32/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN0_2 XI11_2/net21_13_ xsel_32_ XI11_2/XI0/XI0_32/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN0_1 XI11_2/net21_14_ xsel_32_ XI11_2/XI0/XI0_32/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN0_0 XI11_2/net21_15_ xsel_32_ XI11_2/XI0/XI0_32/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN1_15 XI11_2/XI0/XI0_32/d__15_ xsel_32_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN1_14 XI11_2/XI0/XI0_32/d__14_ xsel_32_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN1_13 XI11_2/XI0/XI0_32/d__13_ xsel_32_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN1_12 XI11_2/XI0/XI0_32/d__12_ xsel_32_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN1_11 XI11_2/XI0/XI0_32/d__11_ xsel_32_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN1_10 XI11_2/XI0/XI0_32/d__10_ xsel_32_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN1_9 XI11_2/XI0/XI0_32/d__9_ xsel_32_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN1_8 XI11_2/XI0/XI0_32/d__8_ xsel_32_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN1_7 XI11_2/XI0/XI0_32/d__7_ xsel_32_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN1_6 XI11_2/XI0/XI0_32/d__6_ xsel_32_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN1_5 XI11_2/XI0/XI0_32/d__5_ xsel_32_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN1_4 XI11_2/XI0/XI0_32/d__4_ xsel_32_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN1_3 XI11_2/XI0/XI0_32/d__3_ xsel_32_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN1_2 XI11_2/XI0/XI0_32/d__2_ xsel_32_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN1_1 XI11_2/XI0/XI0_32/d__1_ xsel_32_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_32/MN1_0 XI11_2/XI0/XI0_32/d__0_ xsel_32_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN0_15 XI11_2/net21_0_ xsel_31_ XI11_2/XI0/XI0_31/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN0_14 XI11_2/net21_1_ xsel_31_ XI11_2/XI0/XI0_31/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN0_13 XI11_2/net21_2_ xsel_31_ XI11_2/XI0/XI0_31/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN0_12 XI11_2/net21_3_ xsel_31_ XI11_2/XI0/XI0_31/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN0_11 XI11_2/net21_4_ xsel_31_ XI11_2/XI0/XI0_31/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN0_10 XI11_2/net21_5_ xsel_31_ XI11_2/XI0/XI0_31/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN0_9 XI11_2/net21_6_ xsel_31_ XI11_2/XI0/XI0_31/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN0_8 XI11_2/net21_7_ xsel_31_ XI11_2/XI0/XI0_31/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN0_7 XI11_2/net21_8_ xsel_31_ XI11_2/XI0/XI0_31/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN0_6 XI11_2/net21_9_ xsel_31_ XI11_2/XI0/XI0_31/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN0_5 XI11_2/net21_10_ xsel_31_ XI11_2/XI0/XI0_31/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN0_4 XI11_2/net21_11_ xsel_31_ XI11_2/XI0/XI0_31/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN0_3 XI11_2/net21_12_ xsel_31_ XI11_2/XI0/XI0_31/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN0_2 XI11_2/net21_13_ xsel_31_ XI11_2/XI0/XI0_31/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN0_1 XI11_2/net21_14_ xsel_31_ XI11_2/XI0/XI0_31/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN0_0 XI11_2/net21_15_ xsel_31_ XI11_2/XI0/XI0_31/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN1_15 XI11_2/XI0/XI0_31/d__15_ xsel_31_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN1_14 XI11_2/XI0/XI0_31/d__14_ xsel_31_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN1_13 XI11_2/XI0/XI0_31/d__13_ xsel_31_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN1_12 XI11_2/XI0/XI0_31/d__12_ xsel_31_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN1_11 XI11_2/XI0/XI0_31/d__11_ xsel_31_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN1_10 XI11_2/XI0/XI0_31/d__10_ xsel_31_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN1_9 XI11_2/XI0/XI0_31/d__9_ xsel_31_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN1_8 XI11_2/XI0/XI0_31/d__8_ xsel_31_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN1_7 XI11_2/XI0/XI0_31/d__7_ xsel_31_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN1_6 XI11_2/XI0/XI0_31/d__6_ xsel_31_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN1_5 XI11_2/XI0/XI0_31/d__5_ xsel_31_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN1_4 XI11_2/XI0/XI0_31/d__4_ xsel_31_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN1_3 XI11_2/XI0/XI0_31/d__3_ xsel_31_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN1_2 XI11_2/XI0/XI0_31/d__2_ xsel_31_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN1_1 XI11_2/XI0/XI0_31/d__1_ xsel_31_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_31/MN1_0 XI11_2/XI0/XI0_31/d__0_ xsel_31_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN0_15 XI11_2/net21_0_ xsel_30_ XI11_2/XI0/XI0_30/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN0_14 XI11_2/net21_1_ xsel_30_ XI11_2/XI0/XI0_30/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN0_13 XI11_2/net21_2_ xsel_30_ XI11_2/XI0/XI0_30/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN0_12 XI11_2/net21_3_ xsel_30_ XI11_2/XI0/XI0_30/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN0_11 XI11_2/net21_4_ xsel_30_ XI11_2/XI0/XI0_30/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN0_10 XI11_2/net21_5_ xsel_30_ XI11_2/XI0/XI0_30/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN0_9 XI11_2/net21_6_ xsel_30_ XI11_2/XI0/XI0_30/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN0_8 XI11_2/net21_7_ xsel_30_ XI11_2/XI0/XI0_30/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN0_7 XI11_2/net21_8_ xsel_30_ XI11_2/XI0/XI0_30/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN0_6 XI11_2/net21_9_ xsel_30_ XI11_2/XI0/XI0_30/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN0_5 XI11_2/net21_10_ xsel_30_ XI11_2/XI0/XI0_30/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN0_4 XI11_2/net21_11_ xsel_30_ XI11_2/XI0/XI0_30/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN0_3 XI11_2/net21_12_ xsel_30_ XI11_2/XI0/XI0_30/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN0_2 XI11_2/net21_13_ xsel_30_ XI11_2/XI0/XI0_30/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN0_1 XI11_2/net21_14_ xsel_30_ XI11_2/XI0/XI0_30/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN0_0 XI11_2/net21_15_ xsel_30_ XI11_2/XI0/XI0_30/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN1_15 XI11_2/XI0/XI0_30/d__15_ xsel_30_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN1_14 XI11_2/XI0/XI0_30/d__14_ xsel_30_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN1_13 XI11_2/XI0/XI0_30/d__13_ xsel_30_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN1_12 XI11_2/XI0/XI0_30/d__12_ xsel_30_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN1_11 XI11_2/XI0/XI0_30/d__11_ xsel_30_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN1_10 XI11_2/XI0/XI0_30/d__10_ xsel_30_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN1_9 XI11_2/XI0/XI0_30/d__9_ xsel_30_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN1_8 XI11_2/XI0/XI0_30/d__8_ xsel_30_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN1_7 XI11_2/XI0/XI0_30/d__7_ xsel_30_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN1_6 XI11_2/XI0/XI0_30/d__6_ xsel_30_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN1_5 XI11_2/XI0/XI0_30/d__5_ xsel_30_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN1_4 XI11_2/XI0/XI0_30/d__4_ xsel_30_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN1_3 XI11_2/XI0/XI0_30/d__3_ xsel_30_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN1_2 XI11_2/XI0/XI0_30/d__2_ xsel_30_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN1_1 XI11_2/XI0/XI0_30/d__1_ xsel_30_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_30/MN1_0 XI11_2/XI0/XI0_30/d__0_ xsel_30_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN0_15 XI11_2/net21_0_ xsel_29_ XI11_2/XI0/XI0_29/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN0_14 XI11_2/net21_1_ xsel_29_ XI11_2/XI0/XI0_29/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN0_13 XI11_2/net21_2_ xsel_29_ XI11_2/XI0/XI0_29/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN0_12 XI11_2/net21_3_ xsel_29_ XI11_2/XI0/XI0_29/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN0_11 XI11_2/net21_4_ xsel_29_ XI11_2/XI0/XI0_29/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN0_10 XI11_2/net21_5_ xsel_29_ XI11_2/XI0/XI0_29/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN0_9 XI11_2/net21_6_ xsel_29_ XI11_2/XI0/XI0_29/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN0_8 XI11_2/net21_7_ xsel_29_ XI11_2/XI0/XI0_29/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN0_7 XI11_2/net21_8_ xsel_29_ XI11_2/XI0/XI0_29/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN0_6 XI11_2/net21_9_ xsel_29_ XI11_2/XI0/XI0_29/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN0_5 XI11_2/net21_10_ xsel_29_ XI11_2/XI0/XI0_29/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN0_4 XI11_2/net21_11_ xsel_29_ XI11_2/XI0/XI0_29/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN0_3 XI11_2/net21_12_ xsel_29_ XI11_2/XI0/XI0_29/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN0_2 XI11_2/net21_13_ xsel_29_ XI11_2/XI0/XI0_29/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN0_1 XI11_2/net21_14_ xsel_29_ XI11_2/XI0/XI0_29/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN0_0 XI11_2/net21_15_ xsel_29_ XI11_2/XI0/XI0_29/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN1_15 XI11_2/XI0/XI0_29/d__15_ xsel_29_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN1_14 XI11_2/XI0/XI0_29/d__14_ xsel_29_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN1_13 XI11_2/XI0/XI0_29/d__13_ xsel_29_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN1_12 XI11_2/XI0/XI0_29/d__12_ xsel_29_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN1_11 XI11_2/XI0/XI0_29/d__11_ xsel_29_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN1_10 XI11_2/XI0/XI0_29/d__10_ xsel_29_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN1_9 XI11_2/XI0/XI0_29/d__9_ xsel_29_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN1_8 XI11_2/XI0/XI0_29/d__8_ xsel_29_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN1_7 XI11_2/XI0/XI0_29/d__7_ xsel_29_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN1_6 XI11_2/XI0/XI0_29/d__6_ xsel_29_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN1_5 XI11_2/XI0/XI0_29/d__5_ xsel_29_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN1_4 XI11_2/XI0/XI0_29/d__4_ xsel_29_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN1_3 XI11_2/XI0/XI0_29/d__3_ xsel_29_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN1_2 XI11_2/XI0/XI0_29/d__2_ xsel_29_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN1_1 XI11_2/XI0/XI0_29/d__1_ xsel_29_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_29/MN1_0 XI11_2/XI0/XI0_29/d__0_ xsel_29_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN0_15 XI11_2/net21_0_ xsel_28_ XI11_2/XI0/XI0_28/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN0_14 XI11_2/net21_1_ xsel_28_ XI11_2/XI0/XI0_28/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN0_13 XI11_2/net21_2_ xsel_28_ XI11_2/XI0/XI0_28/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN0_12 XI11_2/net21_3_ xsel_28_ XI11_2/XI0/XI0_28/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN0_11 XI11_2/net21_4_ xsel_28_ XI11_2/XI0/XI0_28/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN0_10 XI11_2/net21_5_ xsel_28_ XI11_2/XI0/XI0_28/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN0_9 XI11_2/net21_6_ xsel_28_ XI11_2/XI0/XI0_28/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN0_8 XI11_2/net21_7_ xsel_28_ XI11_2/XI0/XI0_28/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN0_7 XI11_2/net21_8_ xsel_28_ XI11_2/XI0/XI0_28/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN0_6 XI11_2/net21_9_ xsel_28_ XI11_2/XI0/XI0_28/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN0_5 XI11_2/net21_10_ xsel_28_ XI11_2/XI0/XI0_28/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN0_4 XI11_2/net21_11_ xsel_28_ XI11_2/XI0/XI0_28/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN0_3 XI11_2/net21_12_ xsel_28_ XI11_2/XI0/XI0_28/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN0_2 XI11_2/net21_13_ xsel_28_ XI11_2/XI0/XI0_28/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN0_1 XI11_2/net21_14_ xsel_28_ XI11_2/XI0/XI0_28/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN0_0 XI11_2/net21_15_ xsel_28_ XI11_2/XI0/XI0_28/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN1_15 XI11_2/XI0/XI0_28/d__15_ xsel_28_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN1_14 XI11_2/XI0/XI0_28/d__14_ xsel_28_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN1_13 XI11_2/XI0/XI0_28/d__13_ xsel_28_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN1_12 XI11_2/XI0/XI0_28/d__12_ xsel_28_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN1_11 XI11_2/XI0/XI0_28/d__11_ xsel_28_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN1_10 XI11_2/XI0/XI0_28/d__10_ xsel_28_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN1_9 XI11_2/XI0/XI0_28/d__9_ xsel_28_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN1_8 XI11_2/XI0/XI0_28/d__8_ xsel_28_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN1_7 XI11_2/XI0/XI0_28/d__7_ xsel_28_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN1_6 XI11_2/XI0/XI0_28/d__6_ xsel_28_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN1_5 XI11_2/XI0/XI0_28/d__5_ xsel_28_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN1_4 XI11_2/XI0/XI0_28/d__4_ xsel_28_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN1_3 XI11_2/XI0/XI0_28/d__3_ xsel_28_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN1_2 XI11_2/XI0/XI0_28/d__2_ xsel_28_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN1_1 XI11_2/XI0/XI0_28/d__1_ xsel_28_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_28/MN1_0 XI11_2/XI0/XI0_28/d__0_ xsel_28_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN0_15 XI11_2/net21_0_ xsel_27_ XI11_2/XI0/XI0_27/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN0_14 XI11_2/net21_1_ xsel_27_ XI11_2/XI0/XI0_27/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN0_13 XI11_2/net21_2_ xsel_27_ XI11_2/XI0/XI0_27/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN0_12 XI11_2/net21_3_ xsel_27_ XI11_2/XI0/XI0_27/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN0_11 XI11_2/net21_4_ xsel_27_ XI11_2/XI0/XI0_27/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN0_10 XI11_2/net21_5_ xsel_27_ XI11_2/XI0/XI0_27/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN0_9 XI11_2/net21_6_ xsel_27_ XI11_2/XI0/XI0_27/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN0_8 XI11_2/net21_7_ xsel_27_ XI11_2/XI0/XI0_27/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN0_7 XI11_2/net21_8_ xsel_27_ XI11_2/XI0/XI0_27/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN0_6 XI11_2/net21_9_ xsel_27_ XI11_2/XI0/XI0_27/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN0_5 XI11_2/net21_10_ xsel_27_ XI11_2/XI0/XI0_27/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN0_4 XI11_2/net21_11_ xsel_27_ XI11_2/XI0/XI0_27/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN0_3 XI11_2/net21_12_ xsel_27_ XI11_2/XI0/XI0_27/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN0_2 XI11_2/net21_13_ xsel_27_ XI11_2/XI0/XI0_27/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN0_1 XI11_2/net21_14_ xsel_27_ XI11_2/XI0/XI0_27/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN0_0 XI11_2/net21_15_ xsel_27_ XI11_2/XI0/XI0_27/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN1_15 XI11_2/XI0/XI0_27/d__15_ xsel_27_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN1_14 XI11_2/XI0/XI0_27/d__14_ xsel_27_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN1_13 XI11_2/XI0/XI0_27/d__13_ xsel_27_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN1_12 XI11_2/XI0/XI0_27/d__12_ xsel_27_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN1_11 XI11_2/XI0/XI0_27/d__11_ xsel_27_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN1_10 XI11_2/XI0/XI0_27/d__10_ xsel_27_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN1_9 XI11_2/XI0/XI0_27/d__9_ xsel_27_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN1_8 XI11_2/XI0/XI0_27/d__8_ xsel_27_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN1_7 XI11_2/XI0/XI0_27/d__7_ xsel_27_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN1_6 XI11_2/XI0/XI0_27/d__6_ xsel_27_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN1_5 XI11_2/XI0/XI0_27/d__5_ xsel_27_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN1_4 XI11_2/XI0/XI0_27/d__4_ xsel_27_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN1_3 XI11_2/XI0/XI0_27/d__3_ xsel_27_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN1_2 XI11_2/XI0/XI0_27/d__2_ xsel_27_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN1_1 XI11_2/XI0/XI0_27/d__1_ xsel_27_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_27/MN1_0 XI11_2/XI0/XI0_27/d__0_ xsel_27_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN0_15 XI11_2/net21_0_ xsel_26_ XI11_2/XI0/XI0_26/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN0_14 XI11_2/net21_1_ xsel_26_ XI11_2/XI0/XI0_26/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN0_13 XI11_2/net21_2_ xsel_26_ XI11_2/XI0/XI0_26/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN0_12 XI11_2/net21_3_ xsel_26_ XI11_2/XI0/XI0_26/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN0_11 XI11_2/net21_4_ xsel_26_ XI11_2/XI0/XI0_26/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN0_10 XI11_2/net21_5_ xsel_26_ XI11_2/XI0/XI0_26/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN0_9 XI11_2/net21_6_ xsel_26_ XI11_2/XI0/XI0_26/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN0_8 XI11_2/net21_7_ xsel_26_ XI11_2/XI0/XI0_26/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN0_7 XI11_2/net21_8_ xsel_26_ XI11_2/XI0/XI0_26/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN0_6 XI11_2/net21_9_ xsel_26_ XI11_2/XI0/XI0_26/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN0_5 XI11_2/net21_10_ xsel_26_ XI11_2/XI0/XI0_26/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN0_4 XI11_2/net21_11_ xsel_26_ XI11_2/XI0/XI0_26/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN0_3 XI11_2/net21_12_ xsel_26_ XI11_2/XI0/XI0_26/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN0_2 XI11_2/net21_13_ xsel_26_ XI11_2/XI0/XI0_26/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN0_1 XI11_2/net21_14_ xsel_26_ XI11_2/XI0/XI0_26/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN0_0 XI11_2/net21_15_ xsel_26_ XI11_2/XI0/XI0_26/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN1_15 XI11_2/XI0/XI0_26/d__15_ xsel_26_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN1_14 XI11_2/XI0/XI0_26/d__14_ xsel_26_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN1_13 XI11_2/XI0/XI0_26/d__13_ xsel_26_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN1_12 XI11_2/XI0/XI0_26/d__12_ xsel_26_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN1_11 XI11_2/XI0/XI0_26/d__11_ xsel_26_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN1_10 XI11_2/XI0/XI0_26/d__10_ xsel_26_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN1_9 XI11_2/XI0/XI0_26/d__9_ xsel_26_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN1_8 XI11_2/XI0/XI0_26/d__8_ xsel_26_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN1_7 XI11_2/XI0/XI0_26/d__7_ xsel_26_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN1_6 XI11_2/XI0/XI0_26/d__6_ xsel_26_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN1_5 XI11_2/XI0/XI0_26/d__5_ xsel_26_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN1_4 XI11_2/XI0/XI0_26/d__4_ xsel_26_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN1_3 XI11_2/XI0/XI0_26/d__3_ xsel_26_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN1_2 XI11_2/XI0/XI0_26/d__2_ xsel_26_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN1_1 XI11_2/XI0/XI0_26/d__1_ xsel_26_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_26/MN1_0 XI11_2/XI0/XI0_26/d__0_ xsel_26_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN0_15 XI11_2/net21_0_ xsel_25_ XI11_2/XI0/XI0_25/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN0_14 XI11_2/net21_1_ xsel_25_ XI11_2/XI0/XI0_25/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN0_13 XI11_2/net21_2_ xsel_25_ XI11_2/XI0/XI0_25/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN0_12 XI11_2/net21_3_ xsel_25_ XI11_2/XI0/XI0_25/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN0_11 XI11_2/net21_4_ xsel_25_ XI11_2/XI0/XI0_25/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN0_10 XI11_2/net21_5_ xsel_25_ XI11_2/XI0/XI0_25/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN0_9 XI11_2/net21_6_ xsel_25_ XI11_2/XI0/XI0_25/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN0_8 XI11_2/net21_7_ xsel_25_ XI11_2/XI0/XI0_25/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN0_7 XI11_2/net21_8_ xsel_25_ XI11_2/XI0/XI0_25/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN0_6 XI11_2/net21_9_ xsel_25_ XI11_2/XI0/XI0_25/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN0_5 XI11_2/net21_10_ xsel_25_ XI11_2/XI0/XI0_25/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN0_4 XI11_2/net21_11_ xsel_25_ XI11_2/XI0/XI0_25/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN0_3 XI11_2/net21_12_ xsel_25_ XI11_2/XI0/XI0_25/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN0_2 XI11_2/net21_13_ xsel_25_ XI11_2/XI0/XI0_25/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN0_1 XI11_2/net21_14_ xsel_25_ XI11_2/XI0/XI0_25/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN0_0 XI11_2/net21_15_ xsel_25_ XI11_2/XI0/XI0_25/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN1_15 XI11_2/XI0/XI0_25/d__15_ xsel_25_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN1_14 XI11_2/XI0/XI0_25/d__14_ xsel_25_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN1_13 XI11_2/XI0/XI0_25/d__13_ xsel_25_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN1_12 XI11_2/XI0/XI0_25/d__12_ xsel_25_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN1_11 XI11_2/XI0/XI0_25/d__11_ xsel_25_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN1_10 XI11_2/XI0/XI0_25/d__10_ xsel_25_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN1_9 XI11_2/XI0/XI0_25/d__9_ xsel_25_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN1_8 XI11_2/XI0/XI0_25/d__8_ xsel_25_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN1_7 XI11_2/XI0/XI0_25/d__7_ xsel_25_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN1_6 XI11_2/XI0/XI0_25/d__6_ xsel_25_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN1_5 XI11_2/XI0/XI0_25/d__5_ xsel_25_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN1_4 XI11_2/XI0/XI0_25/d__4_ xsel_25_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN1_3 XI11_2/XI0/XI0_25/d__3_ xsel_25_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN1_2 XI11_2/XI0/XI0_25/d__2_ xsel_25_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN1_1 XI11_2/XI0/XI0_25/d__1_ xsel_25_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_25/MN1_0 XI11_2/XI0/XI0_25/d__0_ xsel_25_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN0_15 XI11_2/net21_0_ xsel_24_ XI11_2/XI0/XI0_24/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN0_14 XI11_2/net21_1_ xsel_24_ XI11_2/XI0/XI0_24/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN0_13 XI11_2/net21_2_ xsel_24_ XI11_2/XI0/XI0_24/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN0_12 XI11_2/net21_3_ xsel_24_ XI11_2/XI0/XI0_24/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN0_11 XI11_2/net21_4_ xsel_24_ XI11_2/XI0/XI0_24/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN0_10 XI11_2/net21_5_ xsel_24_ XI11_2/XI0/XI0_24/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN0_9 XI11_2/net21_6_ xsel_24_ XI11_2/XI0/XI0_24/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN0_8 XI11_2/net21_7_ xsel_24_ XI11_2/XI0/XI0_24/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN0_7 XI11_2/net21_8_ xsel_24_ XI11_2/XI0/XI0_24/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN0_6 XI11_2/net21_9_ xsel_24_ XI11_2/XI0/XI0_24/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN0_5 XI11_2/net21_10_ xsel_24_ XI11_2/XI0/XI0_24/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN0_4 XI11_2/net21_11_ xsel_24_ XI11_2/XI0/XI0_24/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN0_3 XI11_2/net21_12_ xsel_24_ XI11_2/XI0/XI0_24/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN0_2 XI11_2/net21_13_ xsel_24_ XI11_2/XI0/XI0_24/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN0_1 XI11_2/net21_14_ xsel_24_ XI11_2/XI0/XI0_24/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN0_0 XI11_2/net21_15_ xsel_24_ XI11_2/XI0/XI0_24/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN1_15 XI11_2/XI0/XI0_24/d__15_ xsel_24_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN1_14 XI11_2/XI0/XI0_24/d__14_ xsel_24_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN1_13 XI11_2/XI0/XI0_24/d__13_ xsel_24_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN1_12 XI11_2/XI0/XI0_24/d__12_ xsel_24_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN1_11 XI11_2/XI0/XI0_24/d__11_ xsel_24_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN1_10 XI11_2/XI0/XI0_24/d__10_ xsel_24_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN1_9 XI11_2/XI0/XI0_24/d__9_ xsel_24_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN1_8 XI11_2/XI0/XI0_24/d__8_ xsel_24_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN1_7 XI11_2/XI0/XI0_24/d__7_ xsel_24_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN1_6 XI11_2/XI0/XI0_24/d__6_ xsel_24_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN1_5 XI11_2/XI0/XI0_24/d__5_ xsel_24_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN1_4 XI11_2/XI0/XI0_24/d__4_ xsel_24_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN1_3 XI11_2/XI0/XI0_24/d__3_ xsel_24_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN1_2 XI11_2/XI0/XI0_24/d__2_ xsel_24_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN1_1 XI11_2/XI0/XI0_24/d__1_ xsel_24_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_24/MN1_0 XI11_2/XI0/XI0_24/d__0_ xsel_24_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN0_15 XI11_2/net21_0_ xsel_23_ XI11_2/XI0/XI0_23/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN0_14 XI11_2/net21_1_ xsel_23_ XI11_2/XI0/XI0_23/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN0_13 XI11_2/net21_2_ xsel_23_ XI11_2/XI0/XI0_23/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN0_12 XI11_2/net21_3_ xsel_23_ XI11_2/XI0/XI0_23/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN0_11 XI11_2/net21_4_ xsel_23_ XI11_2/XI0/XI0_23/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN0_10 XI11_2/net21_5_ xsel_23_ XI11_2/XI0/XI0_23/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN0_9 XI11_2/net21_6_ xsel_23_ XI11_2/XI0/XI0_23/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN0_8 XI11_2/net21_7_ xsel_23_ XI11_2/XI0/XI0_23/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN0_7 XI11_2/net21_8_ xsel_23_ XI11_2/XI0/XI0_23/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN0_6 XI11_2/net21_9_ xsel_23_ XI11_2/XI0/XI0_23/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN0_5 XI11_2/net21_10_ xsel_23_ XI11_2/XI0/XI0_23/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN0_4 XI11_2/net21_11_ xsel_23_ XI11_2/XI0/XI0_23/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN0_3 XI11_2/net21_12_ xsel_23_ XI11_2/XI0/XI0_23/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN0_2 XI11_2/net21_13_ xsel_23_ XI11_2/XI0/XI0_23/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN0_1 XI11_2/net21_14_ xsel_23_ XI11_2/XI0/XI0_23/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN0_0 XI11_2/net21_15_ xsel_23_ XI11_2/XI0/XI0_23/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN1_15 XI11_2/XI0/XI0_23/d__15_ xsel_23_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN1_14 XI11_2/XI0/XI0_23/d__14_ xsel_23_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN1_13 XI11_2/XI0/XI0_23/d__13_ xsel_23_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN1_12 XI11_2/XI0/XI0_23/d__12_ xsel_23_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN1_11 XI11_2/XI0/XI0_23/d__11_ xsel_23_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN1_10 XI11_2/XI0/XI0_23/d__10_ xsel_23_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN1_9 XI11_2/XI0/XI0_23/d__9_ xsel_23_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN1_8 XI11_2/XI0/XI0_23/d__8_ xsel_23_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN1_7 XI11_2/XI0/XI0_23/d__7_ xsel_23_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN1_6 XI11_2/XI0/XI0_23/d__6_ xsel_23_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN1_5 XI11_2/XI0/XI0_23/d__5_ xsel_23_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN1_4 XI11_2/XI0/XI0_23/d__4_ xsel_23_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN1_3 XI11_2/XI0/XI0_23/d__3_ xsel_23_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN1_2 XI11_2/XI0/XI0_23/d__2_ xsel_23_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN1_1 XI11_2/XI0/XI0_23/d__1_ xsel_23_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_23/MN1_0 XI11_2/XI0/XI0_23/d__0_ xsel_23_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN0_15 XI11_2/net21_0_ xsel_22_ XI11_2/XI0/XI0_22/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN0_14 XI11_2/net21_1_ xsel_22_ XI11_2/XI0/XI0_22/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN0_13 XI11_2/net21_2_ xsel_22_ XI11_2/XI0/XI0_22/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN0_12 XI11_2/net21_3_ xsel_22_ XI11_2/XI0/XI0_22/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN0_11 XI11_2/net21_4_ xsel_22_ XI11_2/XI0/XI0_22/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN0_10 XI11_2/net21_5_ xsel_22_ XI11_2/XI0/XI0_22/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN0_9 XI11_2/net21_6_ xsel_22_ XI11_2/XI0/XI0_22/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN0_8 XI11_2/net21_7_ xsel_22_ XI11_2/XI0/XI0_22/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN0_7 XI11_2/net21_8_ xsel_22_ XI11_2/XI0/XI0_22/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN0_6 XI11_2/net21_9_ xsel_22_ XI11_2/XI0/XI0_22/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN0_5 XI11_2/net21_10_ xsel_22_ XI11_2/XI0/XI0_22/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN0_4 XI11_2/net21_11_ xsel_22_ XI11_2/XI0/XI0_22/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN0_3 XI11_2/net21_12_ xsel_22_ XI11_2/XI0/XI0_22/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN0_2 XI11_2/net21_13_ xsel_22_ XI11_2/XI0/XI0_22/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN0_1 XI11_2/net21_14_ xsel_22_ XI11_2/XI0/XI0_22/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN0_0 XI11_2/net21_15_ xsel_22_ XI11_2/XI0/XI0_22/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN1_15 XI11_2/XI0/XI0_22/d__15_ xsel_22_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN1_14 XI11_2/XI0/XI0_22/d__14_ xsel_22_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN1_13 XI11_2/XI0/XI0_22/d__13_ xsel_22_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN1_12 XI11_2/XI0/XI0_22/d__12_ xsel_22_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN1_11 XI11_2/XI0/XI0_22/d__11_ xsel_22_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN1_10 XI11_2/XI0/XI0_22/d__10_ xsel_22_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN1_9 XI11_2/XI0/XI0_22/d__9_ xsel_22_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN1_8 XI11_2/XI0/XI0_22/d__8_ xsel_22_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN1_7 XI11_2/XI0/XI0_22/d__7_ xsel_22_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN1_6 XI11_2/XI0/XI0_22/d__6_ xsel_22_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN1_5 XI11_2/XI0/XI0_22/d__5_ xsel_22_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN1_4 XI11_2/XI0/XI0_22/d__4_ xsel_22_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN1_3 XI11_2/XI0/XI0_22/d__3_ xsel_22_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN1_2 XI11_2/XI0/XI0_22/d__2_ xsel_22_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN1_1 XI11_2/XI0/XI0_22/d__1_ xsel_22_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_22/MN1_0 XI11_2/XI0/XI0_22/d__0_ xsel_22_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN0_15 XI11_2/net21_0_ xsel_21_ XI11_2/XI0/XI0_21/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN0_14 XI11_2/net21_1_ xsel_21_ XI11_2/XI0/XI0_21/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN0_13 XI11_2/net21_2_ xsel_21_ XI11_2/XI0/XI0_21/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN0_12 XI11_2/net21_3_ xsel_21_ XI11_2/XI0/XI0_21/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN0_11 XI11_2/net21_4_ xsel_21_ XI11_2/XI0/XI0_21/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN0_10 XI11_2/net21_5_ xsel_21_ XI11_2/XI0/XI0_21/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN0_9 XI11_2/net21_6_ xsel_21_ XI11_2/XI0/XI0_21/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN0_8 XI11_2/net21_7_ xsel_21_ XI11_2/XI0/XI0_21/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN0_7 XI11_2/net21_8_ xsel_21_ XI11_2/XI0/XI0_21/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN0_6 XI11_2/net21_9_ xsel_21_ XI11_2/XI0/XI0_21/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN0_5 XI11_2/net21_10_ xsel_21_ XI11_2/XI0/XI0_21/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN0_4 XI11_2/net21_11_ xsel_21_ XI11_2/XI0/XI0_21/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN0_3 XI11_2/net21_12_ xsel_21_ XI11_2/XI0/XI0_21/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN0_2 XI11_2/net21_13_ xsel_21_ XI11_2/XI0/XI0_21/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN0_1 XI11_2/net21_14_ xsel_21_ XI11_2/XI0/XI0_21/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN0_0 XI11_2/net21_15_ xsel_21_ XI11_2/XI0/XI0_21/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN1_15 XI11_2/XI0/XI0_21/d__15_ xsel_21_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN1_14 XI11_2/XI0/XI0_21/d__14_ xsel_21_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN1_13 XI11_2/XI0/XI0_21/d__13_ xsel_21_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN1_12 XI11_2/XI0/XI0_21/d__12_ xsel_21_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN1_11 XI11_2/XI0/XI0_21/d__11_ xsel_21_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN1_10 XI11_2/XI0/XI0_21/d__10_ xsel_21_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN1_9 XI11_2/XI0/XI0_21/d__9_ xsel_21_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN1_8 XI11_2/XI0/XI0_21/d__8_ xsel_21_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN1_7 XI11_2/XI0/XI0_21/d__7_ xsel_21_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN1_6 XI11_2/XI0/XI0_21/d__6_ xsel_21_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN1_5 XI11_2/XI0/XI0_21/d__5_ xsel_21_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN1_4 XI11_2/XI0/XI0_21/d__4_ xsel_21_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN1_3 XI11_2/XI0/XI0_21/d__3_ xsel_21_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN1_2 XI11_2/XI0/XI0_21/d__2_ xsel_21_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN1_1 XI11_2/XI0/XI0_21/d__1_ xsel_21_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_21/MN1_0 XI11_2/XI0/XI0_21/d__0_ xsel_21_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN0_15 XI11_2/net21_0_ xsel_20_ XI11_2/XI0/XI0_20/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN0_14 XI11_2/net21_1_ xsel_20_ XI11_2/XI0/XI0_20/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN0_13 XI11_2/net21_2_ xsel_20_ XI11_2/XI0/XI0_20/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN0_12 XI11_2/net21_3_ xsel_20_ XI11_2/XI0/XI0_20/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN0_11 XI11_2/net21_4_ xsel_20_ XI11_2/XI0/XI0_20/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN0_10 XI11_2/net21_5_ xsel_20_ XI11_2/XI0/XI0_20/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN0_9 XI11_2/net21_6_ xsel_20_ XI11_2/XI0/XI0_20/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN0_8 XI11_2/net21_7_ xsel_20_ XI11_2/XI0/XI0_20/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN0_7 XI11_2/net21_8_ xsel_20_ XI11_2/XI0/XI0_20/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN0_6 XI11_2/net21_9_ xsel_20_ XI11_2/XI0/XI0_20/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN0_5 XI11_2/net21_10_ xsel_20_ XI11_2/XI0/XI0_20/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN0_4 XI11_2/net21_11_ xsel_20_ XI11_2/XI0/XI0_20/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN0_3 XI11_2/net21_12_ xsel_20_ XI11_2/XI0/XI0_20/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN0_2 XI11_2/net21_13_ xsel_20_ XI11_2/XI0/XI0_20/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN0_1 XI11_2/net21_14_ xsel_20_ XI11_2/XI0/XI0_20/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN0_0 XI11_2/net21_15_ xsel_20_ XI11_2/XI0/XI0_20/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN1_15 XI11_2/XI0/XI0_20/d__15_ xsel_20_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN1_14 XI11_2/XI0/XI0_20/d__14_ xsel_20_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN1_13 XI11_2/XI0/XI0_20/d__13_ xsel_20_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN1_12 XI11_2/XI0/XI0_20/d__12_ xsel_20_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN1_11 XI11_2/XI0/XI0_20/d__11_ xsel_20_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN1_10 XI11_2/XI0/XI0_20/d__10_ xsel_20_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN1_9 XI11_2/XI0/XI0_20/d__9_ xsel_20_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN1_8 XI11_2/XI0/XI0_20/d__8_ xsel_20_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN1_7 XI11_2/XI0/XI0_20/d__7_ xsel_20_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN1_6 XI11_2/XI0/XI0_20/d__6_ xsel_20_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN1_5 XI11_2/XI0/XI0_20/d__5_ xsel_20_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN1_4 XI11_2/XI0/XI0_20/d__4_ xsel_20_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN1_3 XI11_2/XI0/XI0_20/d__3_ xsel_20_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN1_2 XI11_2/XI0/XI0_20/d__2_ xsel_20_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN1_1 XI11_2/XI0/XI0_20/d__1_ xsel_20_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_20/MN1_0 XI11_2/XI0/XI0_20/d__0_ xsel_20_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN0_15 XI11_2/net21_0_ xsel_19_ XI11_2/XI0/XI0_19/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN0_14 XI11_2/net21_1_ xsel_19_ XI11_2/XI0/XI0_19/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN0_13 XI11_2/net21_2_ xsel_19_ XI11_2/XI0/XI0_19/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN0_12 XI11_2/net21_3_ xsel_19_ XI11_2/XI0/XI0_19/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN0_11 XI11_2/net21_4_ xsel_19_ XI11_2/XI0/XI0_19/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN0_10 XI11_2/net21_5_ xsel_19_ XI11_2/XI0/XI0_19/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN0_9 XI11_2/net21_6_ xsel_19_ XI11_2/XI0/XI0_19/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN0_8 XI11_2/net21_7_ xsel_19_ XI11_2/XI0/XI0_19/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN0_7 XI11_2/net21_8_ xsel_19_ XI11_2/XI0/XI0_19/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN0_6 XI11_2/net21_9_ xsel_19_ XI11_2/XI0/XI0_19/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN0_5 XI11_2/net21_10_ xsel_19_ XI11_2/XI0/XI0_19/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN0_4 XI11_2/net21_11_ xsel_19_ XI11_2/XI0/XI0_19/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN0_3 XI11_2/net21_12_ xsel_19_ XI11_2/XI0/XI0_19/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN0_2 XI11_2/net21_13_ xsel_19_ XI11_2/XI0/XI0_19/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN0_1 XI11_2/net21_14_ xsel_19_ XI11_2/XI0/XI0_19/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN0_0 XI11_2/net21_15_ xsel_19_ XI11_2/XI0/XI0_19/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN1_15 XI11_2/XI0/XI0_19/d__15_ xsel_19_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN1_14 XI11_2/XI0/XI0_19/d__14_ xsel_19_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN1_13 XI11_2/XI0/XI0_19/d__13_ xsel_19_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN1_12 XI11_2/XI0/XI0_19/d__12_ xsel_19_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN1_11 XI11_2/XI0/XI0_19/d__11_ xsel_19_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN1_10 XI11_2/XI0/XI0_19/d__10_ xsel_19_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN1_9 XI11_2/XI0/XI0_19/d__9_ xsel_19_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN1_8 XI11_2/XI0/XI0_19/d__8_ xsel_19_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN1_7 XI11_2/XI0/XI0_19/d__7_ xsel_19_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN1_6 XI11_2/XI0/XI0_19/d__6_ xsel_19_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN1_5 XI11_2/XI0/XI0_19/d__5_ xsel_19_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN1_4 XI11_2/XI0/XI0_19/d__4_ xsel_19_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN1_3 XI11_2/XI0/XI0_19/d__3_ xsel_19_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN1_2 XI11_2/XI0/XI0_19/d__2_ xsel_19_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN1_1 XI11_2/XI0/XI0_19/d__1_ xsel_19_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_19/MN1_0 XI11_2/XI0/XI0_19/d__0_ xsel_19_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN0_15 XI11_2/net21_0_ xsel_18_ XI11_2/XI0/XI0_18/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN0_14 XI11_2/net21_1_ xsel_18_ XI11_2/XI0/XI0_18/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN0_13 XI11_2/net21_2_ xsel_18_ XI11_2/XI0/XI0_18/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN0_12 XI11_2/net21_3_ xsel_18_ XI11_2/XI0/XI0_18/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN0_11 XI11_2/net21_4_ xsel_18_ XI11_2/XI0/XI0_18/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN0_10 XI11_2/net21_5_ xsel_18_ XI11_2/XI0/XI0_18/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN0_9 XI11_2/net21_6_ xsel_18_ XI11_2/XI0/XI0_18/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN0_8 XI11_2/net21_7_ xsel_18_ XI11_2/XI0/XI0_18/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN0_7 XI11_2/net21_8_ xsel_18_ XI11_2/XI0/XI0_18/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN0_6 XI11_2/net21_9_ xsel_18_ XI11_2/XI0/XI0_18/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN0_5 XI11_2/net21_10_ xsel_18_ XI11_2/XI0/XI0_18/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN0_4 XI11_2/net21_11_ xsel_18_ XI11_2/XI0/XI0_18/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN0_3 XI11_2/net21_12_ xsel_18_ XI11_2/XI0/XI0_18/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN0_2 XI11_2/net21_13_ xsel_18_ XI11_2/XI0/XI0_18/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN0_1 XI11_2/net21_14_ xsel_18_ XI11_2/XI0/XI0_18/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN0_0 XI11_2/net21_15_ xsel_18_ XI11_2/XI0/XI0_18/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN1_15 XI11_2/XI0/XI0_18/d__15_ xsel_18_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN1_14 XI11_2/XI0/XI0_18/d__14_ xsel_18_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN1_13 XI11_2/XI0/XI0_18/d__13_ xsel_18_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN1_12 XI11_2/XI0/XI0_18/d__12_ xsel_18_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN1_11 XI11_2/XI0/XI0_18/d__11_ xsel_18_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN1_10 XI11_2/XI0/XI0_18/d__10_ xsel_18_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN1_9 XI11_2/XI0/XI0_18/d__9_ xsel_18_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN1_8 XI11_2/XI0/XI0_18/d__8_ xsel_18_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN1_7 XI11_2/XI0/XI0_18/d__7_ xsel_18_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN1_6 XI11_2/XI0/XI0_18/d__6_ xsel_18_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN1_5 XI11_2/XI0/XI0_18/d__5_ xsel_18_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN1_4 XI11_2/XI0/XI0_18/d__4_ xsel_18_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN1_3 XI11_2/XI0/XI0_18/d__3_ xsel_18_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN1_2 XI11_2/XI0/XI0_18/d__2_ xsel_18_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN1_1 XI11_2/XI0/XI0_18/d__1_ xsel_18_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_18/MN1_0 XI11_2/XI0/XI0_18/d__0_ xsel_18_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN0_15 XI11_2/net21_0_ xsel_17_ XI11_2/XI0/XI0_17/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN0_14 XI11_2/net21_1_ xsel_17_ XI11_2/XI0/XI0_17/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN0_13 XI11_2/net21_2_ xsel_17_ XI11_2/XI0/XI0_17/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN0_12 XI11_2/net21_3_ xsel_17_ XI11_2/XI0/XI0_17/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN0_11 XI11_2/net21_4_ xsel_17_ XI11_2/XI0/XI0_17/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN0_10 XI11_2/net21_5_ xsel_17_ XI11_2/XI0/XI0_17/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN0_9 XI11_2/net21_6_ xsel_17_ XI11_2/XI0/XI0_17/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN0_8 XI11_2/net21_7_ xsel_17_ XI11_2/XI0/XI0_17/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN0_7 XI11_2/net21_8_ xsel_17_ XI11_2/XI0/XI0_17/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN0_6 XI11_2/net21_9_ xsel_17_ XI11_2/XI0/XI0_17/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN0_5 XI11_2/net21_10_ xsel_17_ XI11_2/XI0/XI0_17/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN0_4 XI11_2/net21_11_ xsel_17_ XI11_2/XI0/XI0_17/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN0_3 XI11_2/net21_12_ xsel_17_ XI11_2/XI0/XI0_17/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN0_2 XI11_2/net21_13_ xsel_17_ XI11_2/XI0/XI0_17/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN0_1 XI11_2/net21_14_ xsel_17_ XI11_2/XI0/XI0_17/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN0_0 XI11_2/net21_15_ xsel_17_ XI11_2/XI0/XI0_17/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN1_15 XI11_2/XI0/XI0_17/d__15_ xsel_17_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN1_14 XI11_2/XI0/XI0_17/d__14_ xsel_17_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN1_13 XI11_2/XI0/XI0_17/d__13_ xsel_17_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN1_12 XI11_2/XI0/XI0_17/d__12_ xsel_17_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN1_11 XI11_2/XI0/XI0_17/d__11_ xsel_17_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN1_10 XI11_2/XI0/XI0_17/d__10_ xsel_17_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN1_9 XI11_2/XI0/XI0_17/d__9_ xsel_17_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN1_8 XI11_2/XI0/XI0_17/d__8_ xsel_17_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN1_7 XI11_2/XI0/XI0_17/d__7_ xsel_17_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN1_6 XI11_2/XI0/XI0_17/d__6_ xsel_17_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN1_5 XI11_2/XI0/XI0_17/d__5_ xsel_17_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN1_4 XI11_2/XI0/XI0_17/d__4_ xsel_17_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN1_3 XI11_2/XI0/XI0_17/d__3_ xsel_17_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN1_2 XI11_2/XI0/XI0_17/d__2_ xsel_17_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN1_1 XI11_2/XI0/XI0_17/d__1_ xsel_17_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_17/MN1_0 XI11_2/XI0/XI0_17/d__0_ xsel_17_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN0_15 XI11_2/net21_0_ xsel_16_ XI11_2/XI0/XI0_16/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN0_14 XI11_2/net21_1_ xsel_16_ XI11_2/XI0/XI0_16/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN0_13 XI11_2/net21_2_ xsel_16_ XI11_2/XI0/XI0_16/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN0_12 XI11_2/net21_3_ xsel_16_ XI11_2/XI0/XI0_16/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN0_11 XI11_2/net21_4_ xsel_16_ XI11_2/XI0/XI0_16/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN0_10 XI11_2/net21_5_ xsel_16_ XI11_2/XI0/XI0_16/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN0_9 XI11_2/net21_6_ xsel_16_ XI11_2/XI0/XI0_16/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN0_8 XI11_2/net21_7_ xsel_16_ XI11_2/XI0/XI0_16/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN0_7 XI11_2/net21_8_ xsel_16_ XI11_2/XI0/XI0_16/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN0_6 XI11_2/net21_9_ xsel_16_ XI11_2/XI0/XI0_16/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN0_5 XI11_2/net21_10_ xsel_16_ XI11_2/XI0/XI0_16/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN0_4 XI11_2/net21_11_ xsel_16_ XI11_2/XI0/XI0_16/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN0_3 XI11_2/net21_12_ xsel_16_ XI11_2/XI0/XI0_16/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN0_2 XI11_2/net21_13_ xsel_16_ XI11_2/XI0/XI0_16/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN0_1 XI11_2/net21_14_ xsel_16_ XI11_2/XI0/XI0_16/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN0_0 XI11_2/net21_15_ xsel_16_ XI11_2/XI0/XI0_16/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN1_15 XI11_2/XI0/XI0_16/d__15_ xsel_16_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN1_14 XI11_2/XI0/XI0_16/d__14_ xsel_16_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN1_13 XI11_2/XI0/XI0_16/d__13_ xsel_16_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN1_12 XI11_2/XI0/XI0_16/d__12_ xsel_16_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN1_11 XI11_2/XI0/XI0_16/d__11_ xsel_16_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN1_10 XI11_2/XI0/XI0_16/d__10_ xsel_16_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN1_9 XI11_2/XI0/XI0_16/d__9_ xsel_16_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN1_8 XI11_2/XI0/XI0_16/d__8_ xsel_16_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN1_7 XI11_2/XI0/XI0_16/d__7_ xsel_16_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN1_6 XI11_2/XI0/XI0_16/d__6_ xsel_16_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN1_5 XI11_2/XI0/XI0_16/d__5_ xsel_16_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN1_4 XI11_2/XI0/XI0_16/d__4_ xsel_16_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN1_3 XI11_2/XI0/XI0_16/d__3_ xsel_16_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN1_2 XI11_2/XI0/XI0_16/d__2_ xsel_16_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN1_1 XI11_2/XI0/XI0_16/d__1_ xsel_16_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_16/MN1_0 XI11_2/XI0/XI0_16/d__0_ xsel_16_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN0_15 XI11_2/net21_0_ xsel_15_ XI11_2/XI0/XI0_15/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN0_14 XI11_2/net21_1_ xsel_15_ XI11_2/XI0/XI0_15/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN0_13 XI11_2/net21_2_ xsel_15_ XI11_2/XI0/XI0_15/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN0_12 XI11_2/net21_3_ xsel_15_ XI11_2/XI0/XI0_15/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN0_11 XI11_2/net21_4_ xsel_15_ XI11_2/XI0/XI0_15/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN0_10 XI11_2/net21_5_ xsel_15_ XI11_2/XI0/XI0_15/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN0_9 XI11_2/net21_6_ xsel_15_ XI11_2/XI0/XI0_15/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN0_8 XI11_2/net21_7_ xsel_15_ XI11_2/XI0/XI0_15/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN0_7 XI11_2/net21_8_ xsel_15_ XI11_2/XI0/XI0_15/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN0_6 XI11_2/net21_9_ xsel_15_ XI11_2/XI0/XI0_15/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN0_5 XI11_2/net21_10_ xsel_15_ XI11_2/XI0/XI0_15/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN0_4 XI11_2/net21_11_ xsel_15_ XI11_2/XI0/XI0_15/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN0_3 XI11_2/net21_12_ xsel_15_ XI11_2/XI0/XI0_15/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN0_2 XI11_2/net21_13_ xsel_15_ XI11_2/XI0/XI0_15/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN0_1 XI11_2/net21_14_ xsel_15_ XI11_2/XI0/XI0_15/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN0_0 XI11_2/net21_15_ xsel_15_ XI11_2/XI0/XI0_15/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN1_15 XI11_2/XI0/XI0_15/d__15_ xsel_15_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN1_14 XI11_2/XI0/XI0_15/d__14_ xsel_15_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN1_13 XI11_2/XI0/XI0_15/d__13_ xsel_15_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN1_12 XI11_2/XI0/XI0_15/d__12_ xsel_15_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN1_11 XI11_2/XI0/XI0_15/d__11_ xsel_15_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN1_10 XI11_2/XI0/XI0_15/d__10_ xsel_15_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN1_9 XI11_2/XI0/XI0_15/d__9_ xsel_15_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN1_8 XI11_2/XI0/XI0_15/d__8_ xsel_15_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN1_7 XI11_2/XI0/XI0_15/d__7_ xsel_15_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN1_6 XI11_2/XI0/XI0_15/d__6_ xsel_15_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN1_5 XI11_2/XI0/XI0_15/d__5_ xsel_15_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN1_4 XI11_2/XI0/XI0_15/d__4_ xsel_15_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN1_3 XI11_2/XI0/XI0_15/d__3_ xsel_15_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN1_2 XI11_2/XI0/XI0_15/d__2_ xsel_15_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN1_1 XI11_2/XI0/XI0_15/d__1_ xsel_15_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_15/MN1_0 XI11_2/XI0/XI0_15/d__0_ xsel_15_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN0_15 XI11_2/net21_0_ xsel_14_ XI11_2/XI0/XI0_14/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN0_14 XI11_2/net21_1_ xsel_14_ XI11_2/XI0/XI0_14/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN0_13 XI11_2/net21_2_ xsel_14_ XI11_2/XI0/XI0_14/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN0_12 XI11_2/net21_3_ xsel_14_ XI11_2/XI0/XI0_14/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN0_11 XI11_2/net21_4_ xsel_14_ XI11_2/XI0/XI0_14/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN0_10 XI11_2/net21_5_ xsel_14_ XI11_2/XI0/XI0_14/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN0_9 XI11_2/net21_6_ xsel_14_ XI11_2/XI0/XI0_14/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN0_8 XI11_2/net21_7_ xsel_14_ XI11_2/XI0/XI0_14/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN0_7 XI11_2/net21_8_ xsel_14_ XI11_2/XI0/XI0_14/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN0_6 XI11_2/net21_9_ xsel_14_ XI11_2/XI0/XI0_14/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN0_5 XI11_2/net21_10_ xsel_14_ XI11_2/XI0/XI0_14/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN0_4 XI11_2/net21_11_ xsel_14_ XI11_2/XI0/XI0_14/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN0_3 XI11_2/net21_12_ xsel_14_ XI11_2/XI0/XI0_14/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN0_2 XI11_2/net21_13_ xsel_14_ XI11_2/XI0/XI0_14/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN0_1 XI11_2/net21_14_ xsel_14_ XI11_2/XI0/XI0_14/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN0_0 XI11_2/net21_15_ xsel_14_ XI11_2/XI0/XI0_14/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN1_15 XI11_2/XI0/XI0_14/d__15_ xsel_14_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN1_14 XI11_2/XI0/XI0_14/d__14_ xsel_14_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN1_13 XI11_2/XI0/XI0_14/d__13_ xsel_14_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN1_12 XI11_2/XI0/XI0_14/d__12_ xsel_14_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN1_11 XI11_2/XI0/XI0_14/d__11_ xsel_14_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN1_10 XI11_2/XI0/XI0_14/d__10_ xsel_14_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN1_9 XI11_2/XI0/XI0_14/d__9_ xsel_14_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN1_8 XI11_2/XI0/XI0_14/d__8_ xsel_14_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN1_7 XI11_2/XI0/XI0_14/d__7_ xsel_14_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN1_6 XI11_2/XI0/XI0_14/d__6_ xsel_14_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN1_5 XI11_2/XI0/XI0_14/d__5_ xsel_14_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN1_4 XI11_2/XI0/XI0_14/d__4_ xsel_14_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN1_3 XI11_2/XI0/XI0_14/d__3_ xsel_14_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN1_2 XI11_2/XI0/XI0_14/d__2_ xsel_14_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN1_1 XI11_2/XI0/XI0_14/d__1_ xsel_14_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_14/MN1_0 XI11_2/XI0/XI0_14/d__0_ xsel_14_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN0_15 XI11_2/net21_0_ xsel_13_ XI11_2/XI0/XI0_13/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN0_14 XI11_2/net21_1_ xsel_13_ XI11_2/XI0/XI0_13/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN0_13 XI11_2/net21_2_ xsel_13_ XI11_2/XI0/XI0_13/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN0_12 XI11_2/net21_3_ xsel_13_ XI11_2/XI0/XI0_13/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN0_11 XI11_2/net21_4_ xsel_13_ XI11_2/XI0/XI0_13/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN0_10 XI11_2/net21_5_ xsel_13_ XI11_2/XI0/XI0_13/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN0_9 XI11_2/net21_6_ xsel_13_ XI11_2/XI0/XI0_13/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN0_8 XI11_2/net21_7_ xsel_13_ XI11_2/XI0/XI0_13/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN0_7 XI11_2/net21_8_ xsel_13_ XI11_2/XI0/XI0_13/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN0_6 XI11_2/net21_9_ xsel_13_ XI11_2/XI0/XI0_13/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN0_5 XI11_2/net21_10_ xsel_13_ XI11_2/XI0/XI0_13/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN0_4 XI11_2/net21_11_ xsel_13_ XI11_2/XI0/XI0_13/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN0_3 XI11_2/net21_12_ xsel_13_ XI11_2/XI0/XI0_13/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN0_2 XI11_2/net21_13_ xsel_13_ XI11_2/XI0/XI0_13/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN0_1 XI11_2/net21_14_ xsel_13_ XI11_2/XI0/XI0_13/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN0_0 XI11_2/net21_15_ xsel_13_ XI11_2/XI0/XI0_13/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN1_15 XI11_2/XI0/XI0_13/d__15_ xsel_13_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN1_14 XI11_2/XI0/XI0_13/d__14_ xsel_13_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN1_13 XI11_2/XI0/XI0_13/d__13_ xsel_13_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN1_12 XI11_2/XI0/XI0_13/d__12_ xsel_13_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN1_11 XI11_2/XI0/XI0_13/d__11_ xsel_13_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN1_10 XI11_2/XI0/XI0_13/d__10_ xsel_13_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN1_9 XI11_2/XI0/XI0_13/d__9_ xsel_13_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN1_8 XI11_2/XI0/XI0_13/d__8_ xsel_13_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN1_7 XI11_2/XI0/XI0_13/d__7_ xsel_13_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN1_6 XI11_2/XI0/XI0_13/d__6_ xsel_13_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN1_5 XI11_2/XI0/XI0_13/d__5_ xsel_13_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN1_4 XI11_2/XI0/XI0_13/d__4_ xsel_13_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN1_3 XI11_2/XI0/XI0_13/d__3_ xsel_13_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN1_2 XI11_2/XI0/XI0_13/d__2_ xsel_13_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN1_1 XI11_2/XI0/XI0_13/d__1_ xsel_13_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_13/MN1_0 XI11_2/XI0/XI0_13/d__0_ xsel_13_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN0_15 XI11_2/net21_0_ xsel_12_ XI11_2/XI0/XI0_12/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN0_14 XI11_2/net21_1_ xsel_12_ XI11_2/XI0/XI0_12/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN0_13 XI11_2/net21_2_ xsel_12_ XI11_2/XI0/XI0_12/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN0_12 XI11_2/net21_3_ xsel_12_ XI11_2/XI0/XI0_12/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN0_11 XI11_2/net21_4_ xsel_12_ XI11_2/XI0/XI0_12/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN0_10 XI11_2/net21_5_ xsel_12_ XI11_2/XI0/XI0_12/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN0_9 XI11_2/net21_6_ xsel_12_ XI11_2/XI0/XI0_12/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN0_8 XI11_2/net21_7_ xsel_12_ XI11_2/XI0/XI0_12/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN0_7 XI11_2/net21_8_ xsel_12_ XI11_2/XI0/XI0_12/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN0_6 XI11_2/net21_9_ xsel_12_ XI11_2/XI0/XI0_12/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN0_5 XI11_2/net21_10_ xsel_12_ XI11_2/XI0/XI0_12/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN0_4 XI11_2/net21_11_ xsel_12_ XI11_2/XI0/XI0_12/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN0_3 XI11_2/net21_12_ xsel_12_ XI11_2/XI0/XI0_12/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN0_2 XI11_2/net21_13_ xsel_12_ XI11_2/XI0/XI0_12/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN0_1 XI11_2/net21_14_ xsel_12_ XI11_2/XI0/XI0_12/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN0_0 XI11_2/net21_15_ xsel_12_ XI11_2/XI0/XI0_12/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN1_15 XI11_2/XI0/XI0_12/d__15_ xsel_12_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN1_14 XI11_2/XI0/XI0_12/d__14_ xsel_12_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN1_13 XI11_2/XI0/XI0_12/d__13_ xsel_12_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN1_12 XI11_2/XI0/XI0_12/d__12_ xsel_12_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN1_11 XI11_2/XI0/XI0_12/d__11_ xsel_12_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN1_10 XI11_2/XI0/XI0_12/d__10_ xsel_12_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN1_9 XI11_2/XI0/XI0_12/d__9_ xsel_12_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN1_8 XI11_2/XI0/XI0_12/d__8_ xsel_12_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN1_7 XI11_2/XI0/XI0_12/d__7_ xsel_12_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN1_6 XI11_2/XI0/XI0_12/d__6_ xsel_12_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN1_5 XI11_2/XI0/XI0_12/d__5_ xsel_12_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN1_4 XI11_2/XI0/XI0_12/d__4_ xsel_12_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN1_3 XI11_2/XI0/XI0_12/d__3_ xsel_12_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN1_2 XI11_2/XI0/XI0_12/d__2_ xsel_12_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN1_1 XI11_2/XI0/XI0_12/d__1_ xsel_12_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_12/MN1_0 XI11_2/XI0/XI0_12/d__0_ xsel_12_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN0_15 XI11_2/net21_0_ xsel_11_ XI11_2/XI0/XI0_11/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN0_14 XI11_2/net21_1_ xsel_11_ XI11_2/XI0/XI0_11/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN0_13 XI11_2/net21_2_ xsel_11_ XI11_2/XI0/XI0_11/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN0_12 XI11_2/net21_3_ xsel_11_ XI11_2/XI0/XI0_11/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN0_11 XI11_2/net21_4_ xsel_11_ XI11_2/XI0/XI0_11/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN0_10 XI11_2/net21_5_ xsel_11_ XI11_2/XI0/XI0_11/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN0_9 XI11_2/net21_6_ xsel_11_ XI11_2/XI0/XI0_11/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN0_8 XI11_2/net21_7_ xsel_11_ XI11_2/XI0/XI0_11/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN0_7 XI11_2/net21_8_ xsel_11_ XI11_2/XI0/XI0_11/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN0_6 XI11_2/net21_9_ xsel_11_ XI11_2/XI0/XI0_11/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN0_5 XI11_2/net21_10_ xsel_11_ XI11_2/XI0/XI0_11/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN0_4 XI11_2/net21_11_ xsel_11_ XI11_2/XI0/XI0_11/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN0_3 XI11_2/net21_12_ xsel_11_ XI11_2/XI0/XI0_11/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN0_2 XI11_2/net21_13_ xsel_11_ XI11_2/XI0/XI0_11/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN0_1 XI11_2/net21_14_ xsel_11_ XI11_2/XI0/XI0_11/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN0_0 XI11_2/net21_15_ xsel_11_ XI11_2/XI0/XI0_11/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN1_15 XI11_2/XI0/XI0_11/d__15_ xsel_11_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN1_14 XI11_2/XI0/XI0_11/d__14_ xsel_11_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN1_13 XI11_2/XI0/XI0_11/d__13_ xsel_11_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN1_12 XI11_2/XI0/XI0_11/d__12_ xsel_11_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN1_11 XI11_2/XI0/XI0_11/d__11_ xsel_11_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN1_10 XI11_2/XI0/XI0_11/d__10_ xsel_11_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN1_9 XI11_2/XI0/XI0_11/d__9_ xsel_11_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN1_8 XI11_2/XI0/XI0_11/d__8_ xsel_11_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN1_7 XI11_2/XI0/XI0_11/d__7_ xsel_11_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN1_6 XI11_2/XI0/XI0_11/d__6_ xsel_11_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN1_5 XI11_2/XI0/XI0_11/d__5_ xsel_11_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN1_4 XI11_2/XI0/XI0_11/d__4_ xsel_11_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN1_3 XI11_2/XI0/XI0_11/d__3_ xsel_11_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN1_2 XI11_2/XI0/XI0_11/d__2_ xsel_11_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN1_1 XI11_2/XI0/XI0_11/d__1_ xsel_11_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_11/MN1_0 XI11_2/XI0/XI0_11/d__0_ xsel_11_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN0_15 XI11_2/net21_0_ xsel_10_ XI11_2/XI0/XI0_10/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN0_14 XI11_2/net21_1_ xsel_10_ XI11_2/XI0/XI0_10/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN0_13 XI11_2/net21_2_ xsel_10_ XI11_2/XI0/XI0_10/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN0_12 XI11_2/net21_3_ xsel_10_ XI11_2/XI0/XI0_10/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN0_11 XI11_2/net21_4_ xsel_10_ XI11_2/XI0/XI0_10/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN0_10 XI11_2/net21_5_ xsel_10_ XI11_2/XI0/XI0_10/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN0_9 XI11_2/net21_6_ xsel_10_ XI11_2/XI0/XI0_10/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN0_8 XI11_2/net21_7_ xsel_10_ XI11_2/XI0/XI0_10/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN0_7 XI11_2/net21_8_ xsel_10_ XI11_2/XI0/XI0_10/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN0_6 XI11_2/net21_9_ xsel_10_ XI11_2/XI0/XI0_10/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN0_5 XI11_2/net21_10_ xsel_10_ XI11_2/XI0/XI0_10/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN0_4 XI11_2/net21_11_ xsel_10_ XI11_2/XI0/XI0_10/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN0_3 XI11_2/net21_12_ xsel_10_ XI11_2/XI0/XI0_10/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN0_2 XI11_2/net21_13_ xsel_10_ XI11_2/XI0/XI0_10/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN0_1 XI11_2/net21_14_ xsel_10_ XI11_2/XI0/XI0_10/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN0_0 XI11_2/net21_15_ xsel_10_ XI11_2/XI0/XI0_10/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN1_15 XI11_2/XI0/XI0_10/d__15_ xsel_10_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN1_14 XI11_2/XI0/XI0_10/d__14_ xsel_10_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN1_13 XI11_2/XI0/XI0_10/d__13_ xsel_10_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN1_12 XI11_2/XI0/XI0_10/d__12_ xsel_10_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN1_11 XI11_2/XI0/XI0_10/d__11_ xsel_10_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN1_10 XI11_2/XI0/XI0_10/d__10_ xsel_10_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN1_9 XI11_2/XI0/XI0_10/d__9_ xsel_10_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN1_8 XI11_2/XI0/XI0_10/d__8_ xsel_10_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN1_7 XI11_2/XI0/XI0_10/d__7_ xsel_10_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN1_6 XI11_2/XI0/XI0_10/d__6_ xsel_10_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN1_5 XI11_2/XI0/XI0_10/d__5_ xsel_10_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN1_4 XI11_2/XI0/XI0_10/d__4_ xsel_10_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN1_3 XI11_2/XI0/XI0_10/d__3_ xsel_10_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN1_2 XI11_2/XI0/XI0_10/d__2_ xsel_10_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN1_1 XI11_2/XI0/XI0_10/d__1_ xsel_10_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_10/MN1_0 XI11_2/XI0/XI0_10/d__0_ xsel_10_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN0_15 XI11_2/net21_0_ xsel_9_ XI11_2/XI0/XI0_9/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN0_14 XI11_2/net21_1_ xsel_9_ XI11_2/XI0/XI0_9/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN0_13 XI11_2/net21_2_ xsel_9_ XI11_2/XI0/XI0_9/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN0_12 XI11_2/net21_3_ xsel_9_ XI11_2/XI0/XI0_9/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN0_11 XI11_2/net21_4_ xsel_9_ XI11_2/XI0/XI0_9/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN0_10 XI11_2/net21_5_ xsel_9_ XI11_2/XI0/XI0_9/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN0_9 XI11_2/net21_6_ xsel_9_ XI11_2/XI0/XI0_9/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN0_8 XI11_2/net21_7_ xsel_9_ XI11_2/XI0/XI0_9/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN0_7 XI11_2/net21_8_ xsel_9_ XI11_2/XI0/XI0_9/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN0_6 XI11_2/net21_9_ xsel_9_ XI11_2/XI0/XI0_9/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN0_5 XI11_2/net21_10_ xsel_9_ XI11_2/XI0/XI0_9/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN0_4 XI11_2/net21_11_ xsel_9_ XI11_2/XI0/XI0_9/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN0_3 XI11_2/net21_12_ xsel_9_ XI11_2/XI0/XI0_9/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN0_2 XI11_2/net21_13_ xsel_9_ XI11_2/XI0/XI0_9/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN0_1 XI11_2/net21_14_ xsel_9_ XI11_2/XI0/XI0_9/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN0_0 XI11_2/net21_15_ xsel_9_ XI11_2/XI0/XI0_9/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN1_15 XI11_2/XI0/XI0_9/d__15_ xsel_9_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN1_14 XI11_2/XI0/XI0_9/d__14_ xsel_9_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN1_13 XI11_2/XI0/XI0_9/d__13_ xsel_9_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN1_12 XI11_2/XI0/XI0_9/d__12_ xsel_9_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN1_11 XI11_2/XI0/XI0_9/d__11_ xsel_9_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN1_10 XI11_2/XI0/XI0_9/d__10_ xsel_9_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN1_9 XI11_2/XI0/XI0_9/d__9_ xsel_9_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN1_8 XI11_2/XI0/XI0_9/d__8_ xsel_9_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN1_7 XI11_2/XI0/XI0_9/d__7_ xsel_9_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN1_6 XI11_2/XI0/XI0_9/d__6_ xsel_9_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN1_5 XI11_2/XI0/XI0_9/d__5_ xsel_9_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN1_4 XI11_2/XI0/XI0_9/d__4_ xsel_9_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN1_3 XI11_2/XI0/XI0_9/d__3_ xsel_9_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN1_2 XI11_2/XI0/XI0_9/d__2_ xsel_9_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN1_1 XI11_2/XI0/XI0_9/d__1_ xsel_9_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_9/MN1_0 XI11_2/XI0/XI0_9/d__0_ xsel_9_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN0_15 XI11_2/net21_0_ xsel_8_ XI11_2/XI0/XI0_8/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN0_14 XI11_2/net21_1_ xsel_8_ XI11_2/XI0/XI0_8/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN0_13 XI11_2/net21_2_ xsel_8_ XI11_2/XI0/XI0_8/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN0_12 XI11_2/net21_3_ xsel_8_ XI11_2/XI0/XI0_8/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN0_11 XI11_2/net21_4_ xsel_8_ XI11_2/XI0/XI0_8/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN0_10 XI11_2/net21_5_ xsel_8_ XI11_2/XI0/XI0_8/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN0_9 XI11_2/net21_6_ xsel_8_ XI11_2/XI0/XI0_8/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN0_8 XI11_2/net21_7_ xsel_8_ XI11_2/XI0/XI0_8/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN0_7 XI11_2/net21_8_ xsel_8_ XI11_2/XI0/XI0_8/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN0_6 XI11_2/net21_9_ xsel_8_ XI11_2/XI0/XI0_8/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN0_5 XI11_2/net21_10_ xsel_8_ XI11_2/XI0/XI0_8/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN0_4 XI11_2/net21_11_ xsel_8_ XI11_2/XI0/XI0_8/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN0_3 XI11_2/net21_12_ xsel_8_ XI11_2/XI0/XI0_8/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN0_2 XI11_2/net21_13_ xsel_8_ XI11_2/XI0/XI0_8/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN0_1 XI11_2/net21_14_ xsel_8_ XI11_2/XI0/XI0_8/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN0_0 XI11_2/net21_15_ xsel_8_ XI11_2/XI0/XI0_8/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN1_15 XI11_2/XI0/XI0_8/d__15_ xsel_8_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN1_14 XI11_2/XI0/XI0_8/d__14_ xsel_8_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN1_13 XI11_2/XI0/XI0_8/d__13_ xsel_8_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN1_12 XI11_2/XI0/XI0_8/d__12_ xsel_8_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN1_11 XI11_2/XI0/XI0_8/d__11_ xsel_8_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN1_10 XI11_2/XI0/XI0_8/d__10_ xsel_8_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN1_9 XI11_2/XI0/XI0_8/d__9_ xsel_8_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN1_8 XI11_2/XI0/XI0_8/d__8_ xsel_8_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN1_7 XI11_2/XI0/XI0_8/d__7_ xsel_8_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN1_6 XI11_2/XI0/XI0_8/d__6_ xsel_8_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN1_5 XI11_2/XI0/XI0_8/d__5_ xsel_8_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN1_4 XI11_2/XI0/XI0_8/d__4_ xsel_8_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN1_3 XI11_2/XI0/XI0_8/d__3_ xsel_8_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN1_2 XI11_2/XI0/XI0_8/d__2_ xsel_8_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN1_1 XI11_2/XI0/XI0_8/d__1_ xsel_8_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_8/MN1_0 XI11_2/XI0/XI0_8/d__0_ xsel_8_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN0_15 XI11_2/net21_0_ xsel_7_ XI11_2/XI0/XI0_7/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN0_14 XI11_2/net21_1_ xsel_7_ XI11_2/XI0/XI0_7/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN0_13 XI11_2/net21_2_ xsel_7_ XI11_2/XI0/XI0_7/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN0_12 XI11_2/net21_3_ xsel_7_ XI11_2/XI0/XI0_7/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN0_11 XI11_2/net21_4_ xsel_7_ XI11_2/XI0/XI0_7/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN0_10 XI11_2/net21_5_ xsel_7_ XI11_2/XI0/XI0_7/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN0_9 XI11_2/net21_6_ xsel_7_ XI11_2/XI0/XI0_7/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN0_8 XI11_2/net21_7_ xsel_7_ XI11_2/XI0/XI0_7/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN0_7 XI11_2/net21_8_ xsel_7_ XI11_2/XI0/XI0_7/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN0_6 XI11_2/net21_9_ xsel_7_ XI11_2/XI0/XI0_7/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN0_5 XI11_2/net21_10_ xsel_7_ XI11_2/XI0/XI0_7/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN0_4 XI11_2/net21_11_ xsel_7_ XI11_2/XI0/XI0_7/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN0_3 XI11_2/net21_12_ xsel_7_ XI11_2/XI0/XI0_7/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN0_2 XI11_2/net21_13_ xsel_7_ XI11_2/XI0/XI0_7/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN0_1 XI11_2/net21_14_ xsel_7_ XI11_2/XI0/XI0_7/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN0_0 XI11_2/net21_15_ xsel_7_ XI11_2/XI0/XI0_7/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN1_15 XI11_2/XI0/XI0_7/d__15_ xsel_7_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN1_14 XI11_2/XI0/XI0_7/d__14_ xsel_7_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN1_13 XI11_2/XI0/XI0_7/d__13_ xsel_7_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN1_12 XI11_2/XI0/XI0_7/d__12_ xsel_7_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN1_11 XI11_2/XI0/XI0_7/d__11_ xsel_7_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN1_10 XI11_2/XI0/XI0_7/d__10_ xsel_7_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN1_9 XI11_2/XI0/XI0_7/d__9_ xsel_7_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN1_8 XI11_2/XI0/XI0_7/d__8_ xsel_7_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN1_7 XI11_2/XI0/XI0_7/d__7_ xsel_7_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN1_6 XI11_2/XI0/XI0_7/d__6_ xsel_7_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN1_5 XI11_2/XI0/XI0_7/d__5_ xsel_7_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN1_4 XI11_2/XI0/XI0_7/d__4_ xsel_7_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN1_3 XI11_2/XI0/XI0_7/d__3_ xsel_7_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN1_2 XI11_2/XI0/XI0_7/d__2_ xsel_7_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN1_1 XI11_2/XI0/XI0_7/d__1_ xsel_7_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_7/MN1_0 XI11_2/XI0/XI0_7/d__0_ xsel_7_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN0_15 XI11_2/net21_0_ xsel_6_ XI11_2/XI0/XI0_6/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN0_14 XI11_2/net21_1_ xsel_6_ XI11_2/XI0/XI0_6/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN0_13 XI11_2/net21_2_ xsel_6_ XI11_2/XI0/XI0_6/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN0_12 XI11_2/net21_3_ xsel_6_ XI11_2/XI0/XI0_6/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN0_11 XI11_2/net21_4_ xsel_6_ XI11_2/XI0/XI0_6/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN0_10 XI11_2/net21_5_ xsel_6_ XI11_2/XI0/XI0_6/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN0_9 XI11_2/net21_6_ xsel_6_ XI11_2/XI0/XI0_6/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN0_8 XI11_2/net21_7_ xsel_6_ XI11_2/XI0/XI0_6/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN0_7 XI11_2/net21_8_ xsel_6_ XI11_2/XI0/XI0_6/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN0_6 XI11_2/net21_9_ xsel_6_ XI11_2/XI0/XI0_6/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN0_5 XI11_2/net21_10_ xsel_6_ XI11_2/XI0/XI0_6/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN0_4 XI11_2/net21_11_ xsel_6_ XI11_2/XI0/XI0_6/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN0_3 XI11_2/net21_12_ xsel_6_ XI11_2/XI0/XI0_6/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN0_2 XI11_2/net21_13_ xsel_6_ XI11_2/XI0/XI0_6/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN0_1 XI11_2/net21_14_ xsel_6_ XI11_2/XI0/XI0_6/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN0_0 XI11_2/net21_15_ xsel_6_ XI11_2/XI0/XI0_6/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN1_15 XI11_2/XI0/XI0_6/d__15_ xsel_6_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN1_14 XI11_2/XI0/XI0_6/d__14_ xsel_6_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN1_13 XI11_2/XI0/XI0_6/d__13_ xsel_6_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN1_12 XI11_2/XI0/XI0_6/d__12_ xsel_6_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN1_11 XI11_2/XI0/XI0_6/d__11_ xsel_6_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN1_10 XI11_2/XI0/XI0_6/d__10_ xsel_6_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN1_9 XI11_2/XI0/XI0_6/d__9_ xsel_6_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN1_8 XI11_2/XI0/XI0_6/d__8_ xsel_6_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN1_7 XI11_2/XI0/XI0_6/d__7_ xsel_6_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN1_6 XI11_2/XI0/XI0_6/d__6_ xsel_6_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN1_5 XI11_2/XI0/XI0_6/d__5_ xsel_6_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN1_4 XI11_2/XI0/XI0_6/d__4_ xsel_6_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN1_3 XI11_2/XI0/XI0_6/d__3_ xsel_6_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN1_2 XI11_2/XI0/XI0_6/d__2_ xsel_6_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN1_1 XI11_2/XI0/XI0_6/d__1_ xsel_6_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_6/MN1_0 XI11_2/XI0/XI0_6/d__0_ xsel_6_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN0_15 XI11_2/net21_0_ xsel_5_ XI11_2/XI0/XI0_5/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN0_14 XI11_2/net21_1_ xsel_5_ XI11_2/XI0/XI0_5/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN0_13 XI11_2/net21_2_ xsel_5_ XI11_2/XI0/XI0_5/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN0_12 XI11_2/net21_3_ xsel_5_ XI11_2/XI0/XI0_5/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN0_11 XI11_2/net21_4_ xsel_5_ XI11_2/XI0/XI0_5/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN0_10 XI11_2/net21_5_ xsel_5_ XI11_2/XI0/XI0_5/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN0_9 XI11_2/net21_6_ xsel_5_ XI11_2/XI0/XI0_5/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN0_8 XI11_2/net21_7_ xsel_5_ XI11_2/XI0/XI0_5/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN0_7 XI11_2/net21_8_ xsel_5_ XI11_2/XI0/XI0_5/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN0_6 XI11_2/net21_9_ xsel_5_ XI11_2/XI0/XI0_5/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN0_5 XI11_2/net21_10_ xsel_5_ XI11_2/XI0/XI0_5/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN0_4 XI11_2/net21_11_ xsel_5_ XI11_2/XI0/XI0_5/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN0_3 XI11_2/net21_12_ xsel_5_ XI11_2/XI0/XI0_5/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN0_2 XI11_2/net21_13_ xsel_5_ XI11_2/XI0/XI0_5/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN0_1 XI11_2/net21_14_ xsel_5_ XI11_2/XI0/XI0_5/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN0_0 XI11_2/net21_15_ xsel_5_ XI11_2/XI0/XI0_5/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN1_15 XI11_2/XI0/XI0_5/d__15_ xsel_5_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN1_14 XI11_2/XI0/XI0_5/d__14_ xsel_5_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN1_13 XI11_2/XI0/XI0_5/d__13_ xsel_5_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN1_12 XI11_2/XI0/XI0_5/d__12_ xsel_5_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN1_11 XI11_2/XI0/XI0_5/d__11_ xsel_5_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN1_10 XI11_2/XI0/XI0_5/d__10_ xsel_5_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN1_9 XI11_2/XI0/XI0_5/d__9_ xsel_5_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN1_8 XI11_2/XI0/XI0_5/d__8_ xsel_5_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN1_7 XI11_2/XI0/XI0_5/d__7_ xsel_5_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN1_6 XI11_2/XI0/XI0_5/d__6_ xsel_5_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN1_5 XI11_2/XI0/XI0_5/d__5_ xsel_5_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN1_4 XI11_2/XI0/XI0_5/d__4_ xsel_5_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN1_3 XI11_2/XI0/XI0_5/d__3_ xsel_5_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN1_2 XI11_2/XI0/XI0_5/d__2_ xsel_5_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN1_1 XI11_2/XI0/XI0_5/d__1_ xsel_5_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_5/MN1_0 XI11_2/XI0/XI0_5/d__0_ xsel_5_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN0_15 XI11_2/net21_0_ xsel_4_ XI11_2/XI0/XI0_4/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN0_14 XI11_2/net21_1_ xsel_4_ XI11_2/XI0/XI0_4/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN0_13 XI11_2/net21_2_ xsel_4_ XI11_2/XI0/XI0_4/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN0_12 XI11_2/net21_3_ xsel_4_ XI11_2/XI0/XI0_4/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN0_11 XI11_2/net21_4_ xsel_4_ XI11_2/XI0/XI0_4/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN0_10 XI11_2/net21_5_ xsel_4_ XI11_2/XI0/XI0_4/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN0_9 XI11_2/net21_6_ xsel_4_ XI11_2/XI0/XI0_4/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN0_8 XI11_2/net21_7_ xsel_4_ XI11_2/XI0/XI0_4/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN0_7 XI11_2/net21_8_ xsel_4_ XI11_2/XI0/XI0_4/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN0_6 XI11_2/net21_9_ xsel_4_ XI11_2/XI0/XI0_4/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN0_5 XI11_2/net21_10_ xsel_4_ XI11_2/XI0/XI0_4/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN0_4 XI11_2/net21_11_ xsel_4_ XI11_2/XI0/XI0_4/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN0_3 XI11_2/net21_12_ xsel_4_ XI11_2/XI0/XI0_4/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN0_2 XI11_2/net21_13_ xsel_4_ XI11_2/XI0/XI0_4/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN0_1 XI11_2/net21_14_ xsel_4_ XI11_2/XI0/XI0_4/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN0_0 XI11_2/net21_15_ xsel_4_ XI11_2/XI0/XI0_4/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN1_15 XI11_2/XI0/XI0_4/d__15_ xsel_4_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN1_14 XI11_2/XI0/XI0_4/d__14_ xsel_4_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN1_13 XI11_2/XI0/XI0_4/d__13_ xsel_4_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN1_12 XI11_2/XI0/XI0_4/d__12_ xsel_4_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN1_11 XI11_2/XI0/XI0_4/d__11_ xsel_4_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN1_10 XI11_2/XI0/XI0_4/d__10_ xsel_4_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN1_9 XI11_2/XI0/XI0_4/d__9_ xsel_4_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN1_8 XI11_2/XI0/XI0_4/d__8_ xsel_4_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN1_7 XI11_2/XI0/XI0_4/d__7_ xsel_4_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN1_6 XI11_2/XI0/XI0_4/d__6_ xsel_4_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN1_5 XI11_2/XI0/XI0_4/d__5_ xsel_4_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN1_4 XI11_2/XI0/XI0_4/d__4_ xsel_4_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN1_3 XI11_2/XI0/XI0_4/d__3_ xsel_4_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN1_2 XI11_2/XI0/XI0_4/d__2_ xsel_4_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN1_1 XI11_2/XI0/XI0_4/d__1_ xsel_4_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_4/MN1_0 XI11_2/XI0/XI0_4/d__0_ xsel_4_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN0_15 XI11_2/net21_0_ xsel_3_ XI11_2/XI0/XI0_3/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN0_14 XI11_2/net21_1_ xsel_3_ XI11_2/XI0/XI0_3/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN0_13 XI11_2/net21_2_ xsel_3_ XI11_2/XI0/XI0_3/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN0_12 XI11_2/net21_3_ xsel_3_ XI11_2/XI0/XI0_3/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN0_11 XI11_2/net21_4_ xsel_3_ XI11_2/XI0/XI0_3/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN0_10 XI11_2/net21_5_ xsel_3_ XI11_2/XI0/XI0_3/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN0_9 XI11_2/net21_6_ xsel_3_ XI11_2/XI0/XI0_3/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN0_8 XI11_2/net21_7_ xsel_3_ XI11_2/XI0/XI0_3/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN0_7 XI11_2/net21_8_ xsel_3_ XI11_2/XI0/XI0_3/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN0_6 XI11_2/net21_9_ xsel_3_ XI11_2/XI0/XI0_3/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN0_5 XI11_2/net21_10_ xsel_3_ XI11_2/XI0/XI0_3/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN0_4 XI11_2/net21_11_ xsel_3_ XI11_2/XI0/XI0_3/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN0_3 XI11_2/net21_12_ xsel_3_ XI11_2/XI0/XI0_3/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN0_2 XI11_2/net21_13_ xsel_3_ XI11_2/XI0/XI0_3/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN0_1 XI11_2/net21_14_ xsel_3_ XI11_2/XI0/XI0_3/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN0_0 XI11_2/net21_15_ xsel_3_ XI11_2/XI0/XI0_3/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN1_15 XI11_2/XI0/XI0_3/d__15_ xsel_3_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN1_14 XI11_2/XI0/XI0_3/d__14_ xsel_3_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN1_13 XI11_2/XI0/XI0_3/d__13_ xsel_3_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN1_12 XI11_2/XI0/XI0_3/d__12_ xsel_3_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN1_11 XI11_2/XI0/XI0_3/d__11_ xsel_3_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN1_10 XI11_2/XI0/XI0_3/d__10_ xsel_3_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN1_9 XI11_2/XI0/XI0_3/d__9_ xsel_3_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN1_8 XI11_2/XI0/XI0_3/d__8_ xsel_3_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN1_7 XI11_2/XI0/XI0_3/d__7_ xsel_3_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN1_6 XI11_2/XI0/XI0_3/d__6_ xsel_3_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN1_5 XI11_2/XI0/XI0_3/d__5_ xsel_3_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN1_4 XI11_2/XI0/XI0_3/d__4_ xsel_3_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN1_3 XI11_2/XI0/XI0_3/d__3_ xsel_3_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN1_2 XI11_2/XI0/XI0_3/d__2_ xsel_3_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN1_1 XI11_2/XI0/XI0_3/d__1_ xsel_3_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_3/MN1_0 XI11_2/XI0/XI0_3/d__0_ xsel_3_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN0_15 XI11_2/net21_0_ xsel_2_ XI11_2/XI0/XI0_2/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN0_14 XI11_2/net21_1_ xsel_2_ XI11_2/XI0/XI0_2/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN0_13 XI11_2/net21_2_ xsel_2_ XI11_2/XI0/XI0_2/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN0_12 XI11_2/net21_3_ xsel_2_ XI11_2/XI0/XI0_2/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN0_11 XI11_2/net21_4_ xsel_2_ XI11_2/XI0/XI0_2/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN0_10 XI11_2/net21_5_ xsel_2_ XI11_2/XI0/XI0_2/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN0_9 XI11_2/net21_6_ xsel_2_ XI11_2/XI0/XI0_2/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN0_8 XI11_2/net21_7_ xsel_2_ XI11_2/XI0/XI0_2/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN0_7 XI11_2/net21_8_ xsel_2_ XI11_2/XI0/XI0_2/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN0_6 XI11_2/net21_9_ xsel_2_ XI11_2/XI0/XI0_2/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN0_5 XI11_2/net21_10_ xsel_2_ XI11_2/XI0/XI0_2/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN0_4 XI11_2/net21_11_ xsel_2_ XI11_2/XI0/XI0_2/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN0_3 XI11_2/net21_12_ xsel_2_ XI11_2/XI0/XI0_2/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN0_2 XI11_2/net21_13_ xsel_2_ XI11_2/XI0/XI0_2/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN0_1 XI11_2/net21_14_ xsel_2_ XI11_2/XI0/XI0_2/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN0_0 XI11_2/net21_15_ xsel_2_ XI11_2/XI0/XI0_2/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN1_15 XI11_2/XI0/XI0_2/d__15_ xsel_2_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN1_14 XI11_2/XI0/XI0_2/d__14_ xsel_2_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN1_13 XI11_2/XI0/XI0_2/d__13_ xsel_2_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN1_12 XI11_2/XI0/XI0_2/d__12_ xsel_2_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN1_11 XI11_2/XI0/XI0_2/d__11_ xsel_2_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN1_10 XI11_2/XI0/XI0_2/d__10_ xsel_2_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN1_9 XI11_2/XI0/XI0_2/d__9_ xsel_2_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN1_8 XI11_2/XI0/XI0_2/d__8_ xsel_2_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN1_7 XI11_2/XI0/XI0_2/d__7_ xsel_2_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN1_6 XI11_2/XI0/XI0_2/d__6_ xsel_2_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN1_5 XI11_2/XI0/XI0_2/d__5_ xsel_2_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN1_4 XI11_2/XI0/XI0_2/d__4_ xsel_2_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN1_3 XI11_2/XI0/XI0_2/d__3_ xsel_2_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN1_2 XI11_2/XI0/XI0_2/d__2_ xsel_2_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN1_1 XI11_2/XI0/XI0_2/d__1_ xsel_2_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_2/MN1_0 XI11_2/XI0/XI0_2/d__0_ xsel_2_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN0_15 XI11_2/net21_0_ xsel_1_ XI11_2/XI0/XI0_1/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN0_14 XI11_2/net21_1_ xsel_1_ XI11_2/XI0/XI0_1/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN0_13 XI11_2/net21_2_ xsel_1_ XI11_2/XI0/XI0_1/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN0_12 XI11_2/net21_3_ xsel_1_ XI11_2/XI0/XI0_1/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN0_11 XI11_2/net21_4_ xsel_1_ XI11_2/XI0/XI0_1/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN0_10 XI11_2/net21_5_ xsel_1_ XI11_2/XI0/XI0_1/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN0_9 XI11_2/net21_6_ xsel_1_ XI11_2/XI0/XI0_1/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN0_8 XI11_2/net21_7_ xsel_1_ XI11_2/XI0/XI0_1/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN0_7 XI11_2/net21_8_ xsel_1_ XI11_2/XI0/XI0_1/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN0_6 XI11_2/net21_9_ xsel_1_ XI11_2/XI0/XI0_1/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN0_5 XI11_2/net21_10_ xsel_1_ XI11_2/XI0/XI0_1/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN0_4 XI11_2/net21_11_ xsel_1_ XI11_2/XI0/XI0_1/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN0_3 XI11_2/net21_12_ xsel_1_ XI11_2/XI0/XI0_1/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN0_2 XI11_2/net21_13_ xsel_1_ XI11_2/XI0/XI0_1/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN0_1 XI11_2/net21_14_ xsel_1_ XI11_2/XI0/XI0_1/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN0_0 XI11_2/net21_15_ xsel_1_ XI11_2/XI0/XI0_1/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN1_15 XI11_2/XI0/XI0_1/d__15_ xsel_1_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN1_14 XI11_2/XI0/XI0_1/d__14_ xsel_1_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN1_13 XI11_2/XI0/XI0_1/d__13_ xsel_1_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN1_12 XI11_2/XI0/XI0_1/d__12_ xsel_1_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN1_11 XI11_2/XI0/XI0_1/d__11_ xsel_1_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN1_10 XI11_2/XI0/XI0_1/d__10_ xsel_1_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN1_9 XI11_2/XI0/XI0_1/d__9_ xsel_1_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN1_8 XI11_2/XI0/XI0_1/d__8_ xsel_1_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN1_7 XI11_2/XI0/XI0_1/d__7_ xsel_1_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN1_6 XI11_2/XI0/XI0_1/d__6_ xsel_1_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN1_5 XI11_2/XI0/XI0_1/d__5_ xsel_1_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN1_4 XI11_2/XI0/XI0_1/d__4_ xsel_1_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN1_3 XI11_2/XI0/XI0_1/d__3_ xsel_1_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN1_2 XI11_2/XI0/XI0_1/d__2_ xsel_1_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN1_1 XI11_2/XI0/XI0_1/d__1_ xsel_1_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_1/MN1_0 XI11_2/XI0/XI0_1/d__0_ xsel_1_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN0_15 XI11_2/net21_0_ xsel_0_ XI11_2/XI0/XI0_0/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN0_14 XI11_2/net21_1_ xsel_0_ XI11_2/XI0/XI0_0/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN0_13 XI11_2/net21_2_ xsel_0_ XI11_2/XI0/XI0_0/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN0_12 XI11_2/net21_3_ xsel_0_ XI11_2/XI0/XI0_0/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN0_11 XI11_2/net21_4_ xsel_0_ XI11_2/XI0/XI0_0/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN0_10 XI11_2/net21_5_ xsel_0_ XI11_2/XI0/XI0_0/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN0_9 XI11_2/net21_6_ xsel_0_ XI11_2/XI0/XI0_0/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN0_8 XI11_2/net21_7_ xsel_0_ XI11_2/XI0/XI0_0/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN0_7 XI11_2/net21_8_ xsel_0_ XI11_2/XI0/XI0_0/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN0_6 XI11_2/net21_9_ xsel_0_ XI11_2/XI0/XI0_0/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN0_5 XI11_2/net21_10_ xsel_0_ XI11_2/XI0/XI0_0/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN0_4 XI11_2/net21_11_ xsel_0_ XI11_2/XI0/XI0_0/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN0_3 XI11_2/net21_12_ xsel_0_ XI11_2/XI0/XI0_0/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN0_2 XI11_2/net21_13_ xsel_0_ XI11_2/XI0/XI0_0/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN0_1 XI11_2/net21_14_ xsel_0_ XI11_2/XI0/XI0_0/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN0_0 XI11_2/net21_15_ xsel_0_ XI11_2/XI0/XI0_0/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN1_15 XI11_2/XI0/XI0_0/d__15_ xsel_0_ XI11_2/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN1_14 XI11_2/XI0/XI0_0/d__14_ xsel_0_ XI11_2/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN1_13 XI11_2/XI0/XI0_0/d__13_ xsel_0_ XI11_2/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN1_12 XI11_2/XI0/XI0_0/d__12_ xsel_0_ XI11_2/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN1_11 XI11_2/XI0/XI0_0/d__11_ xsel_0_ XI11_2/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN1_10 XI11_2/XI0/XI0_0/d__10_ xsel_0_ XI11_2/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN1_9 XI11_2/XI0/XI0_0/d__9_ xsel_0_ XI11_2/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN1_8 XI11_2/XI0/XI0_0/d__8_ xsel_0_ XI11_2/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN1_7 XI11_2/XI0/XI0_0/d__7_ xsel_0_ XI11_2/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN1_6 XI11_2/XI0/XI0_0/d__6_ xsel_0_ XI11_2/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN1_5 XI11_2/XI0/XI0_0/d__5_ xsel_0_ XI11_2/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN1_4 XI11_2/XI0/XI0_0/d__4_ xsel_0_ XI11_2/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN1_3 XI11_2/XI0/XI0_0/d__3_ xsel_0_ XI11_2/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN1_2 XI11_2/XI0/XI0_0/d__2_ xsel_0_ XI11_2/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN1_1 XI11_2/XI0/XI0_0/d__1_ xsel_0_ XI11_2/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_2/XI0/XI0_0/MN1_0 XI11_2/XI0/XI0_0/d__0_ xsel_0_ XI11_2/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI2/MN0_15 XI11_1/net21_0_ ysel_15_ XI11_1/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN0_14 XI11_1/net21_1_ ysel_14_ XI11_1/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN0_13 XI11_1/net21_2_ ysel_13_ XI11_1/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN0_12 XI11_1/net21_3_ ysel_12_ XI11_1/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN0_11 XI11_1/net21_4_ ysel_11_ XI11_1/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN0_10 XI11_1/net21_5_ ysel_10_ XI11_1/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN0_9 XI11_1/net21_6_ ysel_9_ XI11_1/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN0_8 XI11_1/net21_7_ ysel_8_ XI11_1/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN0_7 XI11_1/net21_8_ ysel_7_ XI11_1/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN0_6 XI11_1/net21_9_ ysel_6_ XI11_1/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN0_5 XI11_1/net21_10_ ysel_5_ XI11_1/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN0_4 XI11_1/net21_11_ ysel_4_ XI11_1/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN0_3 XI11_1/net21_12_ ysel_3_ XI11_1/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN0_2 XI11_1/net21_13_ ysel_2_ XI11_1/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN0_1 XI11_1/net21_14_ ysel_1_ XI11_1/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN0_0 XI11_1/net21_15_ ysel_0_ XI11_1/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN1_15 XI11_1/net20_0_ ysel_15_ XI11_1/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN1_14 XI11_1/net20_1_ ysel_14_ XI11_1/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN1_13 XI11_1/net20_2_ ysel_13_ XI11_1/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN1_12 XI11_1/net20_3_ ysel_12_ XI11_1/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN1_11 XI11_1/net20_4_ ysel_11_ XI11_1/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN1_10 XI11_1/net20_5_ ysel_10_ XI11_1/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN1_9 XI11_1/net20_6_ ysel_9_ XI11_1/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN1_8 XI11_1/net20_7_ ysel_8_ XI11_1/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN1_7 XI11_1/net20_8_ ysel_7_ XI11_1/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN1_6 XI11_1/net20_9_ ysel_6_ XI11_1/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN1_5 XI11_1/net20_10_ ysel_5_ XI11_1/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN1_4 XI11_1/net20_11_ ysel_4_ XI11_1/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN1_3 XI11_1/net20_12_ ysel_3_ XI11_1/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN1_2 XI11_1/net20_13_ ysel_2_ XI11_1/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN1_1 XI11_1/net20_14_ ysel_1_ XI11_1/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI2/MN1_0 XI11_1/net20_15_ ysel_0_ XI11_1/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_1/XI4/MN8 vdd XI11_1/XI4/net8 XI11_1/net12 vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_1/XI4/MP0 XI11_1/net9 XI11_1/XI4/net23 vdd vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_1/XI4/MP4 XI11_1/net12 XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI4/MP1 XI11_1/net9 XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI4/MP5 XI11_1/net12 XI11_1/preck XI11_1/net9 vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI4/MN7 vdd XI11_1/XI4/net090 DOUT_1_ vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_1/XI4/MP3 gnd XI11_1/XI4/net089 XI11_1/net12 gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_1/XI4/MN5 XI11_1/net9 XI11_1/XI4/net0103 gnd gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_1/XI4/MN4 XI11_1/XI4/data_out_ XI11_1/XI4/net32 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_1/XI4/MN0 XI11_1/XI4/data_out XI11_1/XI4/net52 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_1/XI4/MN9 gnd XI11_1/XI4/net0112 DOUT_1_ gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_1/XI1_15/MP2 XI11_1/net20_0_ XI11_1/preck XI11_1/net21_0_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI1_15/MP1 XI11_1/net20_0_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_15/MP0 XI11_1/net21_0_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_14/MP2 XI11_1/net20_1_ XI11_1/preck XI11_1/net21_1_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI1_14/MP1 XI11_1/net20_1_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_14/MP0 XI11_1/net21_1_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_13/MP2 XI11_1/net20_2_ XI11_1/preck XI11_1/net21_2_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI1_13/MP1 XI11_1/net20_2_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_13/MP0 XI11_1/net21_2_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_12/MP2 XI11_1/net20_3_ XI11_1/preck XI11_1/net21_3_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI1_12/MP1 XI11_1/net20_3_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_12/MP0 XI11_1/net21_3_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_11/MP2 XI11_1/net20_4_ XI11_1/preck XI11_1/net21_4_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI1_11/MP1 XI11_1/net20_4_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_11/MP0 XI11_1/net21_4_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_10/MP2 XI11_1/net20_5_ XI11_1/preck XI11_1/net21_5_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI1_10/MP1 XI11_1/net20_5_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_10/MP0 XI11_1/net21_5_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_9/MP2 XI11_1/net20_6_ XI11_1/preck XI11_1/net21_6_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI1_9/MP1 XI11_1/net20_6_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_9/MP0 XI11_1/net21_6_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_8/MP2 XI11_1/net20_7_ XI11_1/preck XI11_1/net21_7_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI1_8/MP1 XI11_1/net20_7_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_8/MP0 XI11_1/net21_7_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_7/MP2 XI11_1/net20_8_ XI11_1/preck XI11_1/net21_8_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI1_7/MP1 XI11_1/net20_8_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_7/MP0 XI11_1/net21_8_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_6/MP2 XI11_1/net20_9_ XI11_1/preck XI11_1/net21_9_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI1_6/MP1 XI11_1/net20_9_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_6/MP0 XI11_1/net21_9_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_5/MP2 XI11_1/net20_10_ XI11_1/preck XI11_1/net21_10_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI1_5/MP1 XI11_1/net20_10_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_5/MP0 XI11_1/net21_10_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_4/MP2 XI11_1/net20_11_ XI11_1/preck XI11_1/net21_11_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI1_4/MP1 XI11_1/net20_11_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_4/MP0 XI11_1/net21_11_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_3/MP2 XI11_1/net20_12_ XI11_1/preck XI11_1/net21_12_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI1_3/MP1 XI11_1/net20_12_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_3/MP0 XI11_1/net21_12_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_2/MP2 XI11_1/net20_13_ XI11_1/preck XI11_1/net21_13_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI1_2/MP1 XI11_1/net20_13_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_2/MP0 XI11_1/net21_13_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_1/MP2 XI11_1/net20_14_ XI11_1/preck XI11_1/net21_14_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI1_1/MP1 XI11_1/net20_14_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_1/MP0 XI11_1/net21_14_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_0/MP2 XI11_1/net20_15_ XI11_1/preck XI11_1/net21_15_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_1/XI1_0/MP1 XI11_1/net20_15_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI1_0/MP0 XI11_1/net21_15_ XI11_1/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_1/XI0/MN0_15 gnd gnd XI11_1/net21_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN0_14 gnd gnd XI11_1/net21_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN0_13 gnd gnd XI11_1/net21_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN0_12 gnd gnd XI11_1/net21_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN0_11 gnd gnd XI11_1/net21_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN0_10 gnd gnd XI11_1/net21_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN0_9 gnd gnd XI11_1/net21_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN0_8 gnd gnd XI11_1/net21_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN0_7 gnd gnd XI11_1/net21_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN0_6 gnd gnd XI11_1/net21_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN0_5 gnd gnd XI11_1/net21_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN0_4 gnd gnd XI11_1/net21_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN0_3 gnd gnd XI11_1/net21_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN0_2 gnd gnd XI11_1/net21_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN0_1 gnd gnd XI11_1/net21_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN0_0 gnd gnd XI11_1/net21_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN1_15 gnd gnd XI11_1/net20_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN1_14 gnd gnd XI11_1/net20_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN1_13 gnd gnd XI11_1/net20_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN1_12 gnd gnd XI11_1/net20_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN1_11 gnd gnd XI11_1/net20_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN1_10 gnd gnd XI11_1/net20_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN1_9 gnd gnd XI11_1/net20_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN1_8 gnd gnd XI11_1/net20_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN1_7 gnd gnd XI11_1/net20_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN1_6 gnd gnd XI11_1/net20_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN1_5 gnd gnd XI11_1/net20_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN1_4 gnd gnd XI11_1/net20_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN1_3 gnd gnd XI11_1/net20_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN1_2 gnd gnd XI11_1/net20_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN1_1 gnd gnd XI11_1/net20_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/MN1_0 gnd gnd XI11_1/net20_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN0_15 XI11_1/net21_0_ xsel_63_ XI11_1/XI0/XI0_63/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN0_14 XI11_1/net21_1_ xsel_63_ XI11_1/XI0/XI0_63/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN0_13 XI11_1/net21_2_ xsel_63_ XI11_1/XI0/XI0_63/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN0_12 XI11_1/net21_3_ xsel_63_ XI11_1/XI0/XI0_63/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN0_11 XI11_1/net21_4_ xsel_63_ XI11_1/XI0/XI0_63/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN0_10 XI11_1/net21_5_ xsel_63_ XI11_1/XI0/XI0_63/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN0_9 XI11_1/net21_6_ xsel_63_ XI11_1/XI0/XI0_63/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN0_8 XI11_1/net21_7_ xsel_63_ XI11_1/XI0/XI0_63/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN0_7 XI11_1/net21_8_ xsel_63_ XI11_1/XI0/XI0_63/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN0_6 XI11_1/net21_9_ xsel_63_ XI11_1/XI0/XI0_63/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN0_5 XI11_1/net21_10_ xsel_63_ XI11_1/XI0/XI0_63/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN0_4 XI11_1/net21_11_ xsel_63_ XI11_1/XI0/XI0_63/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN0_3 XI11_1/net21_12_ xsel_63_ XI11_1/XI0/XI0_63/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN0_2 XI11_1/net21_13_ xsel_63_ XI11_1/XI0/XI0_63/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN0_1 XI11_1/net21_14_ xsel_63_ XI11_1/XI0/XI0_63/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN0_0 XI11_1/net21_15_ xsel_63_ XI11_1/XI0/XI0_63/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN1_15 XI11_1/XI0/XI0_63/d__15_ xsel_63_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN1_14 XI11_1/XI0/XI0_63/d__14_ xsel_63_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN1_13 XI11_1/XI0/XI0_63/d__13_ xsel_63_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN1_12 XI11_1/XI0/XI0_63/d__12_ xsel_63_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN1_11 XI11_1/XI0/XI0_63/d__11_ xsel_63_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN1_10 XI11_1/XI0/XI0_63/d__10_ xsel_63_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN1_9 XI11_1/XI0/XI0_63/d__9_ xsel_63_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN1_8 XI11_1/XI0/XI0_63/d__8_ xsel_63_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN1_7 XI11_1/XI0/XI0_63/d__7_ xsel_63_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN1_6 XI11_1/XI0/XI0_63/d__6_ xsel_63_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN1_5 XI11_1/XI0/XI0_63/d__5_ xsel_63_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN1_4 XI11_1/XI0/XI0_63/d__4_ xsel_63_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN1_3 XI11_1/XI0/XI0_63/d__3_ xsel_63_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN1_2 XI11_1/XI0/XI0_63/d__2_ xsel_63_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN1_1 XI11_1/XI0/XI0_63/d__1_ xsel_63_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_63/MN1_0 XI11_1/XI0/XI0_63/d__0_ xsel_63_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN0_15 XI11_1/net21_0_ xsel_62_ XI11_1/XI0/XI0_62/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN0_14 XI11_1/net21_1_ xsel_62_ XI11_1/XI0/XI0_62/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN0_13 XI11_1/net21_2_ xsel_62_ XI11_1/XI0/XI0_62/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN0_12 XI11_1/net21_3_ xsel_62_ XI11_1/XI0/XI0_62/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN0_11 XI11_1/net21_4_ xsel_62_ XI11_1/XI0/XI0_62/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN0_10 XI11_1/net21_5_ xsel_62_ XI11_1/XI0/XI0_62/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN0_9 XI11_1/net21_6_ xsel_62_ XI11_1/XI0/XI0_62/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN0_8 XI11_1/net21_7_ xsel_62_ XI11_1/XI0/XI0_62/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN0_7 XI11_1/net21_8_ xsel_62_ XI11_1/XI0/XI0_62/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN0_6 XI11_1/net21_9_ xsel_62_ XI11_1/XI0/XI0_62/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN0_5 XI11_1/net21_10_ xsel_62_ XI11_1/XI0/XI0_62/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN0_4 XI11_1/net21_11_ xsel_62_ XI11_1/XI0/XI0_62/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN0_3 XI11_1/net21_12_ xsel_62_ XI11_1/XI0/XI0_62/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN0_2 XI11_1/net21_13_ xsel_62_ XI11_1/XI0/XI0_62/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN0_1 XI11_1/net21_14_ xsel_62_ XI11_1/XI0/XI0_62/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN0_0 XI11_1/net21_15_ xsel_62_ XI11_1/XI0/XI0_62/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN1_15 XI11_1/XI0/XI0_62/d__15_ xsel_62_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN1_14 XI11_1/XI0/XI0_62/d__14_ xsel_62_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN1_13 XI11_1/XI0/XI0_62/d__13_ xsel_62_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN1_12 XI11_1/XI0/XI0_62/d__12_ xsel_62_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN1_11 XI11_1/XI0/XI0_62/d__11_ xsel_62_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN1_10 XI11_1/XI0/XI0_62/d__10_ xsel_62_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN1_9 XI11_1/XI0/XI0_62/d__9_ xsel_62_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN1_8 XI11_1/XI0/XI0_62/d__8_ xsel_62_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN1_7 XI11_1/XI0/XI0_62/d__7_ xsel_62_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN1_6 XI11_1/XI0/XI0_62/d__6_ xsel_62_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN1_5 XI11_1/XI0/XI0_62/d__5_ xsel_62_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN1_4 XI11_1/XI0/XI0_62/d__4_ xsel_62_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN1_3 XI11_1/XI0/XI0_62/d__3_ xsel_62_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN1_2 XI11_1/XI0/XI0_62/d__2_ xsel_62_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN1_1 XI11_1/XI0/XI0_62/d__1_ xsel_62_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_62/MN1_0 XI11_1/XI0/XI0_62/d__0_ xsel_62_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN0_15 XI11_1/net21_0_ xsel_61_ XI11_1/XI0/XI0_61/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN0_14 XI11_1/net21_1_ xsel_61_ XI11_1/XI0/XI0_61/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN0_13 XI11_1/net21_2_ xsel_61_ XI11_1/XI0/XI0_61/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN0_12 XI11_1/net21_3_ xsel_61_ XI11_1/XI0/XI0_61/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN0_11 XI11_1/net21_4_ xsel_61_ XI11_1/XI0/XI0_61/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN0_10 XI11_1/net21_5_ xsel_61_ XI11_1/XI0/XI0_61/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN0_9 XI11_1/net21_6_ xsel_61_ XI11_1/XI0/XI0_61/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN0_8 XI11_1/net21_7_ xsel_61_ XI11_1/XI0/XI0_61/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN0_7 XI11_1/net21_8_ xsel_61_ XI11_1/XI0/XI0_61/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN0_6 XI11_1/net21_9_ xsel_61_ XI11_1/XI0/XI0_61/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN0_5 XI11_1/net21_10_ xsel_61_ XI11_1/XI0/XI0_61/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN0_4 XI11_1/net21_11_ xsel_61_ XI11_1/XI0/XI0_61/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN0_3 XI11_1/net21_12_ xsel_61_ XI11_1/XI0/XI0_61/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN0_2 XI11_1/net21_13_ xsel_61_ XI11_1/XI0/XI0_61/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN0_1 XI11_1/net21_14_ xsel_61_ XI11_1/XI0/XI0_61/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN0_0 XI11_1/net21_15_ xsel_61_ XI11_1/XI0/XI0_61/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN1_15 XI11_1/XI0/XI0_61/d__15_ xsel_61_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN1_14 XI11_1/XI0/XI0_61/d__14_ xsel_61_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN1_13 XI11_1/XI0/XI0_61/d__13_ xsel_61_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN1_12 XI11_1/XI0/XI0_61/d__12_ xsel_61_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN1_11 XI11_1/XI0/XI0_61/d__11_ xsel_61_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN1_10 XI11_1/XI0/XI0_61/d__10_ xsel_61_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN1_9 XI11_1/XI0/XI0_61/d__9_ xsel_61_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN1_8 XI11_1/XI0/XI0_61/d__8_ xsel_61_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN1_7 XI11_1/XI0/XI0_61/d__7_ xsel_61_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN1_6 XI11_1/XI0/XI0_61/d__6_ xsel_61_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN1_5 XI11_1/XI0/XI0_61/d__5_ xsel_61_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN1_4 XI11_1/XI0/XI0_61/d__4_ xsel_61_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN1_3 XI11_1/XI0/XI0_61/d__3_ xsel_61_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN1_2 XI11_1/XI0/XI0_61/d__2_ xsel_61_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN1_1 XI11_1/XI0/XI0_61/d__1_ xsel_61_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_61/MN1_0 XI11_1/XI0/XI0_61/d__0_ xsel_61_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN0_15 XI11_1/net21_0_ xsel_60_ XI11_1/XI0/XI0_60/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN0_14 XI11_1/net21_1_ xsel_60_ XI11_1/XI0/XI0_60/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN0_13 XI11_1/net21_2_ xsel_60_ XI11_1/XI0/XI0_60/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN0_12 XI11_1/net21_3_ xsel_60_ XI11_1/XI0/XI0_60/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN0_11 XI11_1/net21_4_ xsel_60_ XI11_1/XI0/XI0_60/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN0_10 XI11_1/net21_5_ xsel_60_ XI11_1/XI0/XI0_60/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN0_9 XI11_1/net21_6_ xsel_60_ XI11_1/XI0/XI0_60/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN0_8 XI11_1/net21_7_ xsel_60_ XI11_1/XI0/XI0_60/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN0_7 XI11_1/net21_8_ xsel_60_ XI11_1/XI0/XI0_60/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN0_6 XI11_1/net21_9_ xsel_60_ XI11_1/XI0/XI0_60/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN0_5 XI11_1/net21_10_ xsel_60_ XI11_1/XI0/XI0_60/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN0_4 XI11_1/net21_11_ xsel_60_ XI11_1/XI0/XI0_60/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN0_3 XI11_1/net21_12_ xsel_60_ XI11_1/XI0/XI0_60/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN0_2 XI11_1/net21_13_ xsel_60_ XI11_1/XI0/XI0_60/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN0_1 XI11_1/net21_14_ xsel_60_ XI11_1/XI0/XI0_60/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN0_0 XI11_1/net21_15_ xsel_60_ XI11_1/XI0/XI0_60/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN1_15 XI11_1/XI0/XI0_60/d__15_ xsel_60_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN1_14 XI11_1/XI0/XI0_60/d__14_ xsel_60_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN1_13 XI11_1/XI0/XI0_60/d__13_ xsel_60_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN1_12 XI11_1/XI0/XI0_60/d__12_ xsel_60_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN1_11 XI11_1/XI0/XI0_60/d__11_ xsel_60_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN1_10 XI11_1/XI0/XI0_60/d__10_ xsel_60_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN1_9 XI11_1/XI0/XI0_60/d__9_ xsel_60_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN1_8 XI11_1/XI0/XI0_60/d__8_ xsel_60_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN1_7 XI11_1/XI0/XI0_60/d__7_ xsel_60_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN1_6 XI11_1/XI0/XI0_60/d__6_ xsel_60_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN1_5 XI11_1/XI0/XI0_60/d__5_ xsel_60_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN1_4 XI11_1/XI0/XI0_60/d__4_ xsel_60_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN1_3 XI11_1/XI0/XI0_60/d__3_ xsel_60_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN1_2 XI11_1/XI0/XI0_60/d__2_ xsel_60_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN1_1 XI11_1/XI0/XI0_60/d__1_ xsel_60_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_60/MN1_0 XI11_1/XI0/XI0_60/d__0_ xsel_60_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN0_15 XI11_1/net21_0_ xsel_59_ XI11_1/XI0/XI0_59/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN0_14 XI11_1/net21_1_ xsel_59_ XI11_1/XI0/XI0_59/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN0_13 XI11_1/net21_2_ xsel_59_ XI11_1/XI0/XI0_59/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN0_12 XI11_1/net21_3_ xsel_59_ XI11_1/XI0/XI0_59/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN0_11 XI11_1/net21_4_ xsel_59_ XI11_1/XI0/XI0_59/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN0_10 XI11_1/net21_5_ xsel_59_ XI11_1/XI0/XI0_59/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN0_9 XI11_1/net21_6_ xsel_59_ XI11_1/XI0/XI0_59/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN0_8 XI11_1/net21_7_ xsel_59_ XI11_1/XI0/XI0_59/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN0_7 XI11_1/net21_8_ xsel_59_ XI11_1/XI0/XI0_59/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN0_6 XI11_1/net21_9_ xsel_59_ XI11_1/XI0/XI0_59/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN0_5 XI11_1/net21_10_ xsel_59_ XI11_1/XI0/XI0_59/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN0_4 XI11_1/net21_11_ xsel_59_ XI11_1/XI0/XI0_59/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN0_3 XI11_1/net21_12_ xsel_59_ XI11_1/XI0/XI0_59/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN0_2 XI11_1/net21_13_ xsel_59_ XI11_1/XI0/XI0_59/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN0_1 XI11_1/net21_14_ xsel_59_ XI11_1/XI0/XI0_59/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN0_0 XI11_1/net21_15_ xsel_59_ XI11_1/XI0/XI0_59/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN1_15 XI11_1/XI0/XI0_59/d__15_ xsel_59_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN1_14 XI11_1/XI0/XI0_59/d__14_ xsel_59_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN1_13 XI11_1/XI0/XI0_59/d__13_ xsel_59_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN1_12 XI11_1/XI0/XI0_59/d__12_ xsel_59_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN1_11 XI11_1/XI0/XI0_59/d__11_ xsel_59_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN1_10 XI11_1/XI0/XI0_59/d__10_ xsel_59_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN1_9 XI11_1/XI0/XI0_59/d__9_ xsel_59_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN1_8 XI11_1/XI0/XI0_59/d__8_ xsel_59_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN1_7 XI11_1/XI0/XI0_59/d__7_ xsel_59_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN1_6 XI11_1/XI0/XI0_59/d__6_ xsel_59_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN1_5 XI11_1/XI0/XI0_59/d__5_ xsel_59_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN1_4 XI11_1/XI0/XI0_59/d__4_ xsel_59_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN1_3 XI11_1/XI0/XI0_59/d__3_ xsel_59_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN1_2 XI11_1/XI0/XI0_59/d__2_ xsel_59_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN1_1 XI11_1/XI0/XI0_59/d__1_ xsel_59_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_59/MN1_0 XI11_1/XI0/XI0_59/d__0_ xsel_59_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN0_15 XI11_1/net21_0_ xsel_58_ XI11_1/XI0/XI0_58/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN0_14 XI11_1/net21_1_ xsel_58_ XI11_1/XI0/XI0_58/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN0_13 XI11_1/net21_2_ xsel_58_ XI11_1/XI0/XI0_58/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN0_12 XI11_1/net21_3_ xsel_58_ XI11_1/XI0/XI0_58/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN0_11 XI11_1/net21_4_ xsel_58_ XI11_1/XI0/XI0_58/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN0_10 XI11_1/net21_5_ xsel_58_ XI11_1/XI0/XI0_58/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN0_9 XI11_1/net21_6_ xsel_58_ XI11_1/XI0/XI0_58/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN0_8 XI11_1/net21_7_ xsel_58_ XI11_1/XI0/XI0_58/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN0_7 XI11_1/net21_8_ xsel_58_ XI11_1/XI0/XI0_58/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN0_6 XI11_1/net21_9_ xsel_58_ XI11_1/XI0/XI0_58/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN0_5 XI11_1/net21_10_ xsel_58_ XI11_1/XI0/XI0_58/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN0_4 XI11_1/net21_11_ xsel_58_ XI11_1/XI0/XI0_58/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN0_3 XI11_1/net21_12_ xsel_58_ XI11_1/XI0/XI0_58/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN0_2 XI11_1/net21_13_ xsel_58_ XI11_1/XI0/XI0_58/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN0_1 XI11_1/net21_14_ xsel_58_ XI11_1/XI0/XI0_58/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN0_0 XI11_1/net21_15_ xsel_58_ XI11_1/XI0/XI0_58/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN1_15 XI11_1/XI0/XI0_58/d__15_ xsel_58_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN1_14 XI11_1/XI0/XI0_58/d__14_ xsel_58_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN1_13 XI11_1/XI0/XI0_58/d__13_ xsel_58_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN1_12 XI11_1/XI0/XI0_58/d__12_ xsel_58_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN1_11 XI11_1/XI0/XI0_58/d__11_ xsel_58_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN1_10 XI11_1/XI0/XI0_58/d__10_ xsel_58_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN1_9 XI11_1/XI0/XI0_58/d__9_ xsel_58_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN1_8 XI11_1/XI0/XI0_58/d__8_ xsel_58_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN1_7 XI11_1/XI0/XI0_58/d__7_ xsel_58_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN1_6 XI11_1/XI0/XI0_58/d__6_ xsel_58_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN1_5 XI11_1/XI0/XI0_58/d__5_ xsel_58_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN1_4 XI11_1/XI0/XI0_58/d__4_ xsel_58_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN1_3 XI11_1/XI0/XI0_58/d__3_ xsel_58_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN1_2 XI11_1/XI0/XI0_58/d__2_ xsel_58_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN1_1 XI11_1/XI0/XI0_58/d__1_ xsel_58_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_58/MN1_0 XI11_1/XI0/XI0_58/d__0_ xsel_58_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN0_15 XI11_1/net21_0_ xsel_57_ XI11_1/XI0/XI0_57/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN0_14 XI11_1/net21_1_ xsel_57_ XI11_1/XI0/XI0_57/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN0_13 XI11_1/net21_2_ xsel_57_ XI11_1/XI0/XI0_57/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN0_12 XI11_1/net21_3_ xsel_57_ XI11_1/XI0/XI0_57/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN0_11 XI11_1/net21_4_ xsel_57_ XI11_1/XI0/XI0_57/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN0_10 XI11_1/net21_5_ xsel_57_ XI11_1/XI0/XI0_57/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN0_9 XI11_1/net21_6_ xsel_57_ XI11_1/XI0/XI0_57/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN0_8 XI11_1/net21_7_ xsel_57_ XI11_1/XI0/XI0_57/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN0_7 XI11_1/net21_8_ xsel_57_ XI11_1/XI0/XI0_57/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN0_6 XI11_1/net21_9_ xsel_57_ XI11_1/XI0/XI0_57/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN0_5 XI11_1/net21_10_ xsel_57_ XI11_1/XI0/XI0_57/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN0_4 XI11_1/net21_11_ xsel_57_ XI11_1/XI0/XI0_57/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN0_3 XI11_1/net21_12_ xsel_57_ XI11_1/XI0/XI0_57/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN0_2 XI11_1/net21_13_ xsel_57_ XI11_1/XI0/XI0_57/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN0_1 XI11_1/net21_14_ xsel_57_ XI11_1/XI0/XI0_57/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN0_0 XI11_1/net21_15_ xsel_57_ XI11_1/XI0/XI0_57/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN1_15 XI11_1/XI0/XI0_57/d__15_ xsel_57_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN1_14 XI11_1/XI0/XI0_57/d__14_ xsel_57_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN1_13 XI11_1/XI0/XI0_57/d__13_ xsel_57_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN1_12 XI11_1/XI0/XI0_57/d__12_ xsel_57_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN1_11 XI11_1/XI0/XI0_57/d__11_ xsel_57_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN1_10 XI11_1/XI0/XI0_57/d__10_ xsel_57_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN1_9 XI11_1/XI0/XI0_57/d__9_ xsel_57_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN1_8 XI11_1/XI0/XI0_57/d__8_ xsel_57_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN1_7 XI11_1/XI0/XI0_57/d__7_ xsel_57_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN1_6 XI11_1/XI0/XI0_57/d__6_ xsel_57_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN1_5 XI11_1/XI0/XI0_57/d__5_ xsel_57_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN1_4 XI11_1/XI0/XI0_57/d__4_ xsel_57_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN1_3 XI11_1/XI0/XI0_57/d__3_ xsel_57_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN1_2 XI11_1/XI0/XI0_57/d__2_ xsel_57_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN1_1 XI11_1/XI0/XI0_57/d__1_ xsel_57_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_57/MN1_0 XI11_1/XI0/XI0_57/d__0_ xsel_57_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN0_15 XI11_1/net21_0_ xsel_56_ XI11_1/XI0/XI0_56/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN0_14 XI11_1/net21_1_ xsel_56_ XI11_1/XI0/XI0_56/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN0_13 XI11_1/net21_2_ xsel_56_ XI11_1/XI0/XI0_56/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN0_12 XI11_1/net21_3_ xsel_56_ XI11_1/XI0/XI0_56/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN0_11 XI11_1/net21_4_ xsel_56_ XI11_1/XI0/XI0_56/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN0_10 XI11_1/net21_5_ xsel_56_ XI11_1/XI0/XI0_56/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN0_9 XI11_1/net21_6_ xsel_56_ XI11_1/XI0/XI0_56/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN0_8 XI11_1/net21_7_ xsel_56_ XI11_1/XI0/XI0_56/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN0_7 XI11_1/net21_8_ xsel_56_ XI11_1/XI0/XI0_56/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN0_6 XI11_1/net21_9_ xsel_56_ XI11_1/XI0/XI0_56/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN0_5 XI11_1/net21_10_ xsel_56_ XI11_1/XI0/XI0_56/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN0_4 XI11_1/net21_11_ xsel_56_ XI11_1/XI0/XI0_56/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN0_3 XI11_1/net21_12_ xsel_56_ XI11_1/XI0/XI0_56/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN0_2 XI11_1/net21_13_ xsel_56_ XI11_1/XI0/XI0_56/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN0_1 XI11_1/net21_14_ xsel_56_ XI11_1/XI0/XI0_56/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN0_0 XI11_1/net21_15_ xsel_56_ XI11_1/XI0/XI0_56/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN1_15 XI11_1/XI0/XI0_56/d__15_ xsel_56_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN1_14 XI11_1/XI0/XI0_56/d__14_ xsel_56_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN1_13 XI11_1/XI0/XI0_56/d__13_ xsel_56_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN1_12 XI11_1/XI0/XI0_56/d__12_ xsel_56_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN1_11 XI11_1/XI0/XI0_56/d__11_ xsel_56_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN1_10 XI11_1/XI0/XI0_56/d__10_ xsel_56_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN1_9 XI11_1/XI0/XI0_56/d__9_ xsel_56_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN1_8 XI11_1/XI0/XI0_56/d__8_ xsel_56_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN1_7 XI11_1/XI0/XI0_56/d__7_ xsel_56_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN1_6 XI11_1/XI0/XI0_56/d__6_ xsel_56_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN1_5 XI11_1/XI0/XI0_56/d__5_ xsel_56_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN1_4 XI11_1/XI0/XI0_56/d__4_ xsel_56_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN1_3 XI11_1/XI0/XI0_56/d__3_ xsel_56_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN1_2 XI11_1/XI0/XI0_56/d__2_ xsel_56_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN1_1 XI11_1/XI0/XI0_56/d__1_ xsel_56_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_56/MN1_0 XI11_1/XI0/XI0_56/d__0_ xsel_56_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN0_15 XI11_1/net21_0_ xsel_55_ XI11_1/XI0/XI0_55/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN0_14 XI11_1/net21_1_ xsel_55_ XI11_1/XI0/XI0_55/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN0_13 XI11_1/net21_2_ xsel_55_ XI11_1/XI0/XI0_55/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN0_12 XI11_1/net21_3_ xsel_55_ XI11_1/XI0/XI0_55/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN0_11 XI11_1/net21_4_ xsel_55_ XI11_1/XI0/XI0_55/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN0_10 XI11_1/net21_5_ xsel_55_ XI11_1/XI0/XI0_55/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN0_9 XI11_1/net21_6_ xsel_55_ XI11_1/XI0/XI0_55/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN0_8 XI11_1/net21_7_ xsel_55_ XI11_1/XI0/XI0_55/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN0_7 XI11_1/net21_8_ xsel_55_ XI11_1/XI0/XI0_55/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN0_6 XI11_1/net21_9_ xsel_55_ XI11_1/XI0/XI0_55/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN0_5 XI11_1/net21_10_ xsel_55_ XI11_1/XI0/XI0_55/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN0_4 XI11_1/net21_11_ xsel_55_ XI11_1/XI0/XI0_55/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN0_3 XI11_1/net21_12_ xsel_55_ XI11_1/XI0/XI0_55/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN0_2 XI11_1/net21_13_ xsel_55_ XI11_1/XI0/XI0_55/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN0_1 XI11_1/net21_14_ xsel_55_ XI11_1/XI0/XI0_55/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN0_0 XI11_1/net21_15_ xsel_55_ XI11_1/XI0/XI0_55/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN1_15 XI11_1/XI0/XI0_55/d__15_ xsel_55_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN1_14 XI11_1/XI0/XI0_55/d__14_ xsel_55_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN1_13 XI11_1/XI0/XI0_55/d__13_ xsel_55_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN1_12 XI11_1/XI0/XI0_55/d__12_ xsel_55_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN1_11 XI11_1/XI0/XI0_55/d__11_ xsel_55_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN1_10 XI11_1/XI0/XI0_55/d__10_ xsel_55_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN1_9 XI11_1/XI0/XI0_55/d__9_ xsel_55_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN1_8 XI11_1/XI0/XI0_55/d__8_ xsel_55_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN1_7 XI11_1/XI0/XI0_55/d__7_ xsel_55_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN1_6 XI11_1/XI0/XI0_55/d__6_ xsel_55_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN1_5 XI11_1/XI0/XI0_55/d__5_ xsel_55_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN1_4 XI11_1/XI0/XI0_55/d__4_ xsel_55_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN1_3 XI11_1/XI0/XI0_55/d__3_ xsel_55_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN1_2 XI11_1/XI0/XI0_55/d__2_ xsel_55_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN1_1 XI11_1/XI0/XI0_55/d__1_ xsel_55_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_55/MN1_0 XI11_1/XI0/XI0_55/d__0_ xsel_55_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN0_15 XI11_1/net21_0_ xsel_54_ XI11_1/XI0/XI0_54/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN0_14 XI11_1/net21_1_ xsel_54_ XI11_1/XI0/XI0_54/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN0_13 XI11_1/net21_2_ xsel_54_ XI11_1/XI0/XI0_54/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN0_12 XI11_1/net21_3_ xsel_54_ XI11_1/XI0/XI0_54/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN0_11 XI11_1/net21_4_ xsel_54_ XI11_1/XI0/XI0_54/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN0_10 XI11_1/net21_5_ xsel_54_ XI11_1/XI0/XI0_54/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN0_9 XI11_1/net21_6_ xsel_54_ XI11_1/XI0/XI0_54/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN0_8 XI11_1/net21_7_ xsel_54_ XI11_1/XI0/XI0_54/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN0_7 XI11_1/net21_8_ xsel_54_ XI11_1/XI0/XI0_54/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN0_6 XI11_1/net21_9_ xsel_54_ XI11_1/XI0/XI0_54/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN0_5 XI11_1/net21_10_ xsel_54_ XI11_1/XI0/XI0_54/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN0_4 XI11_1/net21_11_ xsel_54_ XI11_1/XI0/XI0_54/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN0_3 XI11_1/net21_12_ xsel_54_ XI11_1/XI0/XI0_54/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN0_2 XI11_1/net21_13_ xsel_54_ XI11_1/XI0/XI0_54/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN0_1 XI11_1/net21_14_ xsel_54_ XI11_1/XI0/XI0_54/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN0_0 XI11_1/net21_15_ xsel_54_ XI11_1/XI0/XI0_54/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN1_15 XI11_1/XI0/XI0_54/d__15_ xsel_54_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN1_14 XI11_1/XI0/XI0_54/d__14_ xsel_54_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN1_13 XI11_1/XI0/XI0_54/d__13_ xsel_54_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN1_12 XI11_1/XI0/XI0_54/d__12_ xsel_54_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN1_11 XI11_1/XI0/XI0_54/d__11_ xsel_54_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN1_10 XI11_1/XI0/XI0_54/d__10_ xsel_54_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN1_9 XI11_1/XI0/XI0_54/d__9_ xsel_54_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN1_8 XI11_1/XI0/XI0_54/d__8_ xsel_54_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN1_7 XI11_1/XI0/XI0_54/d__7_ xsel_54_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN1_6 XI11_1/XI0/XI0_54/d__6_ xsel_54_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN1_5 XI11_1/XI0/XI0_54/d__5_ xsel_54_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN1_4 XI11_1/XI0/XI0_54/d__4_ xsel_54_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN1_3 XI11_1/XI0/XI0_54/d__3_ xsel_54_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN1_2 XI11_1/XI0/XI0_54/d__2_ xsel_54_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN1_1 XI11_1/XI0/XI0_54/d__1_ xsel_54_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_54/MN1_0 XI11_1/XI0/XI0_54/d__0_ xsel_54_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN0_15 XI11_1/net21_0_ xsel_53_ XI11_1/XI0/XI0_53/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN0_14 XI11_1/net21_1_ xsel_53_ XI11_1/XI0/XI0_53/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN0_13 XI11_1/net21_2_ xsel_53_ XI11_1/XI0/XI0_53/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN0_12 XI11_1/net21_3_ xsel_53_ XI11_1/XI0/XI0_53/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN0_11 XI11_1/net21_4_ xsel_53_ XI11_1/XI0/XI0_53/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN0_10 XI11_1/net21_5_ xsel_53_ XI11_1/XI0/XI0_53/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN0_9 XI11_1/net21_6_ xsel_53_ XI11_1/XI0/XI0_53/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN0_8 XI11_1/net21_7_ xsel_53_ XI11_1/XI0/XI0_53/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN0_7 XI11_1/net21_8_ xsel_53_ XI11_1/XI0/XI0_53/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN0_6 XI11_1/net21_9_ xsel_53_ XI11_1/XI0/XI0_53/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN0_5 XI11_1/net21_10_ xsel_53_ XI11_1/XI0/XI0_53/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN0_4 XI11_1/net21_11_ xsel_53_ XI11_1/XI0/XI0_53/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN0_3 XI11_1/net21_12_ xsel_53_ XI11_1/XI0/XI0_53/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN0_2 XI11_1/net21_13_ xsel_53_ XI11_1/XI0/XI0_53/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN0_1 XI11_1/net21_14_ xsel_53_ XI11_1/XI0/XI0_53/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN0_0 XI11_1/net21_15_ xsel_53_ XI11_1/XI0/XI0_53/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN1_15 XI11_1/XI0/XI0_53/d__15_ xsel_53_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN1_14 XI11_1/XI0/XI0_53/d__14_ xsel_53_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN1_13 XI11_1/XI0/XI0_53/d__13_ xsel_53_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN1_12 XI11_1/XI0/XI0_53/d__12_ xsel_53_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN1_11 XI11_1/XI0/XI0_53/d__11_ xsel_53_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN1_10 XI11_1/XI0/XI0_53/d__10_ xsel_53_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN1_9 XI11_1/XI0/XI0_53/d__9_ xsel_53_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN1_8 XI11_1/XI0/XI0_53/d__8_ xsel_53_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN1_7 XI11_1/XI0/XI0_53/d__7_ xsel_53_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN1_6 XI11_1/XI0/XI0_53/d__6_ xsel_53_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN1_5 XI11_1/XI0/XI0_53/d__5_ xsel_53_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN1_4 XI11_1/XI0/XI0_53/d__4_ xsel_53_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN1_3 XI11_1/XI0/XI0_53/d__3_ xsel_53_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN1_2 XI11_1/XI0/XI0_53/d__2_ xsel_53_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN1_1 XI11_1/XI0/XI0_53/d__1_ xsel_53_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_53/MN1_0 XI11_1/XI0/XI0_53/d__0_ xsel_53_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN0_15 XI11_1/net21_0_ xsel_52_ XI11_1/XI0/XI0_52/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN0_14 XI11_1/net21_1_ xsel_52_ XI11_1/XI0/XI0_52/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN0_13 XI11_1/net21_2_ xsel_52_ XI11_1/XI0/XI0_52/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN0_12 XI11_1/net21_3_ xsel_52_ XI11_1/XI0/XI0_52/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN0_11 XI11_1/net21_4_ xsel_52_ XI11_1/XI0/XI0_52/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN0_10 XI11_1/net21_5_ xsel_52_ XI11_1/XI0/XI0_52/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN0_9 XI11_1/net21_6_ xsel_52_ XI11_1/XI0/XI0_52/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN0_8 XI11_1/net21_7_ xsel_52_ XI11_1/XI0/XI0_52/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN0_7 XI11_1/net21_8_ xsel_52_ XI11_1/XI0/XI0_52/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN0_6 XI11_1/net21_9_ xsel_52_ XI11_1/XI0/XI0_52/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN0_5 XI11_1/net21_10_ xsel_52_ XI11_1/XI0/XI0_52/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN0_4 XI11_1/net21_11_ xsel_52_ XI11_1/XI0/XI0_52/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN0_3 XI11_1/net21_12_ xsel_52_ XI11_1/XI0/XI0_52/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN0_2 XI11_1/net21_13_ xsel_52_ XI11_1/XI0/XI0_52/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN0_1 XI11_1/net21_14_ xsel_52_ XI11_1/XI0/XI0_52/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN0_0 XI11_1/net21_15_ xsel_52_ XI11_1/XI0/XI0_52/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN1_15 XI11_1/XI0/XI0_52/d__15_ xsel_52_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN1_14 XI11_1/XI0/XI0_52/d__14_ xsel_52_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN1_13 XI11_1/XI0/XI0_52/d__13_ xsel_52_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN1_12 XI11_1/XI0/XI0_52/d__12_ xsel_52_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN1_11 XI11_1/XI0/XI0_52/d__11_ xsel_52_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN1_10 XI11_1/XI0/XI0_52/d__10_ xsel_52_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN1_9 XI11_1/XI0/XI0_52/d__9_ xsel_52_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN1_8 XI11_1/XI0/XI0_52/d__8_ xsel_52_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN1_7 XI11_1/XI0/XI0_52/d__7_ xsel_52_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN1_6 XI11_1/XI0/XI0_52/d__6_ xsel_52_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN1_5 XI11_1/XI0/XI0_52/d__5_ xsel_52_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN1_4 XI11_1/XI0/XI0_52/d__4_ xsel_52_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN1_3 XI11_1/XI0/XI0_52/d__3_ xsel_52_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN1_2 XI11_1/XI0/XI0_52/d__2_ xsel_52_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN1_1 XI11_1/XI0/XI0_52/d__1_ xsel_52_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_52/MN1_0 XI11_1/XI0/XI0_52/d__0_ xsel_52_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN0_15 XI11_1/net21_0_ xsel_51_ XI11_1/XI0/XI0_51/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN0_14 XI11_1/net21_1_ xsel_51_ XI11_1/XI0/XI0_51/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN0_13 XI11_1/net21_2_ xsel_51_ XI11_1/XI0/XI0_51/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN0_12 XI11_1/net21_3_ xsel_51_ XI11_1/XI0/XI0_51/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN0_11 XI11_1/net21_4_ xsel_51_ XI11_1/XI0/XI0_51/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN0_10 XI11_1/net21_5_ xsel_51_ XI11_1/XI0/XI0_51/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN0_9 XI11_1/net21_6_ xsel_51_ XI11_1/XI0/XI0_51/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN0_8 XI11_1/net21_7_ xsel_51_ XI11_1/XI0/XI0_51/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN0_7 XI11_1/net21_8_ xsel_51_ XI11_1/XI0/XI0_51/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN0_6 XI11_1/net21_9_ xsel_51_ XI11_1/XI0/XI0_51/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN0_5 XI11_1/net21_10_ xsel_51_ XI11_1/XI0/XI0_51/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN0_4 XI11_1/net21_11_ xsel_51_ XI11_1/XI0/XI0_51/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN0_3 XI11_1/net21_12_ xsel_51_ XI11_1/XI0/XI0_51/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN0_2 XI11_1/net21_13_ xsel_51_ XI11_1/XI0/XI0_51/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN0_1 XI11_1/net21_14_ xsel_51_ XI11_1/XI0/XI0_51/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN0_0 XI11_1/net21_15_ xsel_51_ XI11_1/XI0/XI0_51/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN1_15 XI11_1/XI0/XI0_51/d__15_ xsel_51_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN1_14 XI11_1/XI0/XI0_51/d__14_ xsel_51_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN1_13 XI11_1/XI0/XI0_51/d__13_ xsel_51_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN1_12 XI11_1/XI0/XI0_51/d__12_ xsel_51_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN1_11 XI11_1/XI0/XI0_51/d__11_ xsel_51_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN1_10 XI11_1/XI0/XI0_51/d__10_ xsel_51_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN1_9 XI11_1/XI0/XI0_51/d__9_ xsel_51_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN1_8 XI11_1/XI0/XI0_51/d__8_ xsel_51_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN1_7 XI11_1/XI0/XI0_51/d__7_ xsel_51_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN1_6 XI11_1/XI0/XI0_51/d__6_ xsel_51_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN1_5 XI11_1/XI0/XI0_51/d__5_ xsel_51_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN1_4 XI11_1/XI0/XI0_51/d__4_ xsel_51_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN1_3 XI11_1/XI0/XI0_51/d__3_ xsel_51_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN1_2 XI11_1/XI0/XI0_51/d__2_ xsel_51_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN1_1 XI11_1/XI0/XI0_51/d__1_ xsel_51_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_51/MN1_0 XI11_1/XI0/XI0_51/d__0_ xsel_51_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN0_15 XI11_1/net21_0_ xsel_50_ XI11_1/XI0/XI0_50/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN0_14 XI11_1/net21_1_ xsel_50_ XI11_1/XI0/XI0_50/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN0_13 XI11_1/net21_2_ xsel_50_ XI11_1/XI0/XI0_50/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN0_12 XI11_1/net21_3_ xsel_50_ XI11_1/XI0/XI0_50/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN0_11 XI11_1/net21_4_ xsel_50_ XI11_1/XI0/XI0_50/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN0_10 XI11_1/net21_5_ xsel_50_ XI11_1/XI0/XI0_50/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN0_9 XI11_1/net21_6_ xsel_50_ XI11_1/XI0/XI0_50/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN0_8 XI11_1/net21_7_ xsel_50_ XI11_1/XI0/XI0_50/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN0_7 XI11_1/net21_8_ xsel_50_ XI11_1/XI0/XI0_50/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN0_6 XI11_1/net21_9_ xsel_50_ XI11_1/XI0/XI0_50/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN0_5 XI11_1/net21_10_ xsel_50_ XI11_1/XI0/XI0_50/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN0_4 XI11_1/net21_11_ xsel_50_ XI11_1/XI0/XI0_50/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN0_3 XI11_1/net21_12_ xsel_50_ XI11_1/XI0/XI0_50/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN0_2 XI11_1/net21_13_ xsel_50_ XI11_1/XI0/XI0_50/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN0_1 XI11_1/net21_14_ xsel_50_ XI11_1/XI0/XI0_50/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN0_0 XI11_1/net21_15_ xsel_50_ XI11_1/XI0/XI0_50/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN1_15 XI11_1/XI0/XI0_50/d__15_ xsel_50_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN1_14 XI11_1/XI0/XI0_50/d__14_ xsel_50_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN1_13 XI11_1/XI0/XI0_50/d__13_ xsel_50_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN1_12 XI11_1/XI0/XI0_50/d__12_ xsel_50_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN1_11 XI11_1/XI0/XI0_50/d__11_ xsel_50_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN1_10 XI11_1/XI0/XI0_50/d__10_ xsel_50_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN1_9 XI11_1/XI0/XI0_50/d__9_ xsel_50_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN1_8 XI11_1/XI0/XI0_50/d__8_ xsel_50_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN1_7 XI11_1/XI0/XI0_50/d__7_ xsel_50_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN1_6 XI11_1/XI0/XI0_50/d__6_ xsel_50_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN1_5 XI11_1/XI0/XI0_50/d__5_ xsel_50_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN1_4 XI11_1/XI0/XI0_50/d__4_ xsel_50_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN1_3 XI11_1/XI0/XI0_50/d__3_ xsel_50_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN1_2 XI11_1/XI0/XI0_50/d__2_ xsel_50_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN1_1 XI11_1/XI0/XI0_50/d__1_ xsel_50_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_50/MN1_0 XI11_1/XI0/XI0_50/d__0_ xsel_50_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN0_15 XI11_1/net21_0_ xsel_49_ XI11_1/XI0/XI0_49/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN0_14 XI11_1/net21_1_ xsel_49_ XI11_1/XI0/XI0_49/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN0_13 XI11_1/net21_2_ xsel_49_ XI11_1/XI0/XI0_49/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN0_12 XI11_1/net21_3_ xsel_49_ XI11_1/XI0/XI0_49/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN0_11 XI11_1/net21_4_ xsel_49_ XI11_1/XI0/XI0_49/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN0_10 XI11_1/net21_5_ xsel_49_ XI11_1/XI0/XI0_49/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN0_9 XI11_1/net21_6_ xsel_49_ XI11_1/XI0/XI0_49/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN0_8 XI11_1/net21_7_ xsel_49_ XI11_1/XI0/XI0_49/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN0_7 XI11_1/net21_8_ xsel_49_ XI11_1/XI0/XI0_49/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN0_6 XI11_1/net21_9_ xsel_49_ XI11_1/XI0/XI0_49/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN0_5 XI11_1/net21_10_ xsel_49_ XI11_1/XI0/XI0_49/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN0_4 XI11_1/net21_11_ xsel_49_ XI11_1/XI0/XI0_49/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN0_3 XI11_1/net21_12_ xsel_49_ XI11_1/XI0/XI0_49/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN0_2 XI11_1/net21_13_ xsel_49_ XI11_1/XI0/XI0_49/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN0_1 XI11_1/net21_14_ xsel_49_ XI11_1/XI0/XI0_49/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN0_0 XI11_1/net21_15_ xsel_49_ XI11_1/XI0/XI0_49/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN1_15 XI11_1/XI0/XI0_49/d__15_ xsel_49_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN1_14 XI11_1/XI0/XI0_49/d__14_ xsel_49_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN1_13 XI11_1/XI0/XI0_49/d__13_ xsel_49_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN1_12 XI11_1/XI0/XI0_49/d__12_ xsel_49_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN1_11 XI11_1/XI0/XI0_49/d__11_ xsel_49_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN1_10 XI11_1/XI0/XI0_49/d__10_ xsel_49_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN1_9 XI11_1/XI0/XI0_49/d__9_ xsel_49_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN1_8 XI11_1/XI0/XI0_49/d__8_ xsel_49_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN1_7 XI11_1/XI0/XI0_49/d__7_ xsel_49_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN1_6 XI11_1/XI0/XI0_49/d__6_ xsel_49_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN1_5 XI11_1/XI0/XI0_49/d__5_ xsel_49_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN1_4 XI11_1/XI0/XI0_49/d__4_ xsel_49_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN1_3 XI11_1/XI0/XI0_49/d__3_ xsel_49_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN1_2 XI11_1/XI0/XI0_49/d__2_ xsel_49_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN1_1 XI11_1/XI0/XI0_49/d__1_ xsel_49_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_49/MN1_0 XI11_1/XI0/XI0_49/d__0_ xsel_49_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN0_15 XI11_1/net21_0_ xsel_48_ XI11_1/XI0/XI0_48/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN0_14 XI11_1/net21_1_ xsel_48_ XI11_1/XI0/XI0_48/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN0_13 XI11_1/net21_2_ xsel_48_ XI11_1/XI0/XI0_48/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN0_12 XI11_1/net21_3_ xsel_48_ XI11_1/XI0/XI0_48/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN0_11 XI11_1/net21_4_ xsel_48_ XI11_1/XI0/XI0_48/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN0_10 XI11_1/net21_5_ xsel_48_ XI11_1/XI0/XI0_48/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN0_9 XI11_1/net21_6_ xsel_48_ XI11_1/XI0/XI0_48/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN0_8 XI11_1/net21_7_ xsel_48_ XI11_1/XI0/XI0_48/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN0_7 XI11_1/net21_8_ xsel_48_ XI11_1/XI0/XI0_48/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN0_6 XI11_1/net21_9_ xsel_48_ XI11_1/XI0/XI0_48/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN0_5 XI11_1/net21_10_ xsel_48_ XI11_1/XI0/XI0_48/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN0_4 XI11_1/net21_11_ xsel_48_ XI11_1/XI0/XI0_48/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN0_3 XI11_1/net21_12_ xsel_48_ XI11_1/XI0/XI0_48/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN0_2 XI11_1/net21_13_ xsel_48_ XI11_1/XI0/XI0_48/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN0_1 XI11_1/net21_14_ xsel_48_ XI11_1/XI0/XI0_48/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN0_0 XI11_1/net21_15_ xsel_48_ XI11_1/XI0/XI0_48/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN1_15 XI11_1/XI0/XI0_48/d__15_ xsel_48_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN1_14 XI11_1/XI0/XI0_48/d__14_ xsel_48_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN1_13 XI11_1/XI0/XI0_48/d__13_ xsel_48_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN1_12 XI11_1/XI0/XI0_48/d__12_ xsel_48_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN1_11 XI11_1/XI0/XI0_48/d__11_ xsel_48_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN1_10 XI11_1/XI0/XI0_48/d__10_ xsel_48_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN1_9 XI11_1/XI0/XI0_48/d__9_ xsel_48_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN1_8 XI11_1/XI0/XI0_48/d__8_ xsel_48_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN1_7 XI11_1/XI0/XI0_48/d__7_ xsel_48_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN1_6 XI11_1/XI0/XI0_48/d__6_ xsel_48_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN1_5 XI11_1/XI0/XI0_48/d__5_ xsel_48_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN1_4 XI11_1/XI0/XI0_48/d__4_ xsel_48_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN1_3 XI11_1/XI0/XI0_48/d__3_ xsel_48_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN1_2 XI11_1/XI0/XI0_48/d__2_ xsel_48_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN1_1 XI11_1/XI0/XI0_48/d__1_ xsel_48_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_48/MN1_0 XI11_1/XI0/XI0_48/d__0_ xsel_48_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN0_15 XI11_1/net21_0_ xsel_47_ XI11_1/XI0/XI0_47/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN0_14 XI11_1/net21_1_ xsel_47_ XI11_1/XI0/XI0_47/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN0_13 XI11_1/net21_2_ xsel_47_ XI11_1/XI0/XI0_47/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN0_12 XI11_1/net21_3_ xsel_47_ XI11_1/XI0/XI0_47/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN0_11 XI11_1/net21_4_ xsel_47_ XI11_1/XI0/XI0_47/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN0_10 XI11_1/net21_5_ xsel_47_ XI11_1/XI0/XI0_47/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN0_9 XI11_1/net21_6_ xsel_47_ XI11_1/XI0/XI0_47/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN0_8 XI11_1/net21_7_ xsel_47_ XI11_1/XI0/XI0_47/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN0_7 XI11_1/net21_8_ xsel_47_ XI11_1/XI0/XI0_47/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN0_6 XI11_1/net21_9_ xsel_47_ XI11_1/XI0/XI0_47/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN0_5 XI11_1/net21_10_ xsel_47_ XI11_1/XI0/XI0_47/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN0_4 XI11_1/net21_11_ xsel_47_ XI11_1/XI0/XI0_47/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN0_3 XI11_1/net21_12_ xsel_47_ XI11_1/XI0/XI0_47/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN0_2 XI11_1/net21_13_ xsel_47_ XI11_1/XI0/XI0_47/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN0_1 XI11_1/net21_14_ xsel_47_ XI11_1/XI0/XI0_47/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN0_0 XI11_1/net21_15_ xsel_47_ XI11_1/XI0/XI0_47/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN1_15 XI11_1/XI0/XI0_47/d__15_ xsel_47_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN1_14 XI11_1/XI0/XI0_47/d__14_ xsel_47_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN1_13 XI11_1/XI0/XI0_47/d__13_ xsel_47_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN1_12 XI11_1/XI0/XI0_47/d__12_ xsel_47_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN1_11 XI11_1/XI0/XI0_47/d__11_ xsel_47_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN1_10 XI11_1/XI0/XI0_47/d__10_ xsel_47_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN1_9 XI11_1/XI0/XI0_47/d__9_ xsel_47_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN1_8 XI11_1/XI0/XI0_47/d__8_ xsel_47_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN1_7 XI11_1/XI0/XI0_47/d__7_ xsel_47_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN1_6 XI11_1/XI0/XI0_47/d__6_ xsel_47_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN1_5 XI11_1/XI0/XI0_47/d__5_ xsel_47_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN1_4 XI11_1/XI0/XI0_47/d__4_ xsel_47_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN1_3 XI11_1/XI0/XI0_47/d__3_ xsel_47_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN1_2 XI11_1/XI0/XI0_47/d__2_ xsel_47_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN1_1 XI11_1/XI0/XI0_47/d__1_ xsel_47_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_47/MN1_0 XI11_1/XI0/XI0_47/d__0_ xsel_47_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN0_15 XI11_1/net21_0_ xsel_46_ XI11_1/XI0/XI0_46/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN0_14 XI11_1/net21_1_ xsel_46_ XI11_1/XI0/XI0_46/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN0_13 XI11_1/net21_2_ xsel_46_ XI11_1/XI0/XI0_46/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN0_12 XI11_1/net21_3_ xsel_46_ XI11_1/XI0/XI0_46/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN0_11 XI11_1/net21_4_ xsel_46_ XI11_1/XI0/XI0_46/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN0_10 XI11_1/net21_5_ xsel_46_ XI11_1/XI0/XI0_46/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN0_9 XI11_1/net21_6_ xsel_46_ XI11_1/XI0/XI0_46/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN0_8 XI11_1/net21_7_ xsel_46_ XI11_1/XI0/XI0_46/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN0_7 XI11_1/net21_8_ xsel_46_ XI11_1/XI0/XI0_46/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN0_6 XI11_1/net21_9_ xsel_46_ XI11_1/XI0/XI0_46/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN0_5 XI11_1/net21_10_ xsel_46_ XI11_1/XI0/XI0_46/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN0_4 XI11_1/net21_11_ xsel_46_ XI11_1/XI0/XI0_46/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN0_3 XI11_1/net21_12_ xsel_46_ XI11_1/XI0/XI0_46/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN0_2 XI11_1/net21_13_ xsel_46_ XI11_1/XI0/XI0_46/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN0_1 XI11_1/net21_14_ xsel_46_ XI11_1/XI0/XI0_46/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN0_0 XI11_1/net21_15_ xsel_46_ XI11_1/XI0/XI0_46/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN1_15 XI11_1/XI0/XI0_46/d__15_ xsel_46_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN1_14 XI11_1/XI0/XI0_46/d__14_ xsel_46_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN1_13 XI11_1/XI0/XI0_46/d__13_ xsel_46_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN1_12 XI11_1/XI0/XI0_46/d__12_ xsel_46_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN1_11 XI11_1/XI0/XI0_46/d__11_ xsel_46_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN1_10 XI11_1/XI0/XI0_46/d__10_ xsel_46_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN1_9 XI11_1/XI0/XI0_46/d__9_ xsel_46_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN1_8 XI11_1/XI0/XI0_46/d__8_ xsel_46_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN1_7 XI11_1/XI0/XI0_46/d__7_ xsel_46_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN1_6 XI11_1/XI0/XI0_46/d__6_ xsel_46_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN1_5 XI11_1/XI0/XI0_46/d__5_ xsel_46_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN1_4 XI11_1/XI0/XI0_46/d__4_ xsel_46_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN1_3 XI11_1/XI0/XI0_46/d__3_ xsel_46_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN1_2 XI11_1/XI0/XI0_46/d__2_ xsel_46_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN1_1 XI11_1/XI0/XI0_46/d__1_ xsel_46_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_46/MN1_0 XI11_1/XI0/XI0_46/d__0_ xsel_46_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN0_15 XI11_1/net21_0_ xsel_45_ XI11_1/XI0/XI0_45/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN0_14 XI11_1/net21_1_ xsel_45_ XI11_1/XI0/XI0_45/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN0_13 XI11_1/net21_2_ xsel_45_ XI11_1/XI0/XI0_45/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN0_12 XI11_1/net21_3_ xsel_45_ XI11_1/XI0/XI0_45/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN0_11 XI11_1/net21_4_ xsel_45_ XI11_1/XI0/XI0_45/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN0_10 XI11_1/net21_5_ xsel_45_ XI11_1/XI0/XI0_45/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN0_9 XI11_1/net21_6_ xsel_45_ XI11_1/XI0/XI0_45/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN0_8 XI11_1/net21_7_ xsel_45_ XI11_1/XI0/XI0_45/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN0_7 XI11_1/net21_8_ xsel_45_ XI11_1/XI0/XI0_45/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN0_6 XI11_1/net21_9_ xsel_45_ XI11_1/XI0/XI0_45/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN0_5 XI11_1/net21_10_ xsel_45_ XI11_1/XI0/XI0_45/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN0_4 XI11_1/net21_11_ xsel_45_ XI11_1/XI0/XI0_45/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN0_3 XI11_1/net21_12_ xsel_45_ XI11_1/XI0/XI0_45/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN0_2 XI11_1/net21_13_ xsel_45_ XI11_1/XI0/XI0_45/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN0_1 XI11_1/net21_14_ xsel_45_ XI11_1/XI0/XI0_45/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN0_0 XI11_1/net21_15_ xsel_45_ XI11_1/XI0/XI0_45/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN1_15 XI11_1/XI0/XI0_45/d__15_ xsel_45_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN1_14 XI11_1/XI0/XI0_45/d__14_ xsel_45_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN1_13 XI11_1/XI0/XI0_45/d__13_ xsel_45_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN1_12 XI11_1/XI0/XI0_45/d__12_ xsel_45_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN1_11 XI11_1/XI0/XI0_45/d__11_ xsel_45_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN1_10 XI11_1/XI0/XI0_45/d__10_ xsel_45_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN1_9 XI11_1/XI0/XI0_45/d__9_ xsel_45_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN1_8 XI11_1/XI0/XI0_45/d__8_ xsel_45_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN1_7 XI11_1/XI0/XI0_45/d__7_ xsel_45_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN1_6 XI11_1/XI0/XI0_45/d__6_ xsel_45_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN1_5 XI11_1/XI0/XI0_45/d__5_ xsel_45_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN1_4 XI11_1/XI0/XI0_45/d__4_ xsel_45_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN1_3 XI11_1/XI0/XI0_45/d__3_ xsel_45_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN1_2 XI11_1/XI0/XI0_45/d__2_ xsel_45_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN1_1 XI11_1/XI0/XI0_45/d__1_ xsel_45_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_45/MN1_0 XI11_1/XI0/XI0_45/d__0_ xsel_45_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN0_15 XI11_1/net21_0_ xsel_44_ XI11_1/XI0/XI0_44/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN0_14 XI11_1/net21_1_ xsel_44_ XI11_1/XI0/XI0_44/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN0_13 XI11_1/net21_2_ xsel_44_ XI11_1/XI0/XI0_44/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN0_12 XI11_1/net21_3_ xsel_44_ XI11_1/XI0/XI0_44/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN0_11 XI11_1/net21_4_ xsel_44_ XI11_1/XI0/XI0_44/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN0_10 XI11_1/net21_5_ xsel_44_ XI11_1/XI0/XI0_44/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN0_9 XI11_1/net21_6_ xsel_44_ XI11_1/XI0/XI0_44/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN0_8 XI11_1/net21_7_ xsel_44_ XI11_1/XI0/XI0_44/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN0_7 XI11_1/net21_8_ xsel_44_ XI11_1/XI0/XI0_44/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN0_6 XI11_1/net21_9_ xsel_44_ XI11_1/XI0/XI0_44/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN0_5 XI11_1/net21_10_ xsel_44_ XI11_1/XI0/XI0_44/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN0_4 XI11_1/net21_11_ xsel_44_ XI11_1/XI0/XI0_44/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN0_3 XI11_1/net21_12_ xsel_44_ XI11_1/XI0/XI0_44/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN0_2 XI11_1/net21_13_ xsel_44_ XI11_1/XI0/XI0_44/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN0_1 XI11_1/net21_14_ xsel_44_ XI11_1/XI0/XI0_44/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN0_0 XI11_1/net21_15_ xsel_44_ XI11_1/XI0/XI0_44/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN1_15 XI11_1/XI0/XI0_44/d__15_ xsel_44_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN1_14 XI11_1/XI0/XI0_44/d__14_ xsel_44_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN1_13 XI11_1/XI0/XI0_44/d__13_ xsel_44_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN1_12 XI11_1/XI0/XI0_44/d__12_ xsel_44_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN1_11 XI11_1/XI0/XI0_44/d__11_ xsel_44_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN1_10 XI11_1/XI0/XI0_44/d__10_ xsel_44_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN1_9 XI11_1/XI0/XI0_44/d__9_ xsel_44_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN1_8 XI11_1/XI0/XI0_44/d__8_ xsel_44_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN1_7 XI11_1/XI0/XI0_44/d__7_ xsel_44_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN1_6 XI11_1/XI0/XI0_44/d__6_ xsel_44_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN1_5 XI11_1/XI0/XI0_44/d__5_ xsel_44_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN1_4 XI11_1/XI0/XI0_44/d__4_ xsel_44_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN1_3 XI11_1/XI0/XI0_44/d__3_ xsel_44_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN1_2 XI11_1/XI0/XI0_44/d__2_ xsel_44_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN1_1 XI11_1/XI0/XI0_44/d__1_ xsel_44_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_44/MN1_0 XI11_1/XI0/XI0_44/d__0_ xsel_44_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN0_15 XI11_1/net21_0_ xsel_43_ XI11_1/XI0/XI0_43/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN0_14 XI11_1/net21_1_ xsel_43_ XI11_1/XI0/XI0_43/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN0_13 XI11_1/net21_2_ xsel_43_ XI11_1/XI0/XI0_43/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN0_12 XI11_1/net21_3_ xsel_43_ XI11_1/XI0/XI0_43/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN0_11 XI11_1/net21_4_ xsel_43_ XI11_1/XI0/XI0_43/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN0_10 XI11_1/net21_5_ xsel_43_ XI11_1/XI0/XI0_43/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN0_9 XI11_1/net21_6_ xsel_43_ XI11_1/XI0/XI0_43/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN0_8 XI11_1/net21_7_ xsel_43_ XI11_1/XI0/XI0_43/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN0_7 XI11_1/net21_8_ xsel_43_ XI11_1/XI0/XI0_43/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN0_6 XI11_1/net21_9_ xsel_43_ XI11_1/XI0/XI0_43/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN0_5 XI11_1/net21_10_ xsel_43_ XI11_1/XI0/XI0_43/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN0_4 XI11_1/net21_11_ xsel_43_ XI11_1/XI0/XI0_43/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN0_3 XI11_1/net21_12_ xsel_43_ XI11_1/XI0/XI0_43/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN0_2 XI11_1/net21_13_ xsel_43_ XI11_1/XI0/XI0_43/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN0_1 XI11_1/net21_14_ xsel_43_ XI11_1/XI0/XI0_43/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN0_0 XI11_1/net21_15_ xsel_43_ XI11_1/XI0/XI0_43/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN1_15 XI11_1/XI0/XI0_43/d__15_ xsel_43_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN1_14 XI11_1/XI0/XI0_43/d__14_ xsel_43_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN1_13 XI11_1/XI0/XI0_43/d__13_ xsel_43_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN1_12 XI11_1/XI0/XI0_43/d__12_ xsel_43_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN1_11 XI11_1/XI0/XI0_43/d__11_ xsel_43_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN1_10 XI11_1/XI0/XI0_43/d__10_ xsel_43_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN1_9 XI11_1/XI0/XI0_43/d__9_ xsel_43_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN1_8 XI11_1/XI0/XI0_43/d__8_ xsel_43_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN1_7 XI11_1/XI0/XI0_43/d__7_ xsel_43_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN1_6 XI11_1/XI0/XI0_43/d__6_ xsel_43_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN1_5 XI11_1/XI0/XI0_43/d__5_ xsel_43_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN1_4 XI11_1/XI0/XI0_43/d__4_ xsel_43_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN1_3 XI11_1/XI0/XI0_43/d__3_ xsel_43_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN1_2 XI11_1/XI0/XI0_43/d__2_ xsel_43_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN1_1 XI11_1/XI0/XI0_43/d__1_ xsel_43_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_43/MN1_0 XI11_1/XI0/XI0_43/d__0_ xsel_43_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN0_15 XI11_1/net21_0_ xsel_42_ XI11_1/XI0/XI0_42/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN0_14 XI11_1/net21_1_ xsel_42_ XI11_1/XI0/XI0_42/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN0_13 XI11_1/net21_2_ xsel_42_ XI11_1/XI0/XI0_42/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN0_12 XI11_1/net21_3_ xsel_42_ XI11_1/XI0/XI0_42/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN0_11 XI11_1/net21_4_ xsel_42_ XI11_1/XI0/XI0_42/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN0_10 XI11_1/net21_5_ xsel_42_ XI11_1/XI0/XI0_42/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN0_9 XI11_1/net21_6_ xsel_42_ XI11_1/XI0/XI0_42/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN0_8 XI11_1/net21_7_ xsel_42_ XI11_1/XI0/XI0_42/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN0_7 XI11_1/net21_8_ xsel_42_ XI11_1/XI0/XI0_42/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN0_6 XI11_1/net21_9_ xsel_42_ XI11_1/XI0/XI0_42/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN0_5 XI11_1/net21_10_ xsel_42_ XI11_1/XI0/XI0_42/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN0_4 XI11_1/net21_11_ xsel_42_ XI11_1/XI0/XI0_42/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN0_3 XI11_1/net21_12_ xsel_42_ XI11_1/XI0/XI0_42/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN0_2 XI11_1/net21_13_ xsel_42_ XI11_1/XI0/XI0_42/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN0_1 XI11_1/net21_14_ xsel_42_ XI11_1/XI0/XI0_42/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN0_0 XI11_1/net21_15_ xsel_42_ XI11_1/XI0/XI0_42/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN1_15 XI11_1/XI0/XI0_42/d__15_ xsel_42_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN1_14 XI11_1/XI0/XI0_42/d__14_ xsel_42_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN1_13 XI11_1/XI0/XI0_42/d__13_ xsel_42_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN1_12 XI11_1/XI0/XI0_42/d__12_ xsel_42_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN1_11 XI11_1/XI0/XI0_42/d__11_ xsel_42_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN1_10 XI11_1/XI0/XI0_42/d__10_ xsel_42_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN1_9 XI11_1/XI0/XI0_42/d__9_ xsel_42_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN1_8 XI11_1/XI0/XI0_42/d__8_ xsel_42_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN1_7 XI11_1/XI0/XI0_42/d__7_ xsel_42_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN1_6 XI11_1/XI0/XI0_42/d__6_ xsel_42_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN1_5 XI11_1/XI0/XI0_42/d__5_ xsel_42_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN1_4 XI11_1/XI0/XI0_42/d__4_ xsel_42_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN1_3 XI11_1/XI0/XI0_42/d__3_ xsel_42_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN1_2 XI11_1/XI0/XI0_42/d__2_ xsel_42_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN1_1 XI11_1/XI0/XI0_42/d__1_ xsel_42_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_42/MN1_0 XI11_1/XI0/XI0_42/d__0_ xsel_42_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN0_15 XI11_1/net21_0_ xsel_41_ XI11_1/XI0/XI0_41/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN0_14 XI11_1/net21_1_ xsel_41_ XI11_1/XI0/XI0_41/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN0_13 XI11_1/net21_2_ xsel_41_ XI11_1/XI0/XI0_41/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN0_12 XI11_1/net21_3_ xsel_41_ XI11_1/XI0/XI0_41/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN0_11 XI11_1/net21_4_ xsel_41_ XI11_1/XI0/XI0_41/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN0_10 XI11_1/net21_5_ xsel_41_ XI11_1/XI0/XI0_41/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN0_9 XI11_1/net21_6_ xsel_41_ XI11_1/XI0/XI0_41/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN0_8 XI11_1/net21_7_ xsel_41_ XI11_1/XI0/XI0_41/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN0_7 XI11_1/net21_8_ xsel_41_ XI11_1/XI0/XI0_41/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN0_6 XI11_1/net21_9_ xsel_41_ XI11_1/XI0/XI0_41/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN0_5 XI11_1/net21_10_ xsel_41_ XI11_1/XI0/XI0_41/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN0_4 XI11_1/net21_11_ xsel_41_ XI11_1/XI0/XI0_41/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN0_3 XI11_1/net21_12_ xsel_41_ XI11_1/XI0/XI0_41/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN0_2 XI11_1/net21_13_ xsel_41_ XI11_1/XI0/XI0_41/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN0_1 XI11_1/net21_14_ xsel_41_ XI11_1/XI0/XI0_41/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN0_0 XI11_1/net21_15_ xsel_41_ XI11_1/XI0/XI0_41/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN1_15 XI11_1/XI0/XI0_41/d__15_ xsel_41_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN1_14 XI11_1/XI0/XI0_41/d__14_ xsel_41_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN1_13 XI11_1/XI0/XI0_41/d__13_ xsel_41_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN1_12 XI11_1/XI0/XI0_41/d__12_ xsel_41_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN1_11 XI11_1/XI0/XI0_41/d__11_ xsel_41_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN1_10 XI11_1/XI0/XI0_41/d__10_ xsel_41_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN1_9 XI11_1/XI0/XI0_41/d__9_ xsel_41_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN1_8 XI11_1/XI0/XI0_41/d__8_ xsel_41_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN1_7 XI11_1/XI0/XI0_41/d__7_ xsel_41_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN1_6 XI11_1/XI0/XI0_41/d__6_ xsel_41_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN1_5 XI11_1/XI0/XI0_41/d__5_ xsel_41_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN1_4 XI11_1/XI0/XI0_41/d__4_ xsel_41_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN1_3 XI11_1/XI0/XI0_41/d__3_ xsel_41_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN1_2 XI11_1/XI0/XI0_41/d__2_ xsel_41_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN1_1 XI11_1/XI0/XI0_41/d__1_ xsel_41_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_41/MN1_0 XI11_1/XI0/XI0_41/d__0_ xsel_41_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN0_15 XI11_1/net21_0_ xsel_40_ XI11_1/XI0/XI0_40/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN0_14 XI11_1/net21_1_ xsel_40_ XI11_1/XI0/XI0_40/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN0_13 XI11_1/net21_2_ xsel_40_ XI11_1/XI0/XI0_40/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN0_12 XI11_1/net21_3_ xsel_40_ XI11_1/XI0/XI0_40/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN0_11 XI11_1/net21_4_ xsel_40_ XI11_1/XI0/XI0_40/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN0_10 XI11_1/net21_5_ xsel_40_ XI11_1/XI0/XI0_40/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN0_9 XI11_1/net21_6_ xsel_40_ XI11_1/XI0/XI0_40/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN0_8 XI11_1/net21_7_ xsel_40_ XI11_1/XI0/XI0_40/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN0_7 XI11_1/net21_8_ xsel_40_ XI11_1/XI0/XI0_40/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN0_6 XI11_1/net21_9_ xsel_40_ XI11_1/XI0/XI0_40/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN0_5 XI11_1/net21_10_ xsel_40_ XI11_1/XI0/XI0_40/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN0_4 XI11_1/net21_11_ xsel_40_ XI11_1/XI0/XI0_40/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN0_3 XI11_1/net21_12_ xsel_40_ XI11_1/XI0/XI0_40/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN0_2 XI11_1/net21_13_ xsel_40_ XI11_1/XI0/XI0_40/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN0_1 XI11_1/net21_14_ xsel_40_ XI11_1/XI0/XI0_40/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN0_0 XI11_1/net21_15_ xsel_40_ XI11_1/XI0/XI0_40/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN1_15 XI11_1/XI0/XI0_40/d__15_ xsel_40_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN1_14 XI11_1/XI0/XI0_40/d__14_ xsel_40_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN1_13 XI11_1/XI0/XI0_40/d__13_ xsel_40_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN1_12 XI11_1/XI0/XI0_40/d__12_ xsel_40_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN1_11 XI11_1/XI0/XI0_40/d__11_ xsel_40_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN1_10 XI11_1/XI0/XI0_40/d__10_ xsel_40_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN1_9 XI11_1/XI0/XI0_40/d__9_ xsel_40_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN1_8 XI11_1/XI0/XI0_40/d__8_ xsel_40_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN1_7 XI11_1/XI0/XI0_40/d__7_ xsel_40_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN1_6 XI11_1/XI0/XI0_40/d__6_ xsel_40_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN1_5 XI11_1/XI0/XI0_40/d__5_ xsel_40_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN1_4 XI11_1/XI0/XI0_40/d__4_ xsel_40_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN1_3 XI11_1/XI0/XI0_40/d__3_ xsel_40_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN1_2 XI11_1/XI0/XI0_40/d__2_ xsel_40_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN1_1 XI11_1/XI0/XI0_40/d__1_ xsel_40_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_40/MN1_0 XI11_1/XI0/XI0_40/d__0_ xsel_40_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN0_15 XI11_1/net21_0_ xsel_39_ XI11_1/XI0/XI0_39/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN0_14 XI11_1/net21_1_ xsel_39_ XI11_1/XI0/XI0_39/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN0_13 XI11_1/net21_2_ xsel_39_ XI11_1/XI0/XI0_39/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN0_12 XI11_1/net21_3_ xsel_39_ XI11_1/XI0/XI0_39/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN0_11 XI11_1/net21_4_ xsel_39_ XI11_1/XI0/XI0_39/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN0_10 XI11_1/net21_5_ xsel_39_ XI11_1/XI0/XI0_39/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN0_9 XI11_1/net21_6_ xsel_39_ XI11_1/XI0/XI0_39/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN0_8 XI11_1/net21_7_ xsel_39_ XI11_1/XI0/XI0_39/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN0_7 XI11_1/net21_8_ xsel_39_ XI11_1/XI0/XI0_39/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN0_6 XI11_1/net21_9_ xsel_39_ XI11_1/XI0/XI0_39/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN0_5 XI11_1/net21_10_ xsel_39_ XI11_1/XI0/XI0_39/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN0_4 XI11_1/net21_11_ xsel_39_ XI11_1/XI0/XI0_39/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN0_3 XI11_1/net21_12_ xsel_39_ XI11_1/XI0/XI0_39/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN0_2 XI11_1/net21_13_ xsel_39_ XI11_1/XI0/XI0_39/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN0_1 XI11_1/net21_14_ xsel_39_ XI11_1/XI0/XI0_39/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN0_0 XI11_1/net21_15_ xsel_39_ XI11_1/XI0/XI0_39/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN1_15 XI11_1/XI0/XI0_39/d__15_ xsel_39_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN1_14 XI11_1/XI0/XI0_39/d__14_ xsel_39_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN1_13 XI11_1/XI0/XI0_39/d__13_ xsel_39_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN1_12 XI11_1/XI0/XI0_39/d__12_ xsel_39_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN1_11 XI11_1/XI0/XI0_39/d__11_ xsel_39_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN1_10 XI11_1/XI0/XI0_39/d__10_ xsel_39_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN1_9 XI11_1/XI0/XI0_39/d__9_ xsel_39_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN1_8 XI11_1/XI0/XI0_39/d__8_ xsel_39_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN1_7 XI11_1/XI0/XI0_39/d__7_ xsel_39_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN1_6 XI11_1/XI0/XI0_39/d__6_ xsel_39_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN1_5 XI11_1/XI0/XI0_39/d__5_ xsel_39_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN1_4 XI11_1/XI0/XI0_39/d__4_ xsel_39_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN1_3 XI11_1/XI0/XI0_39/d__3_ xsel_39_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN1_2 XI11_1/XI0/XI0_39/d__2_ xsel_39_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN1_1 XI11_1/XI0/XI0_39/d__1_ xsel_39_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_39/MN1_0 XI11_1/XI0/XI0_39/d__0_ xsel_39_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN0_15 XI11_1/net21_0_ xsel_38_ XI11_1/XI0/XI0_38/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN0_14 XI11_1/net21_1_ xsel_38_ XI11_1/XI0/XI0_38/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN0_13 XI11_1/net21_2_ xsel_38_ XI11_1/XI0/XI0_38/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN0_12 XI11_1/net21_3_ xsel_38_ XI11_1/XI0/XI0_38/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN0_11 XI11_1/net21_4_ xsel_38_ XI11_1/XI0/XI0_38/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN0_10 XI11_1/net21_5_ xsel_38_ XI11_1/XI0/XI0_38/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN0_9 XI11_1/net21_6_ xsel_38_ XI11_1/XI0/XI0_38/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN0_8 XI11_1/net21_7_ xsel_38_ XI11_1/XI0/XI0_38/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN0_7 XI11_1/net21_8_ xsel_38_ XI11_1/XI0/XI0_38/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN0_6 XI11_1/net21_9_ xsel_38_ XI11_1/XI0/XI0_38/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN0_5 XI11_1/net21_10_ xsel_38_ XI11_1/XI0/XI0_38/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN0_4 XI11_1/net21_11_ xsel_38_ XI11_1/XI0/XI0_38/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN0_3 XI11_1/net21_12_ xsel_38_ XI11_1/XI0/XI0_38/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN0_2 XI11_1/net21_13_ xsel_38_ XI11_1/XI0/XI0_38/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN0_1 XI11_1/net21_14_ xsel_38_ XI11_1/XI0/XI0_38/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN0_0 XI11_1/net21_15_ xsel_38_ XI11_1/XI0/XI0_38/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN1_15 XI11_1/XI0/XI0_38/d__15_ xsel_38_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN1_14 XI11_1/XI0/XI0_38/d__14_ xsel_38_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN1_13 XI11_1/XI0/XI0_38/d__13_ xsel_38_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN1_12 XI11_1/XI0/XI0_38/d__12_ xsel_38_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN1_11 XI11_1/XI0/XI0_38/d__11_ xsel_38_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN1_10 XI11_1/XI0/XI0_38/d__10_ xsel_38_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN1_9 XI11_1/XI0/XI0_38/d__9_ xsel_38_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN1_8 XI11_1/XI0/XI0_38/d__8_ xsel_38_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN1_7 XI11_1/XI0/XI0_38/d__7_ xsel_38_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN1_6 XI11_1/XI0/XI0_38/d__6_ xsel_38_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN1_5 XI11_1/XI0/XI0_38/d__5_ xsel_38_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN1_4 XI11_1/XI0/XI0_38/d__4_ xsel_38_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN1_3 XI11_1/XI0/XI0_38/d__3_ xsel_38_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN1_2 XI11_1/XI0/XI0_38/d__2_ xsel_38_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN1_1 XI11_1/XI0/XI0_38/d__1_ xsel_38_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_38/MN1_0 XI11_1/XI0/XI0_38/d__0_ xsel_38_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN0_15 XI11_1/net21_0_ xsel_37_ XI11_1/XI0/XI0_37/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN0_14 XI11_1/net21_1_ xsel_37_ XI11_1/XI0/XI0_37/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN0_13 XI11_1/net21_2_ xsel_37_ XI11_1/XI0/XI0_37/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN0_12 XI11_1/net21_3_ xsel_37_ XI11_1/XI0/XI0_37/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN0_11 XI11_1/net21_4_ xsel_37_ XI11_1/XI0/XI0_37/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN0_10 XI11_1/net21_5_ xsel_37_ XI11_1/XI0/XI0_37/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN0_9 XI11_1/net21_6_ xsel_37_ XI11_1/XI0/XI0_37/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN0_8 XI11_1/net21_7_ xsel_37_ XI11_1/XI0/XI0_37/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN0_7 XI11_1/net21_8_ xsel_37_ XI11_1/XI0/XI0_37/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN0_6 XI11_1/net21_9_ xsel_37_ XI11_1/XI0/XI0_37/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN0_5 XI11_1/net21_10_ xsel_37_ XI11_1/XI0/XI0_37/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN0_4 XI11_1/net21_11_ xsel_37_ XI11_1/XI0/XI0_37/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN0_3 XI11_1/net21_12_ xsel_37_ XI11_1/XI0/XI0_37/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN0_2 XI11_1/net21_13_ xsel_37_ XI11_1/XI0/XI0_37/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN0_1 XI11_1/net21_14_ xsel_37_ XI11_1/XI0/XI0_37/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN0_0 XI11_1/net21_15_ xsel_37_ XI11_1/XI0/XI0_37/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN1_15 XI11_1/XI0/XI0_37/d__15_ xsel_37_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN1_14 XI11_1/XI0/XI0_37/d__14_ xsel_37_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN1_13 XI11_1/XI0/XI0_37/d__13_ xsel_37_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN1_12 XI11_1/XI0/XI0_37/d__12_ xsel_37_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN1_11 XI11_1/XI0/XI0_37/d__11_ xsel_37_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN1_10 XI11_1/XI0/XI0_37/d__10_ xsel_37_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN1_9 XI11_1/XI0/XI0_37/d__9_ xsel_37_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN1_8 XI11_1/XI0/XI0_37/d__8_ xsel_37_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN1_7 XI11_1/XI0/XI0_37/d__7_ xsel_37_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN1_6 XI11_1/XI0/XI0_37/d__6_ xsel_37_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN1_5 XI11_1/XI0/XI0_37/d__5_ xsel_37_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN1_4 XI11_1/XI0/XI0_37/d__4_ xsel_37_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN1_3 XI11_1/XI0/XI0_37/d__3_ xsel_37_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN1_2 XI11_1/XI0/XI0_37/d__2_ xsel_37_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN1_1 XI11_1/XI0/XI0_37/d__1_ xsel_37_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_37/MN1_0 XI11_1/XI0/XI0_37/d__0_ xsel_37_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN0_15 XI11_1/net21_0_ xsel_36_ XI11_1/XI0/XI0_36/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN0_14 XI11_1/net21_1_ xsel_36_ XI11_1/XI0/XI0_36/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN0_13 XI11_1/net21_2_ xsel_36_ XI11_1/XI0/XI0_36/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN0_12 XI11_1/net21_3_ xsel_36_ XI11_1/XI0/XI0_36/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN0_11 XI11_1/net21_4_ xsel_36_ XI11_1/XI0/XI0_36/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN0_10 XI11_1/net21_5_ xsel_36_ XI11_1/XI0/XI0_36/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN0_9 XI11_1/net21_6_ xsel_36_ XI11_1/XI0/XI0_36/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN0_8 XI11_1/net21_7_ xsel_36_ XI11_1/XI0/XI0_36/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN0_7 XI11_1/net21_8_ xsel_36_ XI11_1/XI0/XI0_36/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN0_6 XI11_1/net21_9_ xsel_36_ XI11_1/XI0/XI0_36/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN0_5 XI11_1/net21_10_ xsel_36_ XI11_1/XI0/XI0_36/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN0_4 XI11_1/net21_11_ xsel_36_ XI11_1/XI0/XI0_36/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN0_3 XI11_1/net21_12_ xsel_36_ XI11_1/XI0/XI0_36/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN0_2 XI11_1/net21_13_ xsel_36_ XI11_1/XI0/XI0_36/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN0_1 XI11_1/net21_14_ xsel_36_ XI11_1/XI0/XI0_36/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN0_0 XI11_1/net21_15_ xsel_36_ XI11_1/XI0/XI0_36/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN1_15 XI11_1/XI0/XI0_36/d__15_ xsel_36_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN1_14 XI11_1/XI0/XI0_36/d__14_ xsel_36_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN1_13 XI11_1/XI0/XI0_36/d__13_ xsel_36_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN1_12 XI11_1/XI0/XI0_36/d__12_ xsel_36_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN1_11 XI11_1/XI0/XI0_36/d__11_ xsel_36_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN1_10 XI11_1/XI0/XI0_36/d__10_ xsel_36_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN1_9 XI11_1/XI0/XI0_36/d__9_ xsel_36_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN1_8 XI11_1/XI0/XI0_36/d__8_ xsel_36_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN1_7 XI11_1/XI0/XI0_36/d__7_ xsel_36_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN1_6 XI11_1/XI0/XI0_36/d__6_ xsel_36_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN1_5 XI11_1/XI0/XI0_36/d__5_ xsel_36_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN1_4 XI11_1/XI0/XI0_36/d__4_ xsel_36_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN1_3 XI11_1/XI0/XI0_36/d__3_ xsel_36_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN1_2 XI11_1/XI0/XI0_36/d__2_ xsel_36_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN1_1 XI11_1/XI0/XI0_36/d__1_ xsel_36_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_36/MN1_0 XI11_1/XI0/XI0_36/d__0_ xsel_36_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN0_15 XI11_1/net21_0_ xsel_35_ XI11_1/XI0/XI0_35/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN0_14 XI11_1/net21_1_ xsel_35_ XI11_1/XI0/XI0_35/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN0_13 XI11_1/net21_2_ xsel_35_ XI11_1/XI0/XI0_35/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN0_12 XI11_1/net21_3_ xsel_35_ XI11_1/XI0/XI0_35/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN0_11 XI11_1/net21_4_ xsel_35_ XI11_1/XI0/XI0_35/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN0_10 XI11_1/net21_5_ xsel_35_ XI11_1/XI0/XI0_35/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN0_9 XI11_1/net21_6_ xsel_35_ XI11_1/XI0/XI0_35/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN0_8 XI11_1/net21_7_ xsel_35_ XI11_1/XI0/XI0_35/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN0_7 XI11_1/net21_8_ xsel_35_ XI11_1/XI0/XI0_35/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN0_6 XI11_1/net21_9_ xsel_35_ XI11_1/XI0/XI0_35/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN0_5 XI11_1/net21_10_ xsel_35_ XI11_1/XI0/XI0_35/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN0_4 XI11_1/net21_11_ xsel_35_ XI11_1/XI0/XI0_35/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN0_3 XI11_1/net21_12_ xsel_35_ XI11_1/XI0/XI0_35/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN0_2 XI11_1/net21_13_ xsel_35_ XI11_1/XI0/XI0_35/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN0_1 XI11_1/net21_14_ xsel_35_ XI11_1/XI0/XI0_35/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN0_0 XI11_1/net21_15_ xsel_35_ XI11_1/XI0/XI0_35/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN1_15 XI11_1/XI0/XI0_35/d__15_ xsel_35_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN1_14 XI11_1/XI0/XI0_35/d__14_ xsel_35_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN1_13 XI11_1/XI0/XI0_35/d__13_ xsel_35_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN1_12 XI11_1/XI0/XI0_35/d__12_ xsel_35_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN1_11 XI11_1/XI0/XI0_35/d__11_ xsel_35_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN1_10 XI11_1/XI0/XI0_35/d__10_ xsel_35_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN1_9 XI11_1/XI0/XI0_35/d__9_ xsel_35_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN1_8 XI11_1/XI0/XI0_35/d__8_ xsel_35_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN1_7 XI11_1/XI0/XI0_35/d__7_ xsel_35_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN1_6 XI11_1/XI0/XI0_35/d__6_ xsel_35_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN1_5 XI11_1/XI0/XI0_35/d__5_ xsel_35_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN1_4 XI11_1/XI0/XI0_35/d__4_ xsel_35_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN1_3 XI11_1/XI0/XI0_35/d__3_ xsel_35_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN1_2 XI11_1/XI0/XI0_35/d__2_ xsel_35_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN1_1 XI11_1/XI0/XI0_35/d__1_ xsel_35_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_35/MN1_0 XI11_1/XI0/XI0_35/d__0_ xsel_35_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN0_15 XI11_1/net21_0_ xsel_34_ XI11_1/XI0/XI0_34/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN0_14 XI11_1/net21_1_ xsel_34_ XI11_1/XI0/XI0_34/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN0_13 XI11_1/net21_2_ xsel_34_ XI11_1/XI0/XI0_34/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN0_12 XI11_1/net21_3_ xsel_34_ XI11_1/XI0/XI0_34/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN0_11 XI11_1/net21_4_ xsel_34_ XI11_1/XI0/XI0_34/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN0_10 XI11_1/net21_5_ xsel_34_ XI11_1/XI0/XI0_34/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN0_9 XI11_1/net21_6_ xsel_34_ XI11_1/XI0/XI0_34/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN0_8 XI11_1/net21_7_ xsel_34_ XI11_1/XI0/XI0_34/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN0_7 XI11_1/net21_8_ xsel_34_ XI11_1/XI0/XI0_34/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN0_6 XI11_1/net21_9_ xsel_34_ XI11_1/XI0/XI0_34/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN0_5 XI11_1/net21_10_ xsel_34_ XI11_1/XI0/XI0_34/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN0_4 XI11_1/net21_11_ xsel_34_ XI11_1/XI0/XI0_34/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN0_3 XI11_1/net21_12_ xsel_34_ XI11_1/XI0/XI0_34/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN0_2 XI11_1/net21_13_ xsel_34_ XI11_1/XI0/XI0_34/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN0_1 XI11_1/net21_14_ xsel_34_ XI11_1/XI0/XI0_34/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN0_0 XI11_1/net21_15_ xsel_34_ XI11_1/XI0/XI0_34/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN1_15 XI11_1/XI0/XI0_34/d__15_ xsel_34_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN1_14 XI11_1/XI0/XI0_34/d__14_ xsel_34_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN1_13 XI11_1/XI0/XI0_34/d__13_ xsel_34_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN1_12 XI11_1/XI0/XI0_34/d__12_ xsel_34_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN1_11 XI11_1/XI0/XI0_34/d__11_ xsel_34_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN1_10 XI11_1/XI0/XI0_34/d__10_ xsel_34_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN1_9 XI11_1/XI0/XI0_34/d__9_ xsel_34_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN1_8 XI11_1/XI0/XI0_34/d__8_ xsel_34_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN1_7 XI11_1/XI0/XI0_34/d__7_ xsel_34_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN1_6 XI11_1/XI0/XI0_34/d__6_ xsel_34_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN1_5 XI11_1/XI0/XI0_34/d__5_ xsel_34_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN1_4 XI11_1/XI0/XI0_34/d__4_ xsel_34_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN1_3 XI11_1/XI0/XI0_34/d__3_ xsel_34_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN1_2 XI11_1/XI0/XI0_34/d__2_ xsel_34_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN1_1 XI11_1/XI0/XI0_34/d__1_ xsel_34_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_34/MN1_0 XI11_1/XI0/XI0_34/d__0_ xsel_34_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN0_15 XI11_1/net21_0_ xsel_33_ XI11_1/XI0/XI0_33/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN0_14 XI11_1/net21_1_ xsel_33_ XI11_1/XI0/XI0_33/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN0_13 XI11_1/net21_2_ xsel_33_ XI11_1/XI0/XI0_33/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN0_12 XI11_1/net21_3_ xsel_33_ XI11_1/XI0/XI0_33/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN0_11 XI11_1/net21_4_ xsel_33_ XI11_1/XI0/XI0_33/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN0_10 XI11_1/net21_5_ xsel_33_ XI11_1/XI0/XI0_33/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN0_9 XI11_1/net21_6_ xsel_33_ XI11_1/XI0/XI0_33/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN0_8 XI11_1/net21_7_ xsel_33_ XI11_1/XI0/XI0_33/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN0_7 XI11_1/net21_8_ xsel_33_ XI11_1/XI0/XI0_33/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN0_6 XI11_1/net21_9_ xsel_33_ XI11_1/XI0/XI0_33/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN0_5 XI11_1/net21_10_ xsel_33_ XI11_1/XI0/XI0_33/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN0_4 XI11_1/net21_11_ xsel_33_ XI11_1/XI0/XI0_33/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN0_3 XI11_1/net21_12_ xsel_33_ XI11_1/XI0/XI0_33/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN0_2 XI11_1/net21_13_ xsel_33_ XI11_1/XI0/XI0_33/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN0_1 XI11_1/net21_14_ xsel_33_ XI11_1/XI0/XI0_33/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN0_0 XI11_1/net21_15_ xsel_33_ XI11_1/XI0/XI0_33/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN1_15 XI11_1/XI0/XI0_33/d__15_ xsel_33_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN1_14 XI11_1/XI0/XI0_33/d__14_ xsel_33_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN1_13 XI11_1/XI0/XI0_33/d__13_ xsel_33_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN1_12 XI11_1/XI0/XI0_33/d__12_ xsel_33_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN1_11 XI11_1/XI0/XI0_33/d__11_ xsel_33_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN1_10 XI11_1/XI0/XI0_33/d__10_ xsel_33_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN1_9 XI11_1/XI0/XI0_33/d__9_ xsel_33_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN1_8 XI11_1/XI0/XI0_33/d__8_ xsel_33_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN1_7 XI11_1/XI0/XI0_33/d__7_ xsel_33_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN1_6 XI11_1/XI0/XI0_33/d__6_ xsel_33_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN1_5 XI11_1/XI0/XI0_33/d__5_ xsel_33_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN1_4 XI11_1/XI0/XI0_33/d__4_ xsel_33_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN1_3 XI11_1/XI0/XI0_33/d__3_ xsel_33_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN1_2 XI11_1/XI0/XI0_33/d__2_ xsel_33_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN1_1 XI11_1/XI0/XI0_33/d__1_ xsel_33_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_33/MN1_0 XI11_1/XI0/XI0_33/d__0_ xsel_33_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN0_15 XI11_1/net21_0_ xsel_32_ XI11_1/XI0/XI0_32/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN0_14 XI11_1/net21_1_ xsel_32_ XI11_1/XI0/XI0_32/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN0_13 XI11_1/net21_2_ xsel_32_ XI11_1/XI0/XI0_32/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN0_12 XI11_1/net21_3_ xsel_32_ XI11_1/XI0/XI0_32/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN0_11 XI11_1/net21_4_ xsel_32_ XI11_1/XI0/XI0_32/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN0_10 XI11_1/net21_5_ xsel_32_ XI11_1/XI0/XI0_32/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN0_9 XI11_1/net21_6_ xsel_32_ XI11_1/XI0/XI0_32/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN0_8 XI11_1/net21_7_ xsel_32_ XI11_1/XI0/XI0_32/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN0_7 XI11_1/net21_8_ xsel_32_ XI11_1/XI0/XI0_32/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN0_6 XI11_1/net21_9_ xsel_32_ XI11_1/XI0/XI0_32/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN0_5 XI11_1/net21_10_ xsel_32_ XI11_1/XI0/XI0_32/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN0_4 XI11_1/net21_11_ xsel_32_ XI11_1/XI0/XI0_32/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN0_3 XI11_1/net21_12_ xsel_32_ XI11_1/XI0/XI0_32/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN0_2 XI11_1/net21_13_ xsel_32_ XI11_1/XI0/XI0_32/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN0_1 XI11_1/net21_14_ xsel_32_ XI11_1/XI0/XI0_32/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN0_0 XI11_1/net21_15_ xsel_32_ XI11_1/XI0/XI0_32/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN1_15 XI11_1/XI0/XI0_32/d__15_ xsel_32_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN1_14 XI11_1/XI0/XI0_32/d__14_ xsel_32_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN1_13 XI11_1/XI0/XI0_32/d__13_ xsel_32_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN1_12 XI11_1/XI0/XI0_32/d__12_ xsel_32_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN1_11 XI11_1/XI0/XI0_32/d__11_ xsel_32_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN1_10 XI11_1/XI0/XI0_32/d__10_ xsel_32_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN1_9 XI11_1/XI0/XI0_32/d__9_ xsel_32_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN1_8 XI11_1/XI0/XI0_32/d__8_ xsel_32_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN1_7 XI11_1/XI0/XI0_32/d__7_ xsel_32_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN1_6 XI11_1/XI0/XI0_32/d__6_ xsel_32_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN1_5 XI11_1/XI0/XI0_32/d__5_ xsel_32_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN1_4 XI11_1/XI0/XI0_32/d__4_ xsel_32_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN1_3 XI11_1/XI0/XI0_32/d__3_ xsel_32_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN1_2 XI11_1/XI0/XI0_32/d__2_ xsel_32_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN1_1 XI11_1/XI0/XI0_32/d__1_ xsel_32_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_32/MN1_0 XI11_1/XI0/XI0_32/d__0_ xsel_32_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN0_15 XI11_1/net21_0_ xsel_31_ XI11_1/XI0/XI0_31/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN0_14 XI11_1/net21_1_ xsel_31_ XI11_1/XI0/XI0_31/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN0_13 XI11_1/net21_2_ xsel_31_ XI11_1/XI0/XI0_31/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN0_12 XI11_1/net21_3_ xsel_31_ XI11_1/XI0/XI0_31/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN0_11 XI11_1/net21_4_ xsel_31_ XI11_1/XI0/XI0_31/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN0_10 XI11_1/net21_5_ xsel_31_ XI11_1/XI0/XI0_31/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN0_9 XI11_1/net21_6_ xsel_31_ XI11_1/XI0/XI0_31/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN0_8 XI11_1/net21_7_ xsel_31_ XI11_1/XI0/XI0_31/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN0_7 XI11_1/net21_8_ xsel_31_ XI11_1/XI0/XI0_31/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN0_6 XI11_1/net21_9_ xsel_31_ XI11_1/XI0/XI0_31/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN0_5 XI11_1/net21_10_ xsel_31_ XI11_1/XI0/XI0_31/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN0_4 XI11_1/net21_11_ xsel_31_ XI11_1/XI0/XI0_31/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN0_3 XI11_1/net21_12_ xsel_31_ XI11_1/XI0/XI0_31/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN0_2 XI11_1/net21_13_ xsel_31_ XI11_1/XI0/XI0_31/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN0_1 XI11_1/net21_14_ xsel_31_ XI11_1/XI0/XI0_31/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN0_0 XI11_1/net21_15_ xsel_31_ XI11_1/XI0/XI0_31/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN1_15 XI11_1/XI0/XI0_31/d__15_ xsel_31_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN1_14 XI11_1/XI0/XI0_31/d__14_ xsel_31_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN1_13 XI11_1/XI0/XI0_31/d__13_ xsel_31_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN1_12 XI11_1/XI0/XI0_31/d__12_ xsel_31_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN1_11 XI11_1/XI0/XI0_31/d__11_ xsel_31_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN1_10 XI11_1/XI0/XI0_31/d__10_ xsel_31_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN1_9 XI11_1/XI0/XI0_31/d__9_ xsel_31_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN1_8 XI11_1/XI0/XI0_31/d__8_ xsel_31_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN1_7 XI11_1/XI0/XI0_31/d__7_ xsel_31_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN1_6 XI11_1/XI0/XI0_31/d__6_ xsel_31_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN1_5 XI11_1/XI0/XI0_31/d__5_ xsel_31_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN1_4 XI11_1/XI0/XI0_31/d__4_ xsel_31_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN1_3 XI11_1/XI0/XI0_31/d__3_ xsel_31_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN1_2 XI11_1/XI0/XI0_31/d__2_ xsel_31_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN1_1 XI11_1/XI0/XI0_31/d__1_ xsel_31_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_31/MN1_0 XI11_1/XI0/XI0_31/d__0_ xsel_31_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN0_15 XI11_1/net21_0_ xsel_30_ XI11_1/XI0/XI0_30/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN0_14 XI11_1/net21_1_ xsel_30_ XI11_1/XI0/XI0_30/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN0_13 XI11_1/net21_2_ xsel_30_ XI11_1/XI0/XI0_30/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN0_12 XI11_1/net21_3_ xsel_30_ XI11_1/XI0/XI0_30/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN0_11 XI11_1/net21_4_ xsel_30_ XI11_1/XI0/XI0_30/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN0_10 XI11_1/net21_5_ xsel_30_ XI11_1/XI0/XI0_30/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN0_9 XI11_1/net21_6_ xsel_30_ XI11_1/XI0/XI0_30/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN0_8 XI11_1/net21_7_ xsel_30_ XI11_1/XI0/XI0_30/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN0_7 XI11_1/net21_8_ xsel_30_ XI11_1/XI0/XI0_30/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN0_6 XI11_1/net21_9_ xsel_30_ XI11_1/XI0/XI0_30/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN0_5 XI11_1/net21_10_ xsel_30_ XI11_1/XI0/XI0_30/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN0_4 XI11_1/net21_11_ xsel_30_ XI11_1/XI0/XI0_30/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN0_3 XI11_1/net21_12_ xsel_30_ XI11_1/XI0/XI0_30/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN0_2 XI11_1/net21_13_ xsel_30_ XI11_1/XI0/XI0_30/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN0_1 XI11_1/net21_14_ xsel_30_ XI11_1/XI0/XI0_30/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN0_0 XI11_1/net21_15_ xsel_30_ XI11_1/XI0/XI0_30/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN1_15 XI11_1/XI0/XI0_30/d__15_ xsel_30_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN1_14 XI11_1/XI0/XI0_30/d__14_ xsel_30_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN1_13 XI11_1/XI0/XI0_30/d__13_ xsel_30_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN1_12 XI11_1/XI0/XI0_30/d__12_ xsel_30_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN1_11 XI11_1/XI0/XI0_30/d__11_ xsel_30_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN1_10 XI11_1/XI0/XI0_30/d__10_ xsel_30_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN1_9 XI11_1/XI0/XI0_30/d__9_ xsel_30_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN1_8 XI11_1/XI0/XI0_30/d__8_ xsel_30_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN1_7 XI11_1/XI0/XI0_30/d__7_ xsel_30_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN1_6 XI11_1/XI0/XI0_30/d__6_ xsel_30_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN1_5 XI11_1/XI0/XI0_30/d__5_ xsel_30_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN1_4 XI11_1/XI0/XI0_30/d__4_ xsel_30_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN1_3 XI11_1/XI0/XI0_30/d__3_ xsel_30_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN1_2 XI11_1/XI0/XI0_30/d__2_ xsel_30_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN1_1 XI11_1/XI0/XI0_30/d__1_ xsel_30_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_30/MN1_0 XI11_1/XI0/XI0_30/d__0_ xsel_30_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN0_15 XI11_1/net21_0_ xsel_29_ XI11_1/XI0/XI0_29/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN0_14 XI11_1/net21_1_ xsel_29_ XI11_1/XI0/XI0_29/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN0_13 XI11_1/net21_2_ xsel_29_ XI11_1/XI0/XI0_29/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN0_12 XI11_1/net21_3_ xsel_29_ XI11_1/XI0/XI0_29/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN0_11 XI11_1/net21_4_ xsel_29_ XI11_1/XI0/XI0_29/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN0_10 XI11_1/net21_5_ xsel_29_ XI11_1/XI0/XI0_29/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN0_9 XI11_1/net21_6_ xsel_29_ XI11_1/XI0/XI0_29/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN0_8 XI11_1/net21_7_ xsel_29_ XI11_1/XI0/XI0_29/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN0_7 XI11_1/net21_8_ xsel_29_ XI11_1/XI0/XI0_29/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN0_6 XI11_1/net21_9_ xsel_29_ XI11_1/XI0/XI0_29/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN0_5 XI11_1/net21_10_ xsel_29_ XI11_1/XI0/XI0_29/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN0_4 XI11_1/net21_11_ xsel_29_ XI11_1/XI0/XI0_29/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN0_3 XI11_1/net21_12_ xsel_29_ XI11_1/XI0/XI0_29/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN0_2 XI11_1/net21_13_ xsel_29_ XI11_1/XI0/XI0_29/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN0_1 XI11_1/net21_14_ xsel_29_ XI11_1/XI0/XI0_29/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN0_0 XI11_1/net21_15_ xsel_29_ XI11_1/XI0/XI0_29/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN1_15 XI11_1/XI0/XI0_29/d__15_ xsel_29_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN1_14 XI11_1/XI0/XI0_29/d__14_ xsel_29_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN1_13 XI11_1/XI0/XI0_29/d__13_ xsel_29_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN1_12 XI11_1/XI0/XI0_29/d__12_ xsel_29_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN1_11 XI11_1/XI0/XI0_29/d__11_ xsel_29_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN1_10 XI11_1/XI0/XI0_29/d__10_ xsel_29_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN1_9 XI11_1/XI0/XI0_29/d__9_ xsel_29_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN1_8 XI11_1/XI0/XI0_29/d__8_ xsel_29_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN1_7 XI11_1/XI0/XI0_29/d__7_ xsel_29_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN1_6 XI11_1/XI0/XI0_29/d__6_ xsel_29_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN1_5 XI11_1/XI0/XI0_29/d__5_ xsel_29_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN1_4 XI11_1/XI0/XI0_29/d__4_ xsel_29_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN1_3 XI11_1/XI0/XI0_29/d__3_ xsel_29_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN1_2 XI11_1/XI0/XI0_29/d__2_ xsel_29_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN1_1 XI11_1/XI0/XI0_29/d__1_ xsel_29_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_29/MN1_0 XI11_1/XI0/XI0_29/d__0_ xsel_29_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN0_15 XI11_1/net21_0_ xsel_28_ XI11_1/XI0/XI0_28/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN0_14 XI11_1/net21_1_ xsel_28_ XI11_1/XI0/XI0_28/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN0_13 XI11_1/net21_2_ xsel_28_ XI11_1/XI0/XI0_28/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN0_12 XI11_1/net21_3_ xsel_28_ XI11_1/XI0/XI0_28/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN0_11 XI11_1/net21_4_ xsel_28_ XI11_1/XI0/XI0_28/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN0_10 XI11_1/net21_5_ xsel_28_ XI11_1/XI0/XI0_28/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN0_9 XI11_1/net21_6_ xsel_28_ XI11_1/XI0/XI0_28/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN0_8 XI11_1/net21_7_ xsel_28_ XI11_1/XI0/XI0_28/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN0_7 XI11_1/net21_8_ xsel_28_ XI11_1/XI0/XI0_28/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN0_6 XI11_1/net21_9_ xsel_28_ XI11_1/XI0/XI0_28/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN0_5 XI11_1/net21_10_ xsel_28_ XI11_1/XI0/XI0_28/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN0_4 XI11_1/net21_11_ xsel_28_ XI11_1/XI0/XI0_28/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN0_3 XI11_1/net21_12_ xsel_28_ XI11_1/XI0/XI0_28/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN0_2 XI11_1/net21_13_ xsel_28_ XI11_1/XI0/XI0_28/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN0_1 XI11_1/net21_14_ xsel_28_ XI11_1/XI0/XI0_28/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN0_0 XI11_1/net21_15_ xsel_28_ XI11_1/XI0/XI0_28/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN1_15 XI11_1/XI0/XI0_28/d__15_ xsel_28_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN1_14 XI11_1/XI0/XI0_28/d__14_ xsel_28_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN1_13 XI11_1/XI0/XI0_28/d__13_ xsel_28_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN1_12 XI11_1/XI0/XI0_28/d__12_ xsel_28_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN1_11 XI11_1/XI0/XI0_28/d__11_ xsel_28_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN1_10 XI11_1/XI0/XI0_28/d__10_ xsel_28_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN1_9 XI11_1/XI0/XI0_28/d__9_ xsel_28_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN1_8 XI11_1/XI0/XI0_28/d__8_ xsel_28_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN1_7 XI11_1/XI0/XI0_28/d__7_ xsel_28_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN1_6 XI11_1/XI0/XI0_28/d__6_ xsel_28_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN1_5 XI11_1/XI0/XI0_28/d__5_ xsel_28_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN1_4 XI11_1/XI0/XI0_28/d__4_ xsel_28_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN1_3 XI11_1/XI0/XI0_28/d__3_ xsel_28_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN1_2 XI11_1/XI0/XI0_28/d__2_ xsel_28_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN1_1 XI11_1/XI0/XI0_28/d__1_ xsel_28_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_28/MN1_0 XI11_1/XI0/XI0_28/d__0_ xsel_28_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN0_15 XI11_1/net21_0_ xsel_27_ XI11_1/XI0/XI0_27/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN0_14 XI11_1/net21_1_ xsel_27_ XI11_1/XI0/XI0_27/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN0_13 XI11_1/net21_2_ xsel_27_ XI11_1/XI0/XI0_27/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN0_12 XI11_1/net21_3_ xsel_27_ XI11_1/XI0/XI0_27/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN0_11 XI11_1/net21_4_ xsel_27_ XI11_1/XI0/XI0_27/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN0_10 XI11_1/net21_5_ xsel_27_ XI11_1/XI0/XI0_27/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN0_9 XI11_1/net21_6_ xsel_27_ XI11_1/XI0/XI0_27/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN0_8 XI11_1/net21_7_ xsel_27_ XI11_1/XI0/XI0_27/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN0_7 XI11_1/net21_8_ xsel_27_ XI11_1/XI0/XI0_27/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN0_6 XI11_1/net21_9_ xsel_27_ XI11_1/XI0/XI0_27/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN0_5 XI11_1/net21_10_ xsel_27_ XI11_1/XI0/XI0_27/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN0_4 XI11_1/net21_11_ xsel_27_ XI11_1/XI0/XI0_27/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN0_3 XI11_1/net21_12_ xsel_27_ XI11_1/XI0/XI0_27/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN0_2 XI11_1/net21_13_ xsel_27_ XI11_1/XI0/XI0_27/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN0_1 XI11_1/net21_14_ xsel_27_ XI11_1/XI0/XI0_27/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN0_0 XI11_1/net21_15_ xsel_27_ XI11_1/XI0/XI0_27/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN1_15 XI11_1/XI0/XI0_27/d__15_ xsel_27_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN1_14 XI11_1/XI0/XI0_27/d__14_ xsel_27_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN1_13 XI11_1/XI0/XI0_27/d__13_ xsel_27_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN1_12 XI11_1/XI0/XI0_27/d__12_ xsel_27_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN1_11 XI11_1/XI0/XI0_27/d__11_ xsel_27_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN1_10 XI11_1/XI0/XI0_27/d__10_ xsel_27_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN1_9 XI11_1/XI0/XI0_27/d__9_ xsel_27_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN1_8 XI11_1/XI0/XI0_27/d__8_ xsel_27_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN1_7 XI11_1/XI0/XI0_27/d__7_ xsel_27_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN1_6 XI11_1/XI0/XI0_27/d__6_ xsel_27_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN1_5 XI11_1/XI0/XI0_27/d__5_ xsel_27_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN1_4 XI11_1/XI0/XI0_27/d__4_ xsel_27_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN1_3 XI11_1/XI0/XI0_27/d__3_ xsel_27_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN1_2 XI11_1/XI0/XI0_27/d__2_ xsel_27_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN1_1 XI11_1/XI0/XI0_27/d__1_ xsel_27_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_27/MN1_0 XI11_1/XI0/XI0_27/d__0_ xsel_27_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN0_15 XI11_1/net21_0_ xsel_26_ XI11_1/XI0/XI0_26/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN0_14 XI11_1/net21_1_ xsel_26_ XI11_1/XI0/XI0_26/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN0_13 XI11_1/net21_2_ xsel_26_ XI11_1/XI0/XI0_26/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN0_12 XI11_1/net21_3_ xsel_26_ XI11_1/XI0/XI0_26/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN0_11 XI11_1/net21_4_ xsel_26_ XI11_1/XI0/XI0_26/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN0_10 XI11_1/net21_5_ xsel_26_ XI11_1/XI0/XI0_26/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN0_9 XI11_1/net21_6_ xsel_26_ XI11_1/XI0/XI0_26/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN0_8 XI11_1/net21_7_ xsel_26_ XI11_1/XI0/XI0_26/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN0_7 XI11_1/net21_8_ xsel_26_ XI11_1/XI0/XI0_26/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN0_6 XI11_1/net21_9_ xsel_26_ XI11_1/XI0/XI0_26/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN0_5 XI11_1/net21_10_ xsel_26_ XI11_1/XI0/XI0_26/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN0_4 XI11_1/net21_11_ xsel_26_ XI11_1/XI0/XI0_26/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN0_3 XI11_1/net21_12_ xsel_26_ XI11_1/XI0/XI0_26/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN0_2 XI11_1/net21_13_ xsel_26_ XI11_1/XI0/XI0_26/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN0_1 XI11_1/net21_14_ xsel_26_ XI11_1/XI0/XI0_26/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN0_0 XI11_1/net21_15_ xsel_26_ XI11_1/XI0/XI0_26/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN1_15 XI11_1/XI0/XI0_26/d__15_ xsel_26_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN1_14 XI11_1/XI0/XI0_26/d__14_ xsel_26_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN1_13 XI11_1/XI0/XI0_26/d__13_ xsel_26_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN1_12 XI11_1/XI0/XI0_26/d__12_ xsel_26_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN1_11 XI11_1/XI0/XI0_26/d__11_ xsel_26_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN1_10 XI11_1/XI0/XI0_26/d__10_ xsel_26_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN1_9 XI11_1/XI0/XI0_26/d__9_ xsel_26_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN1_8 XI11_1/XI0/XI0_26/d__8_ xsel_26_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN1_7 XI11_1/XI0/XI0_26/d__7_ xsel_26_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN1_6 XI11_1/XI0/XI0_26/d__6_ xsel_26_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN1_5 XI11_1/XI0/XI0_26/d__5_ xsel_26_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN1_4 XI11_1/XI0/XI0_26/d__4_ xsel_26_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN1_3 XI11_1/XI0/XI0_26/d__3_ xsel_26_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN1_2 XI11_1/XI0/XI0_26/d__2_ xsel_26_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN1_1 XI11_1/XI0/XI0_26/d__1_ xsel_26_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_26/MN1_0 XI11_1/XI0/XI0_26/d__0_ xsel_26_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN0_15 XI11_1/net21_0_ xsel_25_ XI11_1/XI0/XI0_25/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN0_14 XI11_1/net21_1_ xsel_25_ XI11_1/XI0/XI0_25/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN0_13 XI11_1/net21_2_ xsel_25_ XI11_1/XI0/XI0_25/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN0_12 XI11_1/net21_3_ xsel_25_ XI11_1/XI0/XI0_25/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN0_11 XI11_1/net21_4_ xsel_25_ XI11_1/XI0/XI0_25/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN0_10 XI11_1/net21_5_ xsel_25_ XI11_1/XI0/XI0_25/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN0_9 XI11_1/net21_6_ xsel_25_ XI11_1/XI0/XI0_25/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN0_8 XI11_1/net21_7_ xsel_25_ XI11_1/XI0/XI0_25/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN0_7 XI11_1/net21_8_ xsel_25_ XI11_1/XI0/XI0_25/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN0_6 XI11_1/net21_9_ xsel_25_ XI11_1/XI0/XI0_25/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN0_5 XI11_1/net21_10_ xsel_25_ XI11_1/XI0/XI0_25/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN0_4 XI11_1/net21_11_ xsel_25_ XI11_1/XI0/XI0_25/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN0_3 XI11_1/net21_12_ xsel_25_ XI11_1/XI0/XI0_25/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN0_2 XI11_1/net21_13_ xsel_25_ XI11_1/XI0/XI0_25/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN0_1 XI11_1/net21_14_ xsel_25_ XI11_1/XI0/XI0_25/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN0_0 XI11_1/net21_15_ xsel_25_ XI11_1/XI0/XI0_25/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN1_15 XI11_1/XI0/XI0_25/d__15_ xsel_25_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN1_14 XI11_1/XI0/XI0_25/d__14_ xsel_25_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN1_13 XI11_1/XI0/XI0_25/d__13_ xsel_25_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN1_12 XI11_1/XI0/XI0_25/d__12_ xsel_25_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN1_11 XI11_1/XI0/XI0_25/d__11_ xsel_25_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN1_10 XI11_1/XI0/XI0_25/d__10_ xsel_25_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN1_9 XI11_1/XI0/XI0_25/d__9_ xsel_25_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN1_8 XI11_1/XI0/XI0_25/d__8_ xsel_25_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN1_7 XI11_1/XI0/XI0_25/d__7_ xsel_25_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN1_6 XI11_1/XI0/XI0_25/d__6_ xsel_25_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN1_5 XI11_1/XI0/XI0_25/d__5_ xsel_25_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN1_4 XI11_1/XI0/XI0_25/d__4_ xsel_25_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN1_3 XI11_1/XI0/XI0_25/d__3_ xsel_25_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN1_2 XI11_1/XI0/XI0_25/d__2_ xsel_25_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN1_1 XI11_1/XI0/XI0_25/d__1_ xsel_25_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_25/MN1_0 XI11_1/XI0/XI0_25/d__0_ xsel_25_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN0_15 XI11_1/net21_0_ xsel_24_ XI11_1/XI0/XI0_24/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN0_14 XI11_1/net21_1_ xsel_24_ XI11_1/XI0/XI0_24/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN0_13 XI11_1/net21_2_ xsel_24_ XI11_1/XI0/XI0_24/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN0_12 XI11_1/net21_3_ xsel_24_ XI11_1/XI0/XI0_24/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN0_11 XI11_1/net21_4_ xsel_24_ XI11_1/XI0/XI0_24/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN0_10 XI11_1/net21_5_ xsel_24_ XI11_1/XI0/XI0_24/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN0_9 XI11_1/net21_6_ xsel_24_ XI11_1/XI0/XI0_24/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN0_8 XI11_1/net21_7_ xsel_24_ XI11_1/XI0/XI0_24/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN0_7 XI11_1/net21_8_ xsel_24_ XI11_1/XI0/XI0_24/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN0_6 XI11_1/net21_9_ xsel_24_ XI11_1/XI0/XI0_24/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN0_5 XI11_1/net21_10_ xsel_24_ XI11_1/XI0/XI0_24/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN0_4 XI11_1/net21_11_ xsel_24_ XI11_1/XI0/XI0_24/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN0_3 XI11_1/net21_12_ xsel_24_ XI11_1/XI0/XI0_24/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN0_2 XI11_1/net21_13_ xsel_24_ XI11_1/XI0/XI0_24/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN0_1 XI11_1/net21_14_ xsel_24_ XI11_1/XI0/XI0_24/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN0_0 XI11_1/net21_15_ xsel_24_ XI11_1/XI0/XI0_24/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN1_15 XI11_1/XI0/XI0_24/d__15_ xsel_24_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN1_14 XI11_1/XI0/XI0_24/d__14_ xsel_24_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN1_13 XI11_1/XI0/XI0_24/d__13_ xsel_24_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN1_12 XI11_1/XI0/XI0_24/d__12_ xsel_24_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN1_11 XI11_1/XI0/XI0_24/d__11_ xsel_24_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN1_10 XI11_1/XI0/XI0_24/d__10_ xsel_24_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN1_9 XI11_1/XI0/XI0_24/d__9_ xsel_24_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN1_8 XI11_1/XI0/XI0_24/d__8_ xsel_24_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN1_7 XI11_1/XI0/XI0_24/d__7_ xsel_24_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN1_6 XI11_1/XI0/XI0_24/d__6_ xsel_24_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN1_5 XI11_1/XI0/XI0_24/d__5_ xsel_24_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN1_4 XI11_1/XI0/XI0_24/d__4_ xsel_24_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN1_3 XI11_1/XI0/XI0_24/d__3_ xsel_24_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN1_2 XI11_1/XI0/XI0_24/d__2_ xsel_24_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN1_1 XI11_1/XI0/XI0_24/d__1_ xsel_24_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_24/MN1_0 XI11_1/XI0/XI0_24/d__0_ xsel_24_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN0_15 XI11_1/net21_0_ xsel_23_ XI11_1/XI0/XI0_23/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN0_14 XI11_1/net21_1_ xsel_23_ XI11_1/XI0/XI0_23/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN0_13 XI11_1/net21_2_ xsel_23_ XI11_1/XI0/XI0_23/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN0_12 XI11_1/net21_3_ xsel_23_ XI11_1/XI0/XI0_23/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN0_11 XI11_1/net21_4_ xsel_23_ XI11_1/XI0/XI0_23/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN0_10 XI11_1/net21_5_ xsel_23_ XI11_1/XI0/XI0_23/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN0_9 XI11_1/net21_6_ xsel_23_ XI11_1/XI0/XI0_23/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN0_8 XI11_1/net21_7_ xsel_23_ XI11_1/XI0/XI0_23/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN0_7 XI11_1/net21_8_ xsel_23_ XI11_1/XI0/XI0_23/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN0_6 XI11_1/net21_9_ xsel_23_ XI11_1/XI0/XI0_23/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN0_5 XI11_1/net21_10_ xsel_23_ XI11_1/XI0/XI0_23/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN0_4 XI11_1/net21_11_ xsel_23_ XI11_1/XI0/XI0_23/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN0_3 XI11_1/net21_12_ xsel_23_ XI11_1/XI0/XI0_23/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN0_2 XI11_1/net21_13_ xsel_23_ XI11_1/XI0/XI0_23/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN0_1 XI11_1/net21_14_ xsel_23_ XI11_1/XI0/XI0_23/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN0_0 XI11_1/net21_15_ xsel_23_ XI11_1/XI0/XI0_23/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN1_15 XI11_1/XI0/XI0_23/d__15_ xsel_23_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN1_14 XI11_1/XI0/XI0_23/d__14_ xsel_23_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN1_13 XI11_1/XI0/XI0_23/d__13_ xsel_23_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN1_12 XI11_1/XI0/XI0_23/d__12_ xsel_23_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN1_11 XI11_1/XI0/XI0_23/d__11_ xsel_23_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN1_10 XI11_1/XI0/XI0_23/d__10_ xsel_23_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN1_9 XI11_1/XI0/XI0_23/d__9_ xsel_23_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN1_8 XI11_1/XI0/XI0_23/d__8_ xsel_23_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN1_7 XI11_1/XI0/XI0_23/d__7_ xsel_23_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN1_6 XI11_1/XI0/XI0_23/d__6_ xsel_23_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN1_5 XI11_1/XI0/XI0_23/d__5_ xsel_23_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN1_4 XI11_1/XI0/XI0_23/d__4_ xsel_23_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN1_3 XI11_1/XI0/XI0_23/d__3_ xsel_23_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN1_2 XI11_1/XI0/XI0_23/d__2_ xsel_23_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN1_1 XI11_1/XI0/XI0_23/d__1_ xsel_23_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_23/MN1_0 XI11_1/XI0/XI0_23/d__0_ xsel_23_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN0_15 XI11_1/net21_0_ xsel_22_ XI11_1/XI0/XI0_22/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN0_14 XI11_1/net21_1_ xsel_22_ XI11_1/XI0/XI0_22/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN0_13 XI11_1/net21_2_ xsel_22_ XI11_1/XI0/XI0_22/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN0_12 XI11_1/net21_3_ xsel_22_ XI11_1/XI0/XI0_22/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN0_11 XI11_1/net21_4_ xsel_22_ XI11_1/XI0/XI0_22/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN0_10 XI11_1/net21_5_ xsel_22_ XI11_1/XI0/XI0_22/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN0_9 XI11_1/net21_6_ xsel_22_ XI11_1/XI0/XI0_22/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN0_8 XI11_1/net21_7_ xsel_22_ XI11_1/XI0/XI0_22/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN0_7 XI11_1/net21_8_ xsel_22_ XI11_1/XI0/XI0_22/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN0_6 XI11_1/net21_9_ xsel_22_ XI11_1/XI0/XI0_22/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN0_5 XI11_1/net21_10_ xsel_22_ XI11_1/XI0/XI0_22/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN0_4 XI11_1/net21_11_ xsel_22_ XI11_1/XI0/XI0_22/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN0_3 XI11_1/net21_12_ xsel_22_ XI11_1/XI0/XI0_22/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN0_2 XI11_1/net21_13_ xsel_22_ XI11_1/XI0/XI0_22/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN0_1 XI11_1/net21_14_ xsel_22_ XI11_1/XI0/XI0_22/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN0_0 XI11_1/net21_15_ xsel_22_ XI11_1/XI0/XI0_22/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN1_15 XI11_1/XI0/XI0_22/d__15_ xsel_22_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN1_14 XI11_1/XI0/XI0_22/d__14_ xsel_22_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN1_13 XI11_1/XI0/XI0_22/d__13_ xsel_22_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN1_12 XI11_1/XI0/XI0_22/d__12_ xsel_22_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN1_11 XI11_1/XI0/XI0_22/d__11_ xsel_22_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN1_10 XI11_1/XI0/XI0_22/d__10_ xsel_22_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN1_9 XI11_1/XI0/XI0_22/d__9_ xsel_22_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN1_8 XI11_1/XI0/XI0_22/d__8_ xsel_22_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN1_7 XI11_1/XI0/XI0_22/d__7_ xsel_22_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN1_6 XI11_1/XI0/XI0_22/d__6_ xsel_22_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN1_5 XI11_1/XI0/XI0_22/d__5_ xsel_22_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN1_4 XI11_1/XI0/XI0_22/d__4_ xsel_22_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN1_3 XI11_1/XI0/XI0_22/d__3_ xsel_22_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN1_2 XI11_1/XI0/XI0_22/d__2_ xsel_22_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN1_1 XI11_1/XI0/XI0_22/d__1_ xsel_22_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_22/MN1_0 XI11_1/XI0/XI0_22/d__0_ xsel_22_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN0_15 XI11_1/net21_0_ xsel_21_ XI11_1/XI0/XI0_21/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN0_14 XI11_1/net21_1_ xsel_21_ XI11_1/XI0/XI0_21/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN0_13 XI11_1/net21_2_ xsel_21_ XI11_1/XI0/XI0_21/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN0_12 XI11_1/net21_3_ xsel_21_ XI11_1/XI0/XI0_21/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN0_11 XI11_1/net21_4_ xsel_21_ XI11_1/XI0/XI0_21/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN0_10 XI11_1/net21_5_ xsel_21_ XI11_1/XI0/XI0_21/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN0_9 XI11_1/net21_6_ xsel_21_ XI11_1/XI0/XI0_21/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN0_8 XI11_1/net21_7_ xsel_21_ XI11_1/XI0/XI0_21/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN0_7 XI11_1/net21_8_ xsel_21_ XI11_1/XI0/XI0_21/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN0_6 XI11_1/net21_9_ xsel_21_ XI11_1/XI0/XI0_21/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN0_5 XI11_1/net21_10_ xsel_21_ XI11_1/XI0/XI0_21/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN0_4 XI11_1/net21_11_ xsel_21_ XI11_1/XI0/XI0_21/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN0_3 XI11_1/net21_12_ xsel_21_ XI11_1/XI0/XI0_21/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN0_2 XI11_1/net21_13_ xsel_21_ XI11_1/XI0/XI0_21/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN0_1 XI11_1/net21_14_ xsel_21_ XI11_1/XI0/XI0_21/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN0_0 XI11_1/net21_15_ xsel_21_ XI11_1/XI0/XI0_21/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN1_15 XI11_1/XI0/XI0_21/d__15_ xsel_21_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN1_14 XI11_1/XI0/XI0_21/d__14_ xsel_21_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN1_13 XI11_1/XI0/XI0_21/d__13_ xsel_21_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN1_12 XI11_1/XI0/XI0_21/d__12_ xsel_21_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN1_11 XI11_1/XI0/XI0_21/d__11_ xsel_21_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN1_10 XI11_1/XI0/XI0_21/d__10_ xsel_21_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN1_9 XI11_1/XI0/XI0_21/d__9_ xsel_21_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN1_8 XI11_1/XI0/XI0_21/d__8_ xsel_21_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN1_7 XI11_1/XI0/XI0_21/d__7_ xsel_21_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN1_6 XI11_1/XI0/XI0_21/d__6_ xsel_21_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN1_5 XI11_1/XI0/XI0_21/d__5_ xsel_21_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN1_4 XI11_1/XI0/XI0_21/d__4_ xsel_21_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN1_3 XI11_1/XI0/XI0_21/d__3_ xsel_21_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN1_2 XI11_1/XI0/XI0_21/d__2_ xsel_21_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN1_1 XI11_1/XI0/XI0_21/d__1_ xsel_21_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_21/MN1_0 XI11_1/XI0/XI0_21/d__0_ xsel_21_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN0_15 XI11_1/net21_0_ xsel_20_ XI11_1/XI0/XI0_20/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN0_14 XI11_1/net21_1_ xsel_20_ XI11_1/XI0/XI0_20/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN0_13 XI11_1/net21_2_ xsel_20_ XI11_1/XI0/XI0_20/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN0_12 XI11_1/net21_3_ xsel_20_ XI11_1/XI0/XI0_20/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN0_11 XI11_1/net21_4_ xsel_20_ XI11_1/XI0/XI0_20/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN0_10 XI11_1/net21_5_ xsel_20_ XI11_1/XI0/XI0_20/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN0_9 XI11_1/net21_6_ xsel_20_ XI11_1/XI0/XI0_20/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN0_8 XI11_1/net21_7_ xsel_20_ XI11_1/XI0/XI0_20/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN0_7 XI11_1/net21_8_ xsel_20_ XI11_1/XI0/XI0_20/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN0_6 XI11_1/net21_9_ xsel_20_ XI11_1/XI0/XI0_20/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN0_5 XI11_1/net21_10_ xsel_20_ XI11_1/XI0/XI0_20/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN0_4 XI11_1/net21_11_ xsel_20_ XI11_1/XI0/XI0_20/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN0_3 XI11_1/net21_12_ xsel_20_ XI11_1/XI0/XI0_20/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN0_2 XI11_1/net21_13_ xsel_20_ XI11_1/XI0/XI0_20/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN0_1 XI11_1/net21_14_ xsel_20_ XI11_1/XI0/XI0_20/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN0_0 XI11_1/net21_15_ xsel_20_ XI11_1/XI0/XI0_20/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN1_15 XI11_1/XI0/XI0_20/d__15_ xsel_20_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN1_14 XI11_1/XI0/XI0_20/d__14_ xsel_20_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN1_13 XI11_1/XI0/XI0_20/d__13_ xsel_20_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN1_12 XI11_1/XI0/XI0_20/d__12_ xsel_20_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN1_11 XI11_1/XI0/XI0_20/d__11_ xsel_20_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN1_10 XI11_1/XI0/XI0_20/d__10_ xsel_20_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN1_9 XI11_1/XI0/XI0_20/d__9_ xsel_20_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN1_8 XI11_1/XI0/XI0_20/d__8_ xsel_20_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN1_7 XI11_1/XI0/XI0_20/d__7_ xsel_20_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN1_6 XI11_1/XI0/XI0_20/d__6_ xsel_20_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN1_5 XI11_1/XI0/XI0_20/d__5_ xsel_20_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN1_4 XI11_1/XI0/XI0_20/d__4_ xsel_20_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN1_3 XI11_1/XI0/XI0_20/d__3_ xsel_20_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN1_2 XI11_1/XI0/XI0_20/d__2_ xsel_20_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN1_1 XI11_1/XI0/XI0_20/d__1_ xsel_20_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_20/MN1_0 XI11_1/XI0/XI0_20/d__0_ xsel_20_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN0_15 XI11_1/net21_0_ xsel_19_ XI11_1/XI0/XI0_19/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN0_14 XI11_1/net21_1_ xsel_19_ XI11_1/XI0/XI0_19/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN0_13 XI11_1/net21_2_ xsel_19_ XI11_1/XI0/XI0_19/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN0_12 XI11_1/net21_3_ xsel_19_ XI11_1/XI0/XI0_19/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN0_11 XI11_1/net21_4_ xsel_19_ XI11_1/XI0/XI0_19/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN0_10 XI11_1/net21_5_ xsel_19_ XI11_1/XI0/XI0_19/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN0_9 XI11_1/net21_6_ xsel_19_ XI11_1/XI0/XI0_19/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN0_8 XI11_1/net21_7_ xsel_19_ XI11_1/XI0/XI0_19/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN0_7 XI11_1/net21_8_ xsel_19_ XI11_1/XI0/XI0_19/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN0_6 XI11_1/net21_9_ xsel_19_ XI11_1/XI0/XI0_19/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN0_5 XI11_1/net21_10_ xsel_19_ XI11_1/XI0/XI0_19/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN0_4 XI11_1/net21_11_ xsel_19_ XI11_1/XI0/XI0_19/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN0_3 XI11_1/net21_12_ xsel_19_ XI11_1/XI0/XI0_19/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN0_2 XI11_1/net21_13_ xsel_19_ XI11_1/XI0/XI0_19/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN0_1 XI11_1/net21_14_ xsel_19_ XI11_1/XI0/XI0_19/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN0_0 XI11_1/net21_15_ xsel_19_ XI11_1/XI0/XI0_19/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN1_15 XI11_1/XI0/XI0_19/d__15_ xsel_19_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN1_14 XI11_1/XI0/XI0_19/d__14_ xsel_19_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN1_13 XI11_1/XI0/XI0_19/d__13_ xsel_19_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN1_12 XI11_1/XI0/XI0_19/d__12_ xsel_19_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN1_11 XI11_1/XI0/XI0_19/d__11_ xsel_19_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN1_10 XI11_1/XI0/XI0_19/d__10_ xsel_19_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN1_9 XI11_1/XI0/XI0_19/d__9_ xsel_19_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN1_8 XI11_1/XI0/XI0_19/d__8_ xsel_19_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN1_7 XI11_1/XI0/XI0_19/d__7_ xsel_19_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN1_6 XI11_1/XI0/XI0_19/d__6_ xsel_19_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN1_5 XI11_1/XI0/XI0_19/d__5_ xsel_19_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN1_4 XI11_1/XI0/XI0_19/d__4_ xsel_19_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN1_3 XI11_1/XI0/XI0_19/d__3_ xsel_19_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN1_2 XI11_1/XI0/XI0_19/d__2_ xsel_19_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN1_1 XI11_1/XI0/XI0_19/d__1_ xsel_19_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_19/MN1_0 XI11_1/XI0/XI0_19/d__0_ xsel_19_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN0_15 XI11_1/net21_0_ xsel_18_ XI11_1/XI0/XI0_18/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN0_14 XI11_1/net21_1_ xsel_18_ XI11_1/XI0/XI0_18/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN0_13 XI11_1/net21_2_ xsel_18_ XI11_1/XI0/XI0_18/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN0_12 XI11_1/net21_3_ xsel_18_ XI11_1/XI0/XI0_18/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN0_11 XI11_1/net21_4_ xsel_18_ XI11_1/XI0/XI0_18/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN0_10 XI11_1/net21_5_ xsel_18_ XI11_1/XI0/XI0_18/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN0_9 XI11_1/net21_6_ xsel_18_ XI11_1/XI0/XI0_18/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN0_8 XI11_1/net21_7_ xsel_18_ XI11_1/XI0/XI0_18/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN0_7 XI11_1/net21_8_ xsel_18_ XI11_1/XI0/XI0_18/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN0_6 XI11_1/net21_9_ xsel_18_ XI11_1/XI0/XI0_18/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN0_5 XI11_1/net21_10_ xsel_18_ XI11_1/XI0/XI0_18/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN0_4 XI11_1/net21_11_ xsel_18_ XI11_1/XI0/XI0_18/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN0_3 XI11_1/net21_12_ xsel_18_ XI11_1/XI0/XI0_18/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN0_2 XI11_1/net21_13_ xsel_18_ XI11_1/XI0/XI0_18/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN0_1 XI11_1/net21_14_ xsel_18_ XI11_1/XI0/XI0_18/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN0_0 XI11_1/net21_15_ xsel_18_ XI11_1/XI0/XI0_18/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN1_15 XI11_1/XI0/XI0_18/d__15_ xsel_18_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN1_14 XI11_1/XI0/XI0_18/d__14_ xsel_18_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN1_13 XI11_1/XI0/XI0_18/d__13_ xsel_18_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN1_12 XI11_1/XI0/XI0_18/d__12_ xsel_18_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN1_11 XI11_1/XI0/XI0_18/d__11_ xsel_18_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN1_10 XI11_1/XI0/XI0_18/d__10_ xsel_18_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN1_9 XI11_1/XI0/XI0_18/d__9_ xsel_18_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN1_8 XI11_1/XI0/XI0_18/d__8_ xsel_18_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN1_7 XI11_1/XI0/XI0_18/d__7_ xsel_18_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN1_6 XI11_1/XI0/XI0_18/d__6_ xsel_18_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN1_5 XI11_1/XI0/XI0_18/d__5_ xsel_18_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN1_4 XI11_1/XI0/XI0_18/d__4_ xsel_18_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN1_3 XI11_1/XI0/XI0_18/d__3_ xsel_18_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN1_2 XI11_1/XI0/XI0_18/d__2_ xsel_18_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN1_1 XI11_1/XI0/XI0_18/d__1_ xsel_18_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_18/MN1_0 XI11_1/XI0/XI0_18/d__0_ xsel_18_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN0_15 XI11_1/net21_0_ xsel_17_ XI11_1/XI0/XI0_17/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN0_14 XI11_1/net21_1_ xsel_17_ XI11_1/XI0/XI0_17/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN0_13 XI11_1/net21_2_ xsel_17_ XI11_1/XI0/XI0_17/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN0_12 XI11_1/net21_3_ xsel_17_ XI11_1/XI0/XI0_17/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN0_11 XI11_1/net21_4_ xsel_17_ XI11_1/XI0/XI0_17/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN0_10 XI11_1/net21_5_ xsel_17_ XI11_1/XI0/XI0_17/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN0_9 XI11_1/net21_6_ xsel_17_ XI11_1/XI0/XI0_17/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN0_8 XI11_1/net21_7_ xsel_17_ XI11_1/XI0/XI0_17/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN0_7 XI11_1/net21_8_ xsel_17_ XI11_1/XI0/XI0_17/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN0_6 XI11_1/net21_9_ xsel_17_ XI11_1/XI0/XI0_17/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN0_5 XI11_1/net21_10_ xsel_17_ XI11_1/XI0/XI0_17/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN0_4 XI11_1/net21_11_ xsel_17_ XI11_1/XI0/XI0_17/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN0_3 XI11_1/net21_12_ xsel_17_ XI11_1/XI0/XI0_17/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN0_2 XI11_1/net21_13_ xsel_17_ XI11_1/XI0/XI0_17/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN0_1 XI11_1/net21_14_ xsel_17_ XI11_1/XI0/XI0_17/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN0_0 XI11_1/net21_15_ xsel_17_ XI11_1/XI0/XI0_17/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN1_15 XI11_1/XI0/XI0_17/d__15_ xsel_17_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN1_14 XI11_1/XI0/XI0_17/d__14_ xsel_17_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN1_13 XI11_1/XI0/XI0_17/d__13_ xsel_17_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN1_12 XI11_1/XI0/XI0_17/d__12_ xsel_17_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN1_11 XI11_1/XI0/XI0_17/d__11_ xsel_17_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN1_10 XI11_1/XI0/XI0_17/d__10_ xsel_17_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN1_9 XI11_1/XI0/XI0_17/d__9_ xsel_17_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN1_8 XI11_1/XI0/XI0_17/d__8_ xsel_17_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN1_7 XI11_1/XI0/XI0_17/d__7_ xsel_17_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN1_6 XI11_1/XI0/XI0_17/d__6_ xsel_17_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN1_5 XI11_1/XI0/XI0_17/d__5_ xsel_17_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN1_4 XI11_1/XI0/XI0_17/d__4_ xsel_17_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN1_3 XI11_1/XI0/XI0_17/d__3_ xsel_17_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN1_2 XI11_1/XI0/XI0_17/d__2_ xsel_17_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN1_1 XI11_1/XI0/XI0_17/d__1_ xsel_17_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_17/MN1_0 XI11_1/XI0/XI0_17/d__0_ xsel_17_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN0_15 XI11_1/net21_0_ xsel_16_ XI11_1/XI0/XI0_16/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN0_14 XI11_1/net21_1_ xsel_16_ XI11_1/XI0/XI0_16/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN0_13 XI11_1/net21_2_ xsel_16_ XI11_1/XI0/XI0_16/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN0_12 XI11_1/net21_3_ xsel_16_ XI11_1/XI0/XI0_16/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN0_11 XI11_1/net21_4_ xsel_16_ XI11_1/XI0/XI0_16/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN0_10 XI11_1/net21_5_ xsel_16_ XI11_1/XI0/XI0_16/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN0_9 XI11_1/net21_6_ xsel_16_ XI11_1/XI0/XI0_16/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN0_8 XI11_1/net21_7_ xsel_16_ XI11_1/XI0/XI0_16/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN0_7 XI11_1/net21_8_ xsel_16_ XI11_1/XI0/XI0_16/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN0_6 XI11_1/net21_9_ xsel_16_ XI11_1/XI0/XI0_16/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN0_5 XI11_1/net21_10_ xsel_16_ XI11_1/XI0/XI0_16/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN0_4 XI11_1/net21_11_ xsel_16_ XI11_1/XI0/XI0_16/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN0_3 XI11_1/net21_12_ xsel_16_ XI11_1/XI0/XI0_16/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN0_2 XI11_1/net21_13_ xsel_16_ XI11_1/XI0/XI0_16/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN0_1 XI11_1/net21_14_ xsel_16_ XI11_1/XI0/XI0_16/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN0_0 XI11_1/net21_15_ xsel_16_ XI11_1/XI0/XI0_16/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN1_15 XI11_1/XI0/XI0_16/d__15_ xsel_16_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN1_14 XI11_1/XI0/XI0_16/d__14_ xsel_16_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN1_13 XI11_1/XI0/XI0_16/d__13_ xsel_16_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN1_12 XI11_1/XI0/XI0_16/d__12_ xsel_16_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN1_11 XI11_1/XI0/XI0_16/d__11_ xsel_16_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN1_10 XI11_1/XI0/XI0_16/d__10_ xsel_16_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN1_9 XI11_1/XI0/XI0_16/d__9_ xsel_16_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN1_8 XI11_1/XI0/XI0_16/d__8_ xsel_16_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN1_7 XI11_1/XI0/XI0_16/d__7_ xsel_16_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN1_6 XI11_1/XI0/XI0_16/d__6_ xsel_16_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN1_5 XI11_1/XI0/XI0_16/d__5_ xsel_16_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN1_4 XI11_1/XI0/XI0_16/d__4_ xsel_16_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN1_3 XI11_1/XI0/XI0_16/d__3_ xsel_16_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN1_2 XI11_1/XI0/XI0_16/d__2_ xsel_16_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN1_1 XI11_1/XI0/XI0_16/d__1_ xsel_16_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_16/MN1_0 XI11_1/XI0/XI0_16/d__0_ xsel_16_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN0_15 XI11_1/net21_0_ xsel_15_ XI11_1/XI0/XI0_15/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN0_14 XI11_1/net21_1_ xsel_15_ XI11_1/XI0/XI0_15/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN0_13 XI11_1/net21_2_ xsel_15_ XI11_1/XI0/XI0_15/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN0_12 XI11_1/net21_3_ xsel_15_ XI11_1/XI0/XI0_15/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN0_11 XI11_1/net21_4_ xsel_15_ XI11_1/XI0/XI0_15/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN0_10 XI11_1/net21_5_ xsel_15_ XI11_1/XI0/XI0_15/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN0_9 XI11_1/net21_6_ xsel_15_ XI11_1/XI0/XI0_15/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN0_8 XI11_1/net21_7_ xsel_15_ XI11_1/XI0/XI0_15/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN0_7 XI11_1/net21_8_ xsel_15_ XI11_1/XI0/XI0_15/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN0_6 XI11_1/net21_9_ xsel_15_ XI11_1/XI0/XI0_15/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN0_5 XI11_1/net21_10_ xsel_15_ XI11_1/XI0/XI0_15/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN0_4 XI11_1/net21_11_ xsel_15_ XI11_1/XI0/XI0_15/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN0_3 XI11_1/net21_12_ xsel_15_ XI11_1/XI0/XI0_15/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN0_2 XI11_1/net21_13_ xsel_15_ XI11_1/XI0/XI0_15/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN0_1 XI11_1/net21_14_ xsel_15_ XI11_1/XI0/XI0_15/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN0_0 XI11_1/net21_15_ xsel_15_ XI11_1/XI0/XI0_15/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN1_15 XI11_1/XI0/XI0_15/d__15_ xsel_15_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN1_14 XI11_1/XI0/XI0_15/d__14_ xsel_15_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN1_13 XI11_1/XI0/XI0_15/d__13_ xsel_15_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN1_12 XI11_1/XI0/XI0_15/d__12_ xsel_15_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN1_11 XI11_1/XI0/XI0_15/d__11_ xsel_15_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN1_10 XI11_1/XI0/XI0_15/d__10_ xsel_15_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN1_9 XI11_1/XI0/XI0_15/d__9_ xsel_15_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN1_8 XI11_1/XI0/XI0_15/d__8_ xsel_15_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN1_7 XI11_1/XI0/XI0_15/d__7_ xsel_15_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN1_6 XI11_1/XI0/XI0_15/d__6_ xsel_15_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN1_5 XI11_1/XI0/XI0_15/d__5_ xsel_15_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN1_4 XI11_1/XI0/XI0_15/d__4_ xsel_15_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN1_3 XI11_1/XI0/XI0_15/d__3_ xsel_15_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN1_2 XI11_1/XI0/XI0_15/d__2_ xsel_15_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN1_1 XI11_1/XI0/XI0_15/d__1_ xsel_15_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_15/MN1_0 XI11_1/XI0/XI0_15/d__0_ xsel_15_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN0_15 XI11_1/net21_0_ xsel_14_ XI11_1/XI0/XI0_14/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN0_14 XI11_1/net21_1_ xsel_14_ XI11_1/XI0/XI0_14/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN0_13 XI11_1/net21_2_ xsel_14_ XI11_1/XI0/XI0_14/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN0_12 XI11_1/net21_3_ xsel_14_ XI11_1/XI0/XI0_14/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN0_11 XI11_1/net21_4_ xsel_14_ XI11_1/XI0/XI0_14/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN0_10 XI11_1/net21_5_ xsel_14_ XI11_1/XI0/XI0_14/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN0_9 XI11_1/net21_6_ xsel_14_ XI11_1/XI0/XI0_14/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN0_8 XI11_1/net21_7_ xsel_14_ XI11_1/XI0/XI0_14/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN0_7 XI11_1/net21_8_ xsel_14_ XI11_1/XI0/XI0_14/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN0_6 XI11_1/net21_9_ xsel_14_ XI11_1/XI0/XI0_14/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN0_5 XI11_1/net21_10_ xsel_14_ XI11_1/XI0/XI0_14/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN0_4 XI11_1/net21_11_ xsel_14_ XI11_1/XI0/XI0_14/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN0_3 XI11_1/net21_12_ xsel_14_ XI11_1/XI0/XI0_14/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN0_2 XI11_1/net21_13_ xsel_14_ XI11_1/XI0/XI0_14/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN0_1 XI11_1/net21_14_ xsel_14_ XI11_1/XI0/XI0_14/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN0_0 XI11_1/net21_15_ xsel_14_ XI11_1/XI0/XI0_14/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN1_15 XI11_1/XI0/XI0_14/d__15_ xsel_14_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN1_14 XI11_1/XI0/XI0_14/d__14_ xsel_14_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN1_13 XI11_1/XI0/XI0_14/d__13_ xsel_14_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN1_12 XI11_1/XI0/XI0_14/d__12_ xsel_14_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN1_11 XI11_1/XI0/XI0_14/d__11_ xsel_14_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN1_10 XI11_1/XI0/XI0_14/d__10_ xsel_14_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN1_9 XI11_1/XI0/XI0_14/d__9_ xsel_14_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN1_8 XI11_1/XI0/XI0_14/d__8_ xsel_14_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN1_7 XI11_1/XI0/XI0_14/d__7_ xsel_14_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN1_6 XI11_1/XI0/XI0_14/d__6_ xsel_14_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN1_5 XI11_1/XI0/XI0_14/d__5_ xsel_14_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN1_4 XI11_1/XI0/XI0_14/d__4_ xsel_14_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN1_3 XI11_1/XI0/XI0_14/d__3_ xsel_14_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN1_2 XI11_1/XI0/XI0_14/d__2_ xsel_14_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN1_1 XI11_1/XI0/XI0_14/d__1_ xsel_14_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_14/MN1_0 XI11_1/XI0/XI0_14/d__0_ xsel_14_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN0_15 XI11_1/net21_0_ xsel_13_ XI11_1/XI0/XI0_13/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN0_14 XI11_1/net21_1_ xsel_13_ XI11_1/XI0/XI0_13/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN0_13 XI11_1/net21_2_ xsel_13_ XI11_1/XI0/XI0_13/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN0_12 XI11_1/net21_3_ xsel_13_ XI11_1/XI0/XI0_13/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN0_11 XI11_1/net21_4_ xsel_13_ XI11_1/XI0/XI0_13/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN0_10 XI11_1/net21_5_ xsel_13_ XI11_1/XI0/XI0_13/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN0_9 XI11_1/net21_6_ xsel_13_ XI11_1/XI0/XI0_13/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN0_8 XI11_1/net21_7_ xsel_13_ XI11_1/XI0/XI0_13/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN0_7 XI11_1/net21_8_ xsel_13_ XI11_1/XI0/XI0_13/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN0_6 XI11_1/net21_9_ xsel_13_ XI11_1/XI0/XI0_13/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN0_5 XI11_1/net21_10_ xsel_13_ XI11_1/XI0/XI0_13/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN0_4 XI11_1/net21_11_ xsel_13_ XI11_1/XI0/XI0_13/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN0_3 XI11_1/net21_12_ xsel_13_ XI11_1/XI0/XI0_13/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN0_2 XI11_1/net21_13_ xsel_13_ XI11_1/XI0/XI0_13/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN0_1 XI11_1/net21_14_ xsel_13_ XI11_1/XI0/XI0_13/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN0_0 XI11_1/net21_15_ xsel_13_ XI11_1/XI0/XI0_13/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN1_15 XI11_1/XI0/XI0_13/d__15_ xsel_13_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN1_14 XI11_1/XI0/XI0_13/d__14_ xsel_13_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN1_13 XI11_1/XI0/XI0_13/d__13_ xsel_13_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN1_12 XI11_1/XI0/XI0_13/d__12_ xsel_13_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN1_11 XI11_1/XI0/XI0_13/d__11_ xsel_13_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN1_10 XI11_1/XI0/XI0_13/d__10_ xsel_13_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN1_9 XI11_1/XI0/XI0_13/d__9_ xsel_13_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN1_8 XI11_1/XI0/XI0_13/d__8_ xsel_13_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN1_7 XI11_1/XI0/XI0_13/d__7_ xsel_13_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN1_6 XI11_1/XI0/XI0_13/d__6_ xsel_13_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN1_5 XI11_1/XI0/XI0_13/d__5_ xsel_13_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN1_4 XI11_1/XI0/XI0_13/d__4_ xsel_13_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN1_3 XI11_1/XI0/XI0_13/d__3_ xsel_13_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN1_2 XI11_1/XI0/XI0_13/d__2_ xsel_13_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN1_1 XI11_1/XI0/XI0_13/d__1_ xsel_13_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_13/MN1_0 XI11_1/XI0/XI0_13/d__0_ xsel_13_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN0_15 XI11_1/net21_0_ xsel_12_ XI11_1/XI0/XI0_12/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN0_14 XI11_1/net21_1_ xsel_12_ XI11_1/XI0/XI0_12/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN0_13 XI11_1/net21_2_ xsel_12_ XI11_1/XI0/XI0_12/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN0_12 XI11_1/net21_3_ xsel_12_ XI11_1/XI0/XI0_12/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN0_11 XI11_1/net21_4_ xsel_12_ XI11_1/XI0/XI0_12/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN0_10 XI11_1/net21_5_ xsel_12_ XI11_1/XI0/XI0_12/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN0_9 XI11_1/net21_6_ xsel_12_ XI11_1/XI0/XI0_12/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN0_8 XI11_1/net21_7_ xsel_12_ XI11_1/XI0/XI0_12/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN0_7 XI11_1/net21_8_ xsel_12_ XI11_1/XI0/XI0_12/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN0_6 XI11_1/net21_9_ xsel_12_ XI11_1/XI0/XI0_12/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN0_5 XI11_1/net21_10_ xsel_12_ XI11_1/XI0/XI0_12/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN0_4 XI11_1/net21_11_ xsel_12_ XI11_1/XI0/XI0_12/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN0_3 XI11_1/net21_12_ xsel_12_ XI11_1/XI0/XI0_12/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN0_2 XI11_1/net21_13_ xsel_12_ XI11_1/XI0/XI0_12/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN0_1 XI11_1/net21_14_ xsel_12_ XI11_1/XI0/XI0_12/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN0_0 XI11_1/net21_15_ xsel_12_ XI11_1/XI0/XI0_12/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN1_15 XI11_1/XI0/XI0_12/d__15_ xsel_12_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN1_14 XI11_1/XI0/XI0_12/d__14_ xsel_12_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN1_13 XI11_1/XI0/XI0_12/d__13_ xsel_12_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN1_12 XI11_1/XI0/XI0_12/d__12_ xsel_12_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN1_11 XI11_1/XI0/XI0_12/d__11_ xsel_12_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN1_10 XI11_1/XI0/XI0_12/d__10_ xsel_12_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN1_9 XI11_1/XI0/XI0_12/d__9_ xsel_12_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN1_8 XI11_1/XI0/XI0_12/d__8_ xsel_12_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN1_7 XI11_1/XI0/XI0_12/d__7_ xsel_12_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN1_6 XI11_1/XI0/XI0_12/d__6_ xsel_12_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN1_5 XI11_1/XI0/XI0_12/d__5_ xsel_12_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN1_4 XI11_1/XI0/XI0_12/d__4_ xsel_12_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN1_3 XI11_1/XI0/XI0_12/d__3_ xsel_12_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN1_2 XI11_1/XI0/XI0_12/d__2_ xsel_12_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN1_1 XI11_1/XI0/XI0_12/d__1_ xsel_12_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_12/MN1_0 XI11_1/XI0/XI0_12/d__0_ xsel_12_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN0_15 XI11_1/net21_0_ xsel_11_ XI11_1/XI0/XI0_11/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN0_14 XI11_1/net21_1_ xsel_11_ XI11_1/XI0/XI0_11/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN0_13 XI11_1/net21_2_ xsel_11_ XI11_1/XI0/XI0_11/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN0_12 XI11_1/net21_3_ xsel_11_ XI11_1/XI0/XI0_11/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN0_11 XI11_1/net21_4_ xsel_11_ XI11_1/XI0/XI0_11/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN0_10 XI11_1/net21_5_ xsel_11_ XI11_1/XI0/XI0_11/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN0_9 XI11_1/net21_6_ xsel_11_ XI11_1/XI0/XI0_11/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN0_8 XI11_1/net21_7_ xsel_11_ XI11_1/XI0/XI0_11/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN0_7 XI11_1/net21_8_ xsel_11_ XI11_1/XI0/XI0_11/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN0_6 XI11_1/net21_9_ xsel_11_ XI11_1/XI0/XI0_11/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN0_5 XI11_1/net21_10_ xsel_11_ XI11_1/XI0/XI0_11/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN0_4 XI11_1/net21_11_ xsel_11_ XI11_1/XI0/XI0_11/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN0_3 XI11_1/net21_12_ xsel_11_ XI11_1/XI0/XI0_11/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN0_2 XI11_1/net21_13_ xsel_11_ XI11_1/XI0/XI0_11/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN0_1 XI11_1/net21_14_ xsel_11_ XI11_1/XI0/XI0_11/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN0_0 XI11_1/net21_15_ xsel_11_ XI11_1/XI0/XI0_11/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN1_15 XI11_1/XI0/XI0_11/d__15_ xsel_11_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN1_14 XI11_1/XI0/XI0_11/d__14_ xsel_11_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN1_13 XI11_1/XI0/XI0_11/d__13_ xsel_11_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN1_12 XI11_1/XI0/XI0_11/d__12_ xsel_11_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN1_11 XI11_1/XI0/XI0_11/d__11_ xsel_11_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN1_10 XI11_1/XI0/XI0_11/d__10_ xsel_11_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN1_9 XI11_1/XI0/XI0_11/d__9_ xsel_11_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN1_8 XI11_1/XI0/XI0_11/d__8_ xsel_11_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN1_7 XI11_1/XI0/XI0_11/d__7_ xsel_11_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN1_6 XI11_1/XI0/XI0_11/d__6_ xsel_11_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN1_5 XI11_1/XI0/XI0_11/d__5_ xsel_11_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN1_4 XI11_1/XI0/XI0_11/d__4_ xsel_11_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN1_3 XI11_1/XI0/XI0_11/d__3_ xsel_11_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN1_2 XI11_1/XI0/XI0_11/d__2_ xsel_11_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN1_1 XI11_1/XI0/XI0_11/d__1_ xsel_11_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_11/MN1_0 XI11_1/XI0/XI0_11/d__0_ xsel_11_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN0_15 XI11_1/net21_0_ xsel_10_ XI11_1/XI0/XI0_10/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN0_14 XI11_1/net21_1_ xsel_10_ XI11_1/XI0/XI0_10/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN0_13 XI11_1/net21_2_ xsel_10_ XI11_1/XI0/XI0_10/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN0_12 XI11_1/net21_3_ xsel_10_ XI11_1/XI0/XI0_10/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN0_11 XI11_1/net21_4_ xsel_10_ XI11_1/XI0/XI0_10/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN0_10 XI11_1/net21_5_ xsel_10_ XI11_1/XI0/XI0_10/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN0_9 XI11_1/net21_6_ xsel_10_ XI11_1/XI0/XI0_10/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN0_8 XI11_1/net21_7_ xsel_10_ XI11_1/XI0/XI0_10/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN0_7 XI11_1/net21_8_ xsel_10_ XI11_1/XI0/XI0_10/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN0_6 XI11_1/net21_9_ xsel_10_ XI11_1/XI0/XI0_10/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN0_5 XI11_1/net21_10_ xsel_10_ XI11_1/XI0/XI0_10/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN0_4 XI11_1/net21_11_ xsel_10_ XI11_1/XI0/XI0_10/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN0_3 XI11_1/net21_12_ xsel_10_ XI11_1/XI0/XI0_10/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN0_2 XI11_1/net21_13_ xsel_10_ XI11_1/XI0/XI0_10/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN0_1 XI11_1/net21_14_ xsel_10_ XI11_1/XI0/XI0_10/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN0_0 XI11_1/net21_15_ xsel_10_ XI11_1/XI0/XI0_10/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN1_15 XI11_1/XI0/XI0_10/d__15_ xsel_10_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN1_14 XI11_1/XI0/XI0_10/d__14_ xsel_10_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN1_13 XI11_1/XI0/XI0_10/d__13_ xsel_10_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN1_12 XI11_1/XI0/XI0_10/d__12_ xsel_10_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN1_11 XI11_1/XI0/XI0_10/d__11_ xsel_10_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN1_10 XI11_1/XI0/XI0_10/d__10_ xsel_10_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN1_9 XI11_1/XI0/XI0_10/d__9_ xsel_10_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN1_8 XI11_1/XI0/XI0_10/d__8_ xsel_10_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN1_7 XI11_1/XI0/XI0_10/d__7_ xsel_10_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN1_6 XI11_1/XI0/XI0_10/d__6_ xsel_10_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN1_5 XI11_1/XI0/XI0_10/d__5_ xsel_10_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN1_4 XI11_1/XI0/XI0_10/d__4_ xsel_10_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN1_3 XI11_1/XI0/XI0_10/d__3_ xsel_10_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN1_2 XI11_1/XI0/XI0_10/d__2_ xsel_10_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN1_1 XI11_1/XI0/XI0_10/d__1_ xsel_10_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_10/MN1_0 XI11_1/XI0/XI0_10/d__0_ xsel_10_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN0_15 XI11_1/net21_0_ xsel_9_ XI11_1/XI0/XI0_9/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN0_14 XI11_1/net21_1_ xsel_9_ XI11_1/XI0/XI0_9/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN0_13 XI11_1/net21_2_ xsel_9_ XI11_1/XI0/XI0_9/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN0_12 XI11_1/net21_3_ xsel_9_ XI11_1/XI0/XI0_9/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN0_11 XI11_1/net21_4_ xsel_9_ XI11_1/XI0/XI0_9/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN0_10 XI11_1/net21_5_ xsel_9_ XI11_1/XI0/XI0_9/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN0_9 XI11_1/net21_6_ xsel_9_ XI11_1/XI0/XI0_9/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN0_8 XI11_1/net21_7_ xsel_9_ XI11_1/XI0/XI0_9/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN0_7 XI11_1/net21_8_ xsel_9_ XI11_1/XI0/XI0_9/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN0_6 XI11_1/net21_9_ xsel_9_ XI11_1/XI0/XI0_9/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN0_5 XI11_1/net21_10_ xsel_9_ XI11_1/XI0/XI0_9/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN0_4 XI11_1/net21_11_ xsel_9_ XI11_1/XI0/XI0_9/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN0_3 XI11_1/net21_12_ xsel_9_ XI11_1/XI0/XI0_9/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN0_2 XI11_1/net21_13_ xsel_9_ XI11_1/XI0/XI0_9/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN0_1 XI11_1/net21_14_ xsel_9_ XI11_1/XI0/XI0_9/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN0_0 XI11_1/net21_15_ xsel_9_ XI11_1/XI0/XI0_9/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN1_15 XI11_1/XI0/XI0_9/d__15_ xsel_9_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN1_14 XI11_1/XI0/XI0_9/d__14_ xsel_9_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN1_13 XI11_1/XI0/XI0_9/d__13_ xsel_9_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN1_12 XI11_1/XI0/XI0_9/d__12_ xsel_9_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN1_11 XI11_1/XI0/XI0_9/d__11_ xsel_9_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN1_10 XI11_1/XI0/XI0_9/d__10_ xsel_9_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN1_9 XI11_1/XI0/XI0_9/d__9_ xsel_9_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN1_8 XI11_1/XI0/XI0_9/d__8_ xsel_9_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN1_7 XI11_1/XI0/XI0_9/d__7_ xsel_9_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN1_6 XI11_1/XI0/XI0_9/d__6_ xsel_9_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN1_5 XI11_1/XI0/XI0_9/d__5_ xsel_9_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN1_4 XI11_1/XI0/XI0_9/d__4_ xsel_9_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN1_3 XI11_1/XI0/XI0_9/d__3_ xsel_9_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN1_2 XI11_1/XI0/XI0_9/d__2_ xsel_9_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN1_1 XI11_1/XI0/XI0_9/d__1_ xsel_9_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_9/MN1_0 XI11_1/XI0/XI0_9/d__0_ xsel_9_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN0_15 XI11_1/net21_0_ xsel_8_ XI11_1/XI0/XI0_8/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN0_14 XI11_1/net21_1_ xsel_8_ XI11_1/XI0/XI0_8/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN0_13 XI11_1/net21_2_ xsel_8_ XI11_1/XI0/XI0_8/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN0_12 XI11_1/net21_3_ xsel_8_ XI11_1/XI0/XI0_8/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN0_11 XI11_1/net21_4_ xsel_8_ XI11_1/XI0/XI0_8/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN0_10 XI11_1/net21_5_ xsel_8_ XI11_1/XI0/XI0_8/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN0_9 XI11_1/net21_6_ xsel_8_ XI11_1/XI0/XI0_8/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN0_8 XI11_1/net21_7_ xsel_8_ XI11_1/XI0/XI0_8/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN0_7 XI11_1/net21_8_ xsel_8_ XI11_1/XI0/XI0_8/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN0_6 XI11_1/net21_9_ xsel_8_ XI11_1/XI0/XI0_8/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN0_5 XI11_1/net21_10_ xsel_8_ XI11_1/XI0/XI0_8/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN0_4 XI11_1/net21_11_ xsel_8_ XI11_1/XI0/XI0_8/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN0_3 XI11_1/net21_12_ xsel_8_ XI11_1/XI0/XI0_8/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN0_2 XI11_1/net21_13_ xsel_8_ XI11_1/XI0/XI0_8/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN0_1 XI11_1/net21_14_ xsel_8_ XI11_1/XI0/XI0_8/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN0_0 XI11_1/net21_15_ xsel_8_ XI11_1/XI0/XI0_8/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN1_15 XI11_1/XI0/XI0_8/d__15_ xsel_8_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN1_14 XI11_1/XI0/XI0_8/d__14_ xsel_8_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN1_13 XI11_1/XI0/XI0_8/d__13_ xsel_8_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN1_12 XI11_1/XI0/XI0_8/d__12_ xsel_8_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN1_11 XI11_1/XI0/XI0_8/d__11_ xsel_8_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN1_10 XI11_1/XI0/XI0_8/d__10_ xsel_8_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN1_9 XI11_1/XI0/XI0_8/d__9_ xsel_8_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN1_8 XI11_1/XI0/XI0_8/d__8_ xsel_8_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN1_7 XI11_1/XI0/XI0_8/d__7_ xsel_8_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN1_6 XI11_1/XI0/XI0_8/d__6_ xsel_8_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN1_5 XI11_1/XI0/XI0_8/d__5_ xsel_8_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN1_4 XI11_1/XI0/XI0_8/d__4_ xsel_8_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN1_3 XI11_1/XI0/XI0_8/d__3_ xsel_8_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN1_2 XI11_1/XI0/XI0_8/d__2_ xsel_8_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN1_1 XI11_1/XI0/XI0_8/d__1_ xsel_8_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_8/MN1_0 XI11_1/XI0/XI0_8/d__0_ xsel_8_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN0_15 XI11_1/net21_0_ xsel_7_ XI11_1/XI0/XI0_7/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN0_14 XI11_1/net21_1_ xsel_7_ XI11_1/XI0/XI0_7/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN0_13 XI11_1/net21_2_ xsel_7_ XI11_1/XI0/XI0_7/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN0_12 XI11_1/net21_3_ xsel_7_ XI11_1/XI0/XI0_7/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN0_11 XI11_1/net21_4_ xsel_7_ XI11_1/XI0/XI0_7/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN0_10 XI11_1/net21_5_ xsel_7_ XI11_1/XI0/XI0_7/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN0_9 XI11_1/net21_6_ xsel_7_ XI11_1/XI0/XI0_7/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN0_8 XI11_1/net21_7_ xsel_7_ XI11_1/XI0/XI0_7/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN0_7 XI11_1/net21_8_ xsel_7_ XI11_1/XI0/XI0_7/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN0_6 XI11_1/net21_9_ xsel_7_ XI11_1/XI0/XI0_7/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN0_5 XI11_1/net21_10_ xsel_7_ XI11_1/XI0/XI0_7/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN0_4 XI11_1/net21_11_ xsel_7_ XI11_1/XI0/XI0_7/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN0_3 XI11_1/net21_12_ xsel_7_ XI11_1/XI0/XI0_7/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN0_2 XI11_1/net21_13_ xsel_7_ XI11_1/XI0/XI0_7/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN0_1 XI11_1/net21_14_ xsel_7_ XI11_1/XI0/XI0_7/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN0_0 XI11_1/net21_15_ xsel_7_ XI11_1/XI0/XI0_7/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN1_15 XI11_1/XI0/XI0_7/d__15_ xsel_7_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN1_14 XI11_1/XI0/XI0_7/d__14_ xsel_7_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN1_13 XI11_1/XI0/XI0_7/d__13_ xsel_7_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN1_12 XI11_1/XI0/XI0_7/d__12_ xsel_7_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN1_11 XI11_1/XI0/XI0_7/d__11_ xsel_7_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN1_10 XI11_1/XI0/XI0_7/d__10_ xsel_7_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN1_9 XI11_1/XI0/XI0_7/d__9_ xsel_7_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN1_8 XI11_1/XI0/XI0_7/d__8_ xsel_7_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN1_7 XI11_1/XI0/XI0_7/d__7_ xsel_7_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN1_6 XI11_1/XI0/XI0_7/d__6_ xsel_7_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN1_5 XI11_1/XI0/XI0_7/d__5_ xsel_7_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN1_4 XI11_1/XI0/XI0_7/d__4_ xsel_7_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN1_3 XI11_1/XI0/XI0_7/d__3_ xsel_7_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN1_2 XI11_1/XI0/XI0_7/d__2_ xsel_7_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN1_1 XI11_1/XI0/XI0_7/d__1_ xsel_7_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_7/MN1_0 XI11_1/XI0/XI0_7/d__0_ xsel_7_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN0_15 XI11_1/net21_0_ xsel_6_ XI11_1/XI0/XI0_6/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN0_14 XI11_1/net21_1_ xsel_6_ XI11_1/XI0/XI0_6/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN0_13 XI11_1/net21_2_ xsel_6_ XI11_1/XI0/XI0_6/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN0_12 XI11_1/net21_3_ xsel_6_ XI11_1/XI0/XI0_6/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN0_11 XI11_1/net21_4_ xsel_6_ XI11_1/XI0/XI0_6/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN0_10 XI11_1/net21_5_ xsel_6_ XI11_1/XI0/XI0_6/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN0_9 XI11_1/net21_6_ xsel_6_ XI11_1/XI0/XI0_6/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN0_8 XI11_1/net21_7_ xsel_6_ XI11_1/XI0/XI0_6/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN0_7 XI11_1/net21_8_ xsel_6_ XI11_1/XI0/XI0_6/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN0_6 XI11_1/net21_9_ xsel_6_ XI11_1/XI0/XI0_6/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN0_5 XI11_1/net21_10_ xsel_6_ XI11_1/XI0/XI0_6/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN0_4 XI11_1/net21_11_ xsel_6_ XI11_1/XI0/XI0_6/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN0_3 XI11_1/net21_12_ xsel_6_ XI11_1/XI0/XI0_6/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN0_2 XI11_1/net21_13_ xsel_6_ XI11_1/XI0/XI0_6/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN0_1 XI11_1/net21_14_ xsel_6_ XI11_1/XI0/XI0_6/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN0_0 XI11_1/net21_15_ xsel_6_ XI11_1/XI0/XI0_6/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN1_15 XI11_1/XI0/XI0_6/d__15_ xsel_6_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN1_14 XI11_1/XI0/XI0_6/d__14_ xsel_6_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN1_13 XI11_1/XI0/XI0_6/d__13_ xsel_6_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN1_12 XI11_1/XI0/XI0_6/d__12_ xsel_6_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN1_11 XI11_1/XI0/XI0_6/d__11_ xsel_6_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN1_10 XI11_1/XI0/XI0_6/d__10_ xsel_6_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN1_9 XI11_1/XI0/XI0_6/d__9_ xsel_6_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN1_8 XI11_1/XI0/XI0_6/d__8_ xsel_6_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN1_7 XI11_1/XI0/XI0_6/d__7_ xsel_6_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN1_6 XI11_1/XI0/XI0_6/d__6_ xsel_6_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN1_5 XI11_1/XI0/XI0_6/d__5_ xsel_6_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN1_4 XI11_1/XI0/XI0_6/d__4_ xsel_6_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN1_3 XI11_1/XI0/XI0_6/d__3_ xsel_6_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN1_2 XI11_1/XI0/XI0_6/d__2_ xsel_6_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN1_1 XI11_1/XI0/XI0_6/d__1_ xsel_6_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_6/MN1_0 XI11_1/XI0/XI0_6/d__0_ xsel_6_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN0_15 XI11_1/net21_0_ xsel_5_ XI11_1/XI0/XI0_5/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN0_14 XI11_1/net21_1_ xsel_5_ XI11_1/XI0/XI0_5/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN0_13 XI11_1/net21_2_ xsel_5_ XI11_1/XI0/XI0_5/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN0_12 XI11_1/net21_3_ xsel_5_ XI11_1/XI0/XI0_5/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN0_11 XI11_1/net21_4_ xsel_5_ XI11_1/XI0/XI0_5/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN0_10 XI11_1/net21_5_ xsel_5_ XI11_1/XI0/XI0_5/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN0_9 XI11_1/net21_6_ xsel_5_ XI11_1/XI0/XI0_5/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN0_8 XI11_1/net21_7_ xsel_5_ XI11_1/XI0/XI0_5/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN0_7 XI11_1/net21_8_ xsel_5_ XI11_1/XI0/XI0_5/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN0_6 XI11_1/net21_9_ xsel_5_ XI11_1/XI0/XI0_5/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN0_5 XI11_1/net21_10_ xsel_5_ XI11_1/XI0/XI0_5/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN0_4 XI11_1/net21_11_ xsel_5_ XI11_1/XI0/XI0_5/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN0_3 XI11_1/net21_12_ xsel_5_ XI11_1/XI0/XI0_5/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN0_2 XI11_1/net21_13_ xsel_5_ XI11_1/XI0/XI0_5/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN0_1 XI11_1/net21_14_ xsel_5_ XI11_1/XI0/XI0_5/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN0_0 XI11_1/net21_15_ xsel_5_ XI11_1/XI0/XI0_5/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN1_15 XI11_1/XI0/XI0_5/d__15_ xsel_5_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN1_14 XI11_1/XI0/XI0_5/d__14_ xsel_5_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN1_13 XI11_1/XI0/XI0_5/d__13_ xsel_5_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN1_12 XI11_1/XI0/XI0_5/d__12_ xsel_5_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN1_11 XI11_1/XI0/XI0_5/d__11_ xsel_5_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN1_10 XI11_1/XI0/XI0_5/d__10_ xsel_5_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN1_9 XI11_1/XI0/XI0_5/d__9_ xsel_5_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN1_8 XI11_1/XI0/XI0_5/d__8_ xsel_5_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN1_7 XI11_1/XI0/XI0_5/d__7_ xsel_5_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN1_6 XI11_1/XI0/XI0_5/d__6_ xsel_5_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN1_5 XI11_1/XI0/XI0_5/d__5_ xsel_5_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN1_4 XI11_1/XI0/XI0_5/d__4_ xsel_5_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN1_3 XI11_1/XI0/XI0_5/d__3_ xsel_5_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN1_2 XI11_1/XI0/XI0_5/d__2_ xsel_5_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN1_1 XI11_1/XI0/XI0_5/d__1_ xsel_5_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_5/MN1_0 XI11_1/XI0/XI0_5/d__0_ xsel_5_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN0_15 XI11_1/net21_0_ xsel_4_ XI11_1/XI0/XI0_4/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN0_14 XI11_1/net21_1_ xsel_4_ XI11_1/XI0/XI0_4/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN0_13 XI11_1/net21_2_ xsel_4_ XI11_1/XI0/XI0_4/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN0_12 XI11_1/net21_3_ xsel_4_ XI11_1/XI0/XI0_4/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN0_11 XI11_1/net21_4_ xsel_4_ XI11_1/XI0/XI0_4/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN0_10 XI11_1/net21_5_ xsel_4_ XI11_1/XI0/XI0_4/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN0_9 XI11_1/net21_6_ xsel_4_ XI11_1/XI0/XI0_4/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN0_8 XI11_1/net21_7_ xsel_4_ XI11_1/XI0/XI0_4/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN0_7 XI11_1/net21_8_ xsel_4_ XI11_1/XI0/XI0_4/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN0_6 XI11_1/net21_9_ xsel_4_ XI11_1/XI0/XI0_4/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN0_5 XI11_1/net21_10_ xsel_4_ XI11_1/XI0/XI0_4/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN0_4 XI11_1/net21_11_ xsel_4_ XI11_1/XI0/XI0_4/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN0_3 XI11_1/net21_12_ xsel_4_ XI11_1/XI0/XI0_4/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN0_2 XI11_1/net21_13_ xsel_4_ XI11_1/XI0/XI0_4/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN0_1 XI11_1/net21_14_ xsel_4_ XI11_1/XI0/XI0_4/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN0_0 XI11_1/net21_15_ xsel_4_ XI11_1/XI0/XI0_4/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN1_15 XI11_1/XI0/XI0_4/d__15_ xsel_4_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN1_14 XI11_1/XI0/XI0_4/d__14_ xsel_4_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN1_13 XI11_1/XI0/XI0_4/d__13_ xsel_4_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN1_12 XI11_1/XI0/XI0_4/d__12_ xsel_4_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN1_11 XI11_1/XI0/XI0_4/d__11_ xsel_4_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN1_10 XI11_1/XI0/XI0_4/d__10_ xsel_4_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN1_9 XI11_1/XI0/XI0_4/d__9_ xsel_4_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN1_8 XI11_1/XI0/XI0_4/d__8_ xsel_4_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN1_7 XI11_1/XI0/XI0_4/d__7_ xsel_4_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN1_6 XI11_1/XI0/XI0_4/d__6_ xsel_4_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN1_5 XI11_1/XI0/XI0_4/d__5_ xsel_4_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN1_4 XI11_1/XI0/XI0_4/d__4_ xsel_4_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN1_3 XI11_1/XI0/XI0_4/d__3_ xsel_4_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN1_2 XI11_1/XI0/XI0_4/d__2_ xsel_4_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN1_1 XI11_1/XI0/XI0_4/d__1_ xsel_4_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_4/MN1_0 XI11_1/XI0/XI0_4/d__0_ xsel_4_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN0_15 XI11_1/net21_0_ xsel_3_ XI11_1/XI0/XI0_3/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN0_14 XI11_1/net21_1_ xsel_3_ XI11_1/XI0/XI0_3/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN0_13 XI11_1/net21_2_ xsel_3_ XI11_1/XI0/XI0_3/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN0_12 XI11_1/net21_3_ xsel_3_ XI11_1/XI0/XI0_3/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN0_11 XI11_1/net21_4_ xsel_3_ XI11_1/XI0/XI0_3/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN0_10 XI11_1/net21_5_ xsel_3_ XI11_1/XI0/XI0_3/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN0_9 XI11_1/net21_6_ xsel_3_ XI11_1/XI0/XI0_3/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN0_8 XI11_1/net21_7_ xsel_3_ XI11_1/XI0/XI0_3/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN0_7 XI11_1/net21_8_ xsel_3_ XI11_1/XI0/XI0_3/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN0_6 XI11_1/net21_9_ xsel_3_ XI11_1/XI0/XI0_3/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN0_5 XI11_1/net21_10_ xsel_3_ XI11_1/XI0/XI0_3/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN0_4 XI11_1/net21_11_ xsel_3_ XI11_1/XI0/XI0_3/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN0_3 XI11_1/net21_12_ xsel_3_ XI11_1/XI0/XI0_3/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN0_2 XI11_1/net21_13_ xsel_3_ XI11_1/XI0/XI0_3/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN0_1 XI11_1/net21_14_ xsel_3_ XI11_1/XI0/XI0_3/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN0_0 XI11_1/net21_15_ xsel_3_ XI11_1/XI0/XI0_3/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN1_15 XI11_1/XI0/XI0_3/d__15_ xsel_3_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN1_14 XI11_1/XI0/XI0_3/d__14_ xsel_3_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN1_13 XI11_1/XI0/XI0_3/d__13_ xsel_3_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN1_12 XI11_1/XI0/XI0_3/d__12_ xsel_3_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN1_11 XI11_1/XI0/XI0_3/d__11_ xsel_3_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN1_10 XI11_1/XI0/XI0_3/d__10_ xsel_3_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN1_9 XI11_1/XI0/XI0_3/d__9_ xsel_3_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN1_8 XI11_1/XI0/XI0_3/d__8_ xsel_3_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN1_7 XI11_1/XI0/XI0_3/d__7_ xsel_3_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN1_6 XI11_1/XI0/XI0_3/d__6_ xsel_3_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN1_5 XI11_1/XI0/XI0_3/d__5_ xsel_3_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN1_4 XI11_1/XI0/XI0_3/d__4_ xsel_3_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN1_3 XI11_1/XI0/XI0_3/d__3_ xsel_3_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN1_2 XI11_1/XI0/XI0_3/d__2_ xsel_3_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN1_1 XI11_1/XI0/XI0_3/d__1_ xsel_3_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_3/MN1_0 XI11_1/XI0/XI0_3/d__0_ xsel_3_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN0_15 XI11_1/net21_0_ xsel_2_ XI11_1/XI0/XI0_2/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN0_14 XI11_1/net21_1_ xsel_2_ XI11_1/XI0/XI0_2/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN0_13 XI11_1/net21_2_ xsel_2_ XI11_1/XI0/XI0_2/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN0_12 XI11_1/net21_3_ xsel_2_ XI11_1/XI0/XI0_2/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN0_11 XI11_1/net21_4_ xsel_2_ XI11_1/XI0/XI0_2/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN0_10 XI11_1/net21_5_ xsel_2_ XI11_1/XI0/XI0_2/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN0_9 XI11_1/net21_6_ xsel_2_ XI11_1/XI0/XI0_2/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN0_8 XI11_1/net21_7_ xsel_2_ XI11_1/XI0/XI0_2/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN0_7 XI11_1/net21_8_ xsel_2_ XI11_1/XI0/XI0_2/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN0_6 XI11_1/net21_9_ xsel_2_ XI11_1/XI0/XI0_2/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN0_5 XI11_1/net21_10_ xsel_2_ XI11_1/XI0/XI0_2/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN0_4 XI11_1/net21_11_ xsel_2_ XI11_1/XI0/XI0_2/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN0_3 XI11_1/net21_12_ xsel_2_ XI11_1/XI0/XI0_2/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN0_2 XI11_1/net21_13_ xsel_2_ XI11_1/XI0/XI0_2/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN0_1 XI11_1/net21_14_ xsel_2_ XI11_1/XI0/XI0_2/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN0_0 XI11_1/net21_15_ xsel_2_ XI11_1/XI0/XI0_2/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN1_15 XI11_1/XI0/XI0_2/d__15_ xsel_2_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN1_14 XI11_1/XI0/XI0_2/d__14_ xsel_2_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN1_13 XI11_1/XI0/XI0_2/d__13_ xsel_2_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN1_12 XI11_1/XI0/XI0_2/d__12_ xsel_2_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN1_11 XI11_1/XI0/XI0_2/d__11_ xsel_2_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN1_10 XI11_1/XI0/XI0_2/d__10_ xsel_2_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN1_9 XI11_1/XI0/XI0_2/d__9_ xsel_2_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN1_8 XI11_1/XI0/XI0_2/d__8_ xsel_2_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN1_7 XI11_1/XI0/XI0_2/d__7_ xsel_2_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN1_6 XI11_1/XI0/XI0_2/d__6_ xsel_2_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN1_5 XI11_1/XI0/XI0_2/d__5_ xsel_2_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN1_4 XI11_1/XI0/XI0_2/d__4_ xsel_2_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN1_3 XI11_1/XI0/XI0_2/d__3_ xsel_2_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN1_2 XI11_1/XI0/XI0_2/d__2_ xsel_2_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN1_1 XI11_1/XI0/XI0_2/d__1_ xsel_2_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_2/MN1_0 XI11_1/XI0/XI0_2/d__0_ xsel_2_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN0_15 XI11_1/net21_0_ xsel_1_ XI11_1/XI0/XI0_1/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN0_14 XI11_1/net21_1_ xsel_1_ XI11_1/XI0/XI0_1/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN0_13 XI11_1/net21_2_ xsel_1_ XI11_1/XI0/XI0_1/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN0_12 XI11_1/net21_3_ xsel_1_ XI11_1/XI0/XI0_1/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN0_11 XI11_1/net21_4_ xsel_1_ XI11_1/XI0/XI0_1/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN0_10 XI11_1/net21_5_ xsel_1_ XI11_1/XI0/XI0_1/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN0_9 XI11_1/net21_6_ xsel_1_ XI11_1/XI0/XI0_1/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN0_8 XI11_1/net21_7_ xsel_1_ XI11_1/XI0/XI0_1/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN0_7 XI11_1/net21_8_ xsel_1_ XI11_1/XI0/XI0_1/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN0_6 XI11_1/net21_9_ xsel_1_ XI11_1/XI0/XI0_1/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN0_5 XI11_1/net21_10_ xsel_1_ XI11_1/XI0/XI0_1/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN0_4 XI11_1/net21_11_ xsel_1_ XI11_1/XI0/XI0_1/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN0_3 XI11_1/net21_12_ xsel_1_ XI11_1/XI0/XI0_1/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN0_2 XI11_1/net21_13_ xsel_1_ XI11_1/XI0/XI0_1/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN0_1 XI11_1/net21_14_ xsel_1_ XI11_1/XI0/XI0_1/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN0_0 XI11_1/net21_15_ xsel_1_ XI11_1/XI0/XI0_1/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN1_15 XI11_1/XI0/XI0_1/d__15_ xsel_1_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN1_14 XI11_1/XI0/XI0_1/d__14_ xsel_1_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN1_13 XI11_1/XI0/XI0_1/d__13_ xsel_1_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN1_12 XI11_1/XI0/XI0_1/d__12_ xsel_1_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN1_11 XI11_1/XI0/XI0_1/d__11_ xsel_1_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN1_10 XI11_1/XI0/XI0_1/d__10_ xsel_1_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN1_9 XI11_1/XI0/XI0_1/d__9_ xsel_1_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN1_8 XI11_1/XI0/XI0_1/d__8_ xsel_1_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN1_7 XI11_1/XI0/XI0_1/d__7_ xsel_1_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN1_6 XI11_1/XI0/XI0_1/d__6_ xsel_1_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN1_5 XI11_1/XI0/XI0_1/d__5_ xsel_1_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN1_4 XI11_1/XI0/XI0_1/d__4_ xsel_1_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN1_3 XI11_1/XI0/XI0_1/d__3_ xsel_1_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN1_2 XI11_1/XI0/XI0_1/d__2_ xsel_1_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN1_1 XI11_1/XI0/XI0_1/d__1_ xsel_1_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_1/MN1_0 XI11_1/XI0/XI0_1/d__0_ xsel_1_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN0_15 XI11_1/net21_0_ xsel_0_ XI11_1/XI0/XI0_0/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN0_14 XI11_1/net21_1_ xsel_0_ XI11_1/XI0/XI0_0/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN0_13 XI11_1/net21_2_ xsel_0_ XI11_1/XI0/XI0_0/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN0_12 XI11_1/net21_3_ xsel_0_ XI11_1/XI0/XI0_0/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN0_11 XI11_1/net21_4_ xsel_0_ XI11_1/XI0/XI0_0/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN0_10 XI11_1/net21_5_ xsel_0_ XI11_1/XI0/XI0_0/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN0_9 XI11_1/net21_6_ xsel_0_ XI11_1/XI0/XI0_0/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN0_8 XI11_1/net21_7_ xsel_0_ XI11_1/XI0/XI0_0/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN0_7 XI11_1/net21_8_ xsel_0_ XI11_1/XI0/XI0_0/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN0_6 XI11_1/net21_9_ xsel_0_ XI11_1/XI0/XI0_0/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN0_5 XI11_1/net21_10_ xsel_0_ XI11_1/XI0/XI0_0/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN0_4 XI11_1/net21_11_ xsel_0_ XI11_1/XI0/XI0_0/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN0_3 XI11_1/net21_12_ xsel_0_ XI11_1/XI0/XI0_0/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN0_2 XI11_1/net21_13_ xsel_0_ XI11_1/XI0/XI0_0/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN0_1 XI11_1/net21_14_ xsel_0_ XI11_1/XI0/XI0_0/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN0_0 XI11_1/net21_15_ xsel_0_ XI11_1/XI0/XI0_0/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN1_15 XI11_1/XI0/XI0_0/d__15_ xsel_0_ XI11_1/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN1_14 XI11_1/XI0/XI0_0/d__14_ xsel_0_ XI11_1/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN1_13 XI11_1/XI0/XI0_0/d__13_ xsel_0_ XI11_1/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN1_12 XI11_1/XI0/XI0_0/d__12_ xsel_0_ XI11_1/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN1_11 XI11_1/XI0/XI0_0/d__11_ xsel_0_ XI11_1/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN1_10 XI11_1/XI0/XI0_0/d__10_ xsel_0_ XI11_1/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN1_9 XI11_1/XI0/XI0_0/d__9_ xsel_0_ XI11_1/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN1_8 XI11_1/XI0/XI0_0/d__8_ xsel_0_ XI11_1/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN1_7 XI11_1/XI0/XI0_0/d__7_ xsel_0_ XI11_1/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN1_6 XI11_1/XI0/XI0_0/d__6_ xsel_0_ XI11_1/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN1_5 XI11_1/XI0/XI0_0/d__5_ xsel_0_ XI11_1/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN1_4 XI11_1/XI0/XI0_0/d__4_ xsel_0_ XI11_1/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN1_3 XI11_1/XI0/XI0_0/d__3_ xsel_0_ XI11_1/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN1_2 XI11_1/XI0/XI0_0/d__2_ xsel_0_ XI11_1/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN1_1 XI11_1/XI0/XI0_0/d__1_ xsel_0_ XI11_1/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_1/XI0/XI0_0/MN1_0 XI11_1/XI0/XI0_0/d__0_ xsel_0_ XI11_1/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI2/MN0_15 XI11_0/net21_0_ ysel_15_ XI11_0/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN0_14 XI11_0/net21_1_ ysel_14_ XI11_0/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN0_13 XI11_0/net21_2_ ysel_13_ XI11_0/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN0_12 XI11_0/net21_3_ ysel_12_ XI11_0/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN0_11 XI11_0/net21_4_ ysel_11_ XI11_0/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN0_10 XI11_0/net21_5_ ysel_10_ XI11_0/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN0_9 XI11_0/net21_6_ ysel_9_ XI11_0/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN0_8 XI11_0/net21_7_ ysel_8_ XI11_0/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN0_7 XI11_0/net21_8_ ysel_7_ XI11_0/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN0_6 XI11_0/net21_9_ ysel_6_ XI11_0/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN0_5 XI11_0/net21_10_ ysel_5_ XI11_0/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN0_4 XI11_0/net21_11_ ysel_4_ XI11_0/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN0_3 XI11_0/net21_12_ ysel_3_ XI11_0/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN0_2 XI11_0/net21_13_ ysel_2_ XI11_0/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN0_1 XI11_0/net21_14_ ysel_1_ XI11_0/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN0_0 XI11_0/net21_15_ ysel_0_ XI11_0/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN1_15 XI11_0/net20_0_ ysel_15_ XI11_0/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN1_14 XI11_0/net20_1_ ysel_14_ XI11_0/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN1_13 XI11_0/net20_2_ ysel_13_ XI11_0/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN1_12 XI11_0/net20_3_ ysel_12_ XI11_0/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN1_11 XI11_0/net20_4_ ysel_11_ XI11_0/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN1_10 XI11_0/net20_5_ ysel_10_ XI11_0/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN1_9 XI11_0/net20_6_ ysel_9_ XI11_0/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN1_8 XI11_0/net20_7_ ysel_8_ XI11_0/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN1_7 XI11_0/net20_8_ ysel_7_ XI11_0/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN1_6 XI11_0/net20_9_ ysel_6_ XI11_0/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN1_5 XI11_0/net20_10_ ysel_5_ XI11_0/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN1_4 XI11_0/net20_11_ ysel_4_ XI11_0/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN1_3 XI11_0/net20_12_ ysel_3_ XI11_0/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN1_2 XI11_0/net20_13_ ysel_2_ XI11_0/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN1_1 XI11_0/net20_14_ ysel_1_ XI11_0/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI2/MN1_0 XI11_0/net20_15_ ysel_0_ XI11_0/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_0/XI4/MN8 vdd XI11_0/XI4/net8 XI11_0/net12 vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_0/XI4/MP0 XI11_0/net9 XI11_0/XI4/net23 vdd vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_0/XI4/MP4 XI11_0/net12 XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI4/MP1 XI11_0/net9 XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI4/MP5 XI11_0/net12 XI11_0/preck XI11_0/net9 vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI4/MN7 vdd XI11_0/XI4/net090 DOUT_0_ vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_0/XI4/MP3 gnd XI11_0/XI4/net089 XI11_0/net12 gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_0/XI4/MN5 XI11_0/net9 XI11_0/XI4/net0103 gnd gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_0/XI4/MN4 XI11_0/XI4/data_out_ XI11_0/XI4/net32 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_0/XI4/MN0 XI11_0/XI4/data_out XI11_0/XI4/net52 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_0/XI4/MN9 gnd XI11_0/XI4/net0112 DOUT_0_ gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_0/XI1_15/MP2 XI11_0/net20_0_ XI11_0/preck XI11_0/net21_0_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI1_15/MP1 XI11_0/net20_0_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_15/MP0 XI11_0/net21_0_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_14/MP2 XI11_0/net20_1_ XI11_0/preck XI11_0/net21_1_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI1_14/MP1 XI11_0/net20_1_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_14/MP0 XI11_0/net21_1_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_13/MP2 XI11_0/net20_2_ XI11_0/preck XI11_0/net21_2_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI1_13/MP1 XI11_0/net20_2_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_13/MP0 XI11_0/net21_2_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_12/MP2 XI11_0/net20_3_ XI11_0/preck XI11_0/net21_3_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI1_12/MP1 XI11_0/net20_3_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_12/MP0 XI11_0/net21_3_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_11/MP2 XI11_0/net20_4_ XI11_0/preck XI11_0/net21_4_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI1_11/MP1 XI11_0/net20_4_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_11/MP0 XI11_0/net21_4_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_10/MP2 XI11_0/net20_5_ XI11_0/preck XI11_0/net21_5_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI1_10/MP1 XI11_0/net20_5_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_10/MP0 XI11_0/net21_5_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_9/MP2 XI11_0/net20_6_ XI11_0/preck XI11_0/net21_6_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI1_9/MP1 XI11_0/net20_6_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_9/MP0 XI11_0/net21_6_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_8/MP2 XI11_0/net20_7_ XI11_0/preck XI11_0/net21_7_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI1_8/MP1 XI11_0/net20_7_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_8/MP0 XI11_0/net21_7_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_7/MP2 XI11_0/net20_8_ XI11_0/preck XI11_0/net21_8_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI1_7/MP1 XI11_0/net20_8_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_7/MP0 XI11_0/net21_8_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_6/MP2 XI11_0/net20_9_ XI11_0/preck XI11_0/net21_9_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI1_6/MP1 XI11_0/net20_9_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_6/MP0 XI11_0/net21_9_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_5/MP2 XI11_0/net20_10_ XI11_0/preck XI11_0/net21_10_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI1_5/MP1 XI11_0/net20_10_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_5/MP0 XI11_0/net21_10_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_4/MP2 XI11_0/net20_11_ XI11_0/preck XI11_0/net21_11_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI1_4/MP1 XI11_0/net20_11_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_4/MP0 XI11_0/net21_11_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_3/MP2 XI11_0/net20_12_ XI11_0/preck XI11_0/net21_12_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI1_3/MP1 XI11_0/net20_12_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_3/MP0 XI11_0/net21_12_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_2/MP2 XI11_0/net20_13_ XI11_0/preck XI11_0/net21_13_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI1_2/MP1 XI11_0/net20_13_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_2/MP0 XI11_0/net21_13_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_1/MP2 XI11_0/net20_14_ XI11_0/preck XI11_0/net21_14_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI1_1/MP1 XI11_0/net20_14_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_1/MP0 XI11_0/net21_14_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_0/MP2 XI11_0/net20_15_ XI11_0/preck XI11_0/net21_15_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_0/XI1_0/MP1 XI11_0/net20_15_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI1_0/MP0 XI11_0/net21_15_ XI11_0/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_0/XI0/MN0_15 gnd gnd XI11_0/net21_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN0_14 gnd gnd XI11_0/net21_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN0_13 gnd gnd XI11_0/net21_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN0_12 gnd gnd XI11_0/net21_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN0_11 gnd gnd XI11_0/net21_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN0_10 gnd gnd XI11_0/net21_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN0_9 gnd gnd XI11_0/net21_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN0_8 gnd gnd XI11_0/net21_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN0_7 gnd gnd XI11_0/net21_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN0_6 gnd gnd XI11_0/net21_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN0_5 gnd gnd XI11_0/net21_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN0_4 gnd gnd XI11_0/net21_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN0_3 gnd gnd XI11_0/net21_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN0_2 gnd gnd XI11_0/net21_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN0_1 gnd gnd XI11_0/net21_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN0_0 gnd gnd XI11_0/net21_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN1_15 gnd gnd XI11_0/net20_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN1_14 gnd gnd XI11_0/net20_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN1_13 gnd gnd XI11_0/net20_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN1_12 gnd gnd XI11_0/net20_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN1_11 gnd gnd XI11_0/net20_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN1_10 gnd gnd XI11_0/net20_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN1_9 gnd gnd XI11_0/net20_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN1_8 gnd gnd XI11_0/net20_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN1_7 gnd gnd XI11_0/net20_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN1_6 gnd gnd XI11_0/net20_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN1_5 gnd gnd XI11_0/net20_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN1_4 gnd gnd XI11_0/net20_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN1_3 gnd gnd XI11_0/net20_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN1_2 gnd gnd XI11_0/net20_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN1_1 gnd gnd XI11_0/net20_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/MN1_0 gnd gnd XI11_0/net20_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN0_15 XI11_0/net21_0_ xsel_63_ XI11_0/XI0/XI0_63/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN0_14 XI11_0/net21_1_ xsel_63_ XI11_0/XI0/XI0_63/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN0_13 XI11_0/net21_2_ xsel_63_ XI11_0/XI0/XI0_63/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN0_12 XI11_0/net21_3_ xsel_63_ XI11_0/XI0/XI0_63/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN0_11 XI11_0/net21_4_ xsel_63_ XI11_0/XI0/XI0_63/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN0_10 XI11_0/net21_5_ xsel_63_ XI11_0/XI0/XI0_63/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN0_9 XI11_0/net21_6_ xsel_63_ XI11_0/XI0/XI0_63/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN0_8 XI11_0/net21_7_ xsel_63_ XI11_0/XI0/XI0_63/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN0_7 XI11_0/net21_8_ xsel_63_ XI11_0/XI0/XI0_63/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN0_6 XI11_0/net21_9_ xsel_63_ XI11_0/XI0/XI0_63/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN0_5 XI11_0/net21_10_ xsel_63_ XI11_0/XI0/XI0_63/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN0_4 XI11_0/net21_11_ xsel_63_ XI11_0/XI0/XI0_63/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN0_3 XI11_0/net21_12_ xsel_63_ XI11_0/XI0/XI0_63/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN0_2 XI11_0/net21_13_ xsel_63_ XI11_0/XI0/XI0_63/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN0_1 XI11_0/net21_14_ xsel_63_ XI11_0/XI0/XI0_63/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN0_0 XI11_0/net21_15_ xsel_63_ XI11_0/XI0/XI0_63/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN1_15 XI11_0/XI0/XI0_63/d__15_ xsel_63_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN1_14 XI11_0/XI0/XI0_63/d__14_ xsel_63_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN1_13 XI11_0/XI0/XI0_63/d__13_ xsel_63_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN1_12 XI11_0/XI0/XI0_63/d__12_ xsel_63_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN1_11 XI11_0/XI0/XI0_63/d__11_ xsel_63_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN1_10 XI11_0/XI0/XI0_63/d__10_ xsel_63_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN1_9 XI11_0/XI0/XI0_63/d__9_ xsel_63_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN1_8 XI11_0/XI0/XI0_63/d__8_ xsel_63_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN1_7 XI11_0/XI0/XI0_63/d__7_ xsel_63_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN1_6 XI11_0/XI0/XI0_63/d__6_ xsel_63_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN1_5 XI11_0/XI0/XI0_63/d__5_ xsel_63_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN1_4 XI11_0/XI0/XI0_63/d__4_ xsel_63_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN1_3 XI11_0/XI0/XI0_63/d__3_ xsel_63_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN1_2 XI11_0/XI0/XI0_63/d__2_ xsel_63_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN1_1 XI11_0/XI0/XI0_63/d__1_ xsel_63_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_63/MN1_0 XI11_0/XI0/XI0_63/d__0_ xsel_63_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN0_15 XI11_0/net21_0_ xsel_62_ XI11_0/XI0/XI0_62/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN0_14 XI11_0/net21_1_ xsel_62_ XI11_0/XI0/XI0_62/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN0_13 XI11_0/net21_2_ xsel_62_ XI11_0/XI0/XI0_62/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN0_12 XI11_0/net21_3_ xsel_62_ XI11_0/XI0/XI0_62/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN0_11 XI11_0/net21_4_ xsel_62_ XI11_0/XI0/XI0_62/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN0_10 XI11_0/net21_5_ xsel_62_ XI11_0/XI0/XI0_62/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN0_9 XI11_0/net21_6_ xsel_62_ XI11_0/XI0/XI0_62/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN0_8 XI11_0/net21_7_ xsel_62_ XI11_0/XI0/XI0_62/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN0_7 XI11_0/net21_8_ xsel_62_ XI11_0/XI0/XI0_62/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN0_6 XI11_0/net21_9_ xsel_62_ XI11_0/XI0/XI0_62/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN0_5 XI11_0/net21_10_ xsel_62_ XI11_0/XI0/XI0_62/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN0_4 XI11_0/net21_11_ xsel_62_ XI11_0/XI0/XI0_62/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN0_3 XI11_0/net21_12_ xsel_62_ XI11_0/XI0/XI0_62/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN0_2 XI11_0/net21_13_ xsel_62_ XI11_0/XI0/XI0_62/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN0_1 XI11_0/net21_14_ xsel_62_ XI11_0/XI0/XI0_62/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN0_0 XI11_0/net21_15_ xsel_62_ XI11_0/XI0/XI0_62/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN1_15 XI11_0/XI0/XI0_62/d__15_ xsel_62_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN1_14 XI11_0/XI0/XI0_62/d__14_ xsel_62_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN1_13 XI11_0/XI0/XI0_62/d__13_ xsel_62_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN1_12 XI11_0/XI0/XI0_62/d__12_ xsel_62_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN1_11 XI11_0/XI0/XI0_62/d__11_ xsel_62_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN1_10 XI11_0/XI0/XI0_62/d__10_ xsel_62_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN1_9 XI11_0/XI0/XI0_62/d__9_ xsel_62_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN1_8 XI11_0/XI0/XI0_62/d__8_ xsel_62_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN1_7 XI11_0/XI0/XI0_62/d__7_ xsel_62_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN1_6 XI11_0/XI0/XI0_62/d__6_ xsel_62_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN1_5 XI11_0/XI0/XI0_62/d__5_ xsel_62_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN1_4 XI11_0/XI0/XI0_62/d__4_ xsel_62_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN1_3 XI11_0/XI0/XI0_62/d__3_ xsel_62_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN1_2 XI11_0/XI0/XI0_62/d__2_ xsel_62_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN1_1 XI11_0/XI0/XI0_62/d__1_ xsel_62_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_62/MN1_0 XI11_0/XI0/XI0_62/d__0_ xsel_62_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN0_15 XI11_0/net21_0_ xsel_61_ XI11_0/XI0/XI0_61/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN0_14 XI11_0/net21_1_ xsel_61_ XI11_0/XI0/XI0_61/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN0_13 XI11_0/net21_2_ xsel_61_ XI11_0/XI0/XI0_61/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN0_12 XI11_0/net21_3_ xsel_61_ XI11_0/XI0/XI0_61/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN0_11 XI11_0/net21_4_ xsel_61_ XI11_0/XI0/XI0_61/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN0_10 XI11_0/net21_5_ xsel_61_ XI11_0/XI0/XI0_61/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN0_9 XI11_0/net21_6_ xsel_61_ XI11_0/XI0/XI0_61/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN0_8 XI11_0/net21_7_ xsel_61_ XI11_0/XI0/XI0_61/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN0_7 XI11_0/net21_8_ xsel_61_ XI11_0/XI0/XI0_61/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN0_6 XI11_0/net21_9_ xsel_61_ XI11_0/XI0/XI0_61/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN0_5 XI11_0/net21_10_ xsel_61_ XI11_0/XI0/XI0_61/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN0_4 XI11_0/net21_11_ xsel_61_ XI11_0/XI0/XI0_61/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN0_3 XI11_0/net21_12_ xsel_61_ XI11_0/XI0/XI0_61/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN0_2 XI11_0/net21_13_ xsel_61_ XI11_0/XI0/XI0_61/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN0_1 XI11_0/net21_14_ xsel_61_ XI11_0/XI0/XI0_61/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN0_0 XI11_0/net21_15_ xsel_61_ XI11_0/XI0/XI0_61/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN1_15 XI11_0/XI0/XI0_61/d__15_ xsel_61_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN1_14 XI11_0/XI0/XI0_61/d__14_ xsel_61_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN1_13 XI11_0/XI0/XI0_61/d__13_ xsel_61_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN1_12 XI11_0/XI0/XI0_61/d__12_ xsel_61_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN1_11 XI11_0/XI0/XI0_61/d__11_ xsel_61_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN1_10 XI11_0/XI0/XI0_61/d__10_ xsel_61_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN1_9 XI11_0/XI0/XI0_61/d__9_ xsel_61_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN1_8 XI11_0/XI0/XI0_61/d__8_ xsel_61_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN1_7 XI11_0/XI0/XI0_61/d__7_ xsel_61_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN1_6 XI11_0/XI0/XI0_61/d__6_ xsel_61_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN1_5 XI11_0/XI0/XI0_61/d__5_ xsel_61_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN1_4 XI11_0/XI0/XI0_61/d__4_ xsel_61_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN1_3 XI11_0/XI0/XI0_61/d__3_ xsel_61_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN1_2 XI11_0/XI0/XI0_61/d__2_ xsel_61_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN1_1 XI11_0/XI0/XI0_61/d__1_ xsel_61_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_61/MN1_0 XI11_0/XI0/XI0_61/d__0_ xsel_61_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN0_15 XI11_0/net21_0_ xsel_60_ XI11_0/XI0/XI0_60/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN0_14 XI11_0/net21_1_ xsel_60_ XI11_0/XI0/XI0_60/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN0_13 XI11_0/net21_2_ xsel_60_ XI11_0/XI0/XI0_60/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN0_12 XI11_0/net21_3_ xsel_60_ XI11_0/XI0/XI0_60/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN0_11 XI11_0/net21_4_ xsel_60_ XI11_0/XI0/XI0_60/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN0_10 XI11_0/net21_5_ xsel_60_ XI11_0/XI0/XI0_60/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN0_9 XI11_0/net21_6_ xsel_60_ XI11_0/XI0/XI0_60/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN0_8 XI11_0/net21_7_ xsel_60_ XI11_0/XI0/XI0_60/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN0_7 XI11_0/net21_8_ xsel_60_ XI11_0/XI0/XI0_60/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN0_6 XI11_0/net21_9_ xsel_60_ XI11_0/XI0/XI0_60/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN0_5 XI11_0/net21_10_ xsel_60_ XI11_0/XI0/XI0_60/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN0_4 XI11_0/net21_11_ xsel_60_ XI11_0/XI0/XI0_60/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN0_3 XI11_0/net21_12_ xsel_60_ XI11_0/XI0/XI0_60/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN0_2 XI11_0/net21_13_ xsel_60_ XI11_0/XI0/XI0_60/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN0_1 XI11_0/net21_14_ xsel_60_ XI11_0/XI0/XI0_60/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN0_0 XI11_0/net21_15_ xsel_60_ XI11_0/XI0/XI0_60/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN1_15 XI11_0/XI0/XI0_60/d__15_ xsel_60_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN1_14 XI11_0/XI0/XI0_60/d__14_ xsel_60_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN1_13 XI11_0/XI0/XI0_60/d__13_ xsel_60_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN1_12 XI11_0/XI0/XI0_60/d__12_ xsel_60_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN1_11 XI11_0/XI0/XI0_60/d__11_ xsel_60_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN1_10 XI11_0/XI0/XI0_60/d__10_ xsel_60_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN1_9 XI11_0/XI0/XI0_60/d__9_ xsel_60_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN1_8 XI11_0/XI0/XI0_60/d__8_ xsel_60_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN1_7 XI11_0/XI0/XI0_60/d__7_ xsel_60_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN1_6 XI11_0/XI0/XI0_60/d__6_ xsel_60_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN1_5 XI11_0/XI0/XI0_60/d__5_ xsel_60_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN1_4 XI11_0/XI0/XI0_60/d__4_ xsel_60_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN1_3 XI11_0/XI0/XI0_60/d__3_ xsel_60_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN1_2 XI11_0/XI0/XI0_60/d__2_ xsel_60_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN1_1 XI11_0/XI0/XI0_60/d__1_ xsel_60_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_60/MN1_0 XI11_0/XI0/XI0_60/d__0_ xsel_60_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN0_15 XI11_0/net21_0_ xsel_59_ XI11_0/XI0/XI0_59/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN0_14 XI11_0/net21_1_ xsel_59_ XI11_0/XI0/XI0_59/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN0_13 XI11_0/net21_2_ xsel_59_ XI11_0/XI0/XI0_59/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN0_12 XI11_0/net21_3_ xsel_59_ XI11_0/XI0/XI0_59/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN0_11 XI11_0/net21_4_ xsel_59_ XI11_0/XI0/XI0_59/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN0_10 XI11_0/net21_5_ xsel_59_ XI11_0/XI0/XI0_59/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN0_9 XI11_0/net21_6_ xsel_59_ XI11_0/XI0/XI0_59/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN0_8 XI11_0/net21_7_ xsel_59_ XI11_0/XI0/XI0_59/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN0_7 XI11_0/net21_8_ xsel_59_ XI11_0/XI0/XI0_59/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN0_6 XI11_0/net21_9_ xsel_59_ XI11_0/XI0/XI0_59/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN0_5 XI11_0/net21_10_ xsel_59_ XI11_0/XI0/XI0_59/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN0_4 XI11_0/net21_11_ xsel_59_ XI11_0/XI0/XI0_59/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN0_3 XI11_0/net21_12_ xsel_59_ XI11_0/XI0/XI0_59/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN0_2 XI11_0/net21_13_ xsel_59_ XI11_0/XI0/XI0_59/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN0_1 XI11_0/net21_14_ xsel_59_ XI11_0/XI0/XI0_59/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN0_0 XI11_0/net21_15_ xsel_59_ XI11_0/XI0/XI0_59/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN1_15 XI11_0/XI0/XI0_59/d__15_ xsel_59_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN1_14 XI11_0/XI0/XI0_59/d__14_ xsel_59_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN1_13 XI11_0/XI0/XI0_59/d__13_ xsel_59_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN1_12 XI11_0/XI0/XI0_59/d__12_ xsel_59_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN1_11 XI11_0/XI0/XI0_59/d__11_ xsel_59_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN1_10 XI11_0/XI0/XI0_59/d__10_ xsel_59_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN1_9 XI11_0/XI0/XI0_59/d__9_ xsel_59_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN1_8 XI11_0/XI0/XI0_59/d__8_ xsel_59_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN1_7 XI11_0/XI0/XI0_59/d__7_ xsel_59_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN1_6 XI11_0/XI0/XI0_59/d__6_ xsel_59_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN1_5 XI11_0/XI0/XI0_59/d__5_ xsel_59_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN1_4 XI11_0/XI0/XI0_59/d__4_ xsel_59_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN1_3 XI11_0/XI0/XI0_59/d__3_ xsel_59_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN1_2 XI11_0/XI0/XI0_59/d__2_ xsel_59_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN1_1 XI11_0/XI0/XI0_59/d__1_ xsel_59_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_59/MN1_0 XI11_0/XI0/XI0_59/d__0_ xsel_59_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN0_15 XI11_0/net21_0_ xsel_58_ XI11_0/XI0/XI0_58/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN0_14 XI11_0/net21_1_ xsel_58_ XI11_0/XI0/XI0_58/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN0_13 XI11_0/net21_2_ xsel_58_ XI11_0/XI0/XI0_58/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN0_12 XI11_0/net21_3_ xsel_58_ XI11_0/XI0/XI0_58/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN0_11 XI11_0/net21_4_ xsel_58_ XI11_0/XI0/XI0_58/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN0_10 XI11_0/net21_5_ xsel_58_ XI11_0/XI0/XI0_58/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN0_9 XI11_0/net21_6_ xsel_58_ XI11_0/XI0/XI0_58/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN0_8 XI11_0/net21_7_ xsel_58_ XI11_0/XI0/XI0_58/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN0_7 XI11_0/net21_8_ xsel_58_ XI11_0/XI0/XI0_58/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN0_6 XI11_0/net21_9_ xsel_58_ XI11_0/XI0/XI0_58/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN0_5 XI11_0/net21_10_ xsel_58_ XI11_0/XI0/XI0_58/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN0_4 XI11_0/net21_11_ xsel_58_ XI11_0/XI0/XI0_58/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN0_3 XI11_0/net21_12_ xsel_58_ XI11_0/XI0/XI0_58/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN0_2 XI11_0/net21_13_ xsel_58_ XI11_0/XI0/XI0_58/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN0_1 XI11_0/net21_14_ xsel_58_ XI11_0/XI0/XI0_58/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN0_0 XI11_0/net21_15_ xsel_58_ XI11_0/XI0/XI0_58/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN1_15 XI11_0/XI0/XI0_58/d__15_ xsel_58_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN1_14 XI11_0/XI0/XI0_58/d__14_ xsel_58_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN1_13 XI11_0/XI0/XI0_58/d__13_ xsel_58_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN1_12 XI11_0/XI0/XI0_58/d__12_ xsel_58_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN1_11 XI11_0/XI0/XI0_58/d__11_ xsel_58_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN1_10 XI11_0/XI0/XI0_58/d__10_ xsel_58_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN1_9 XI11_0/XI0/XI0_58/d__9_ xsel_58_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN1_8 XI11_0/XI0/XI0_58/d__8_ xsel_58_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN1_7 XI11_0/XI0/XI0_58/d__7_ xsel_58_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN1_6 XI11_0/XI0/XI0_58/d__6_ xsel_58_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN1_5 XI11_0/XI0/XI0_58/d__5_ xsel_58_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN1_4 XI11_0/XI0/XI0_58/d__4_ xsel_58_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN1_3 XI11_0/XI0/XI0_58/d__3_ xsel_58_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN1_2 XI11_0/XI0/XI0_58/d__2_ xsel_58_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN1_1 XI11_0/XI0/XI0_58/d__1_ xsel_58_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_58/MN1_0 XI11_0/XI0/XI0_58/d__0_ xsel_58_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN0_15 XI11_0/net21_0_ xsel_57_ XI11_0/XI0/XI0_57/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN0_14 XI11_0/net21_1_ xsel_57_ XI11_0/XI0/XI0_57/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN0_13 XI11_0/net21_2_ xsel_57_ XI11_0/XI0/XI0_57/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN0_12 XI11_0/net21_3_ xsel_57_ XI11_0/XI0/XI0_57/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN0_11 XI11_0/net21_4_ xsel_57_ XI11_0/XI0/XI0_57/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN0_10 XI11_0/net21_5_ xsel_57_ XI11_0/XI0/XI0_57/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN0_9 XI11_0/net21_6_ xsel_57_ XI11_0/XI0/XI0_57/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN0_8 XI11_0/net21_7_ xsel_57_ XI11_0/XI0/XI0_57/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN0_7 XI11_0/net21_8_ xsel_57_ XI11_0/XI0/XI0_57/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN0_6 XI11_0/net21_9_ xsel_57_ XI11_0/XI0/XI0_57/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN0_5 XI11_0/net21_10_ xsel_57_ XI11_0/XI0/XI0_57/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN0_4 XI11_0/net21_11_ xsel_57_ XI11_0/XI0/XI0_57/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN0_3 XI11_0/net21_12_ xsel_57_ XI11_0/XI0/XI0_57/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN0_2 XI11_0/net21_13_ xsel_57_ XI11_0/XI0/XI0_57/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN0_1 XI11_0/net21_14_ xsel_57_ XI11_0/XI0/XI0_57/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN0_0 XI11_0/net21_15_ xsel_57_ XI11_0/XI0/XI0_57/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN1_15 XI11_0/XI0/XI0_57/d__15_ xsel_57_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN1_14 XI11_0/XI0/XI0_57/d__14_ xsel_57_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN1_13 XI11_0/XI0/XI0_57/d__13_ xsel_57_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN1_12 XI11_0/XI0/XI0_57/d__12_ xsel_57_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN1_11 XI11_0/XI0/XI0_57/d__11_ xsel_57_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN1_10 XI11_0/XI0/XI0_57/d__10_ xsel_57_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN1_9 XI11_0/XI0/XI0_57/d__9_ xsel_57_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN1_8 XI11_0/XI0/XI0_57/d__8_ xsel_57_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN1_7 XI11_0/XI0/XI0_57/d__7_ xsel_57_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN1_6 XI11_0/XI0/XI0_57/d__6_ xsel_57_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN1_5 XI11_0/XI0/XI0_57/d__5_ xsel_57_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN1_4 XI11_0/XI0/XI0_57/d__4_ xsel_57_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN1_3 XI11_0/XI0/XI0_57/d__3_ xsel_57_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN1_2 XI11_0/XI0/XI0_57/d__2_ xsel_57_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN1_1 XI11_0/XI0/XI0_57/d__1_ xsel_57_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_57/MN1_0 XI11_0/XI0/XI0_57/d__0_ xsel_57_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN0_15 XI11_0/net21_0_ xsel_56_ XI11_0/XI0/XI0_56/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN0_14 XI11_0/net21_1_ xsel_56_ XI11_0/XI0/XI0_56/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN0_13 XI11_0/net21_2_ xsel_56_ XI11_0/XI0/XI0_56/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN0_12 XI11_0/net21_3_ xsel_56_ XI11_0/XI0/XI0_56/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN0_11 XI11_0/net21_4_ xsel_56_ XI11_0/XI0/XI0_56/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN0_10 XI11_0/net21_5_ xsel_56_ XI11_0/XI0/XI0_56/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN0_9 XI11_0/net21_6_ xsel_56_ XI11_0/XI0/XI0_56/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN0_8 XI11_0/net21_7_ xsel_56_ XI11_0/XI0/XI0_56/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN0_7 XI11_0/net21_8_ xsel_56_ XI11_0/XI0/XI0_56/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN0_6 XI11_0/net21_9_ xsel_56_ XI11_0/XI0/XI0_56/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN0_5 XI11_0/net21_10_ xsel_56_ XI11_0/XI0/XI0_56/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN0_4 XI11_0/net21_11_ xsel_56_ XI11_0/XI0/XI0_56/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN0_3 XI11_0/net21_12_ xsel_56_ XI11_0/XI0/XI0_56/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN0_2 XI11_0/net21_13_ xsel_56_ XI11_0/XI0/XI0_56/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN0_1 XI11_0/net21_14_ xsel_56_ XI11_0/XI0/XI0_56/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN0_0 XI11_0/net21_15_ xsel_56_ XI11_0/XI0/XI0_56/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN1_15 XI11_0/XI0/XI0_56/d__15_ xsel_56_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN1_14 XI11_0/XI0/XI0_56/d__14_ xsel_56_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN1_13 XI11_0/XI0/XI0_56/d__13_ xsel_56_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN1_12 XI11_0/XI0/XI0_56/d__12_ xsel_56_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN1_11 XI11_0/XI0/XI0_56/d__11_ xsel_56_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN1_10 XI11_0/XI0/XI0_56/d__10_ xsel_56_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN1_9 XI11_0/XI0/XI0_56/d__9_ xsel_56_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN1_8 XI11_0/XI0/XI0_56/d__8_ xsel_56_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN1_7 XI11_0/XI0/XI0_56/d__7_ xsel_56_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN1_6 XI11_0/XI0/XI0_56/d__6_ xsel_56_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN1_5 XI11_0/XI0/XI0_56/d__5_ xsel_56_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN1_4 XI11_0/XI0/XI0_56/d__4_ xsel_56_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN1_3 XI11_0/XI0/XI0_56/d__3_ xsel_56_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN1_2 XI11_0/XI0/XI0_56/d__2_ xsel_56_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN1_1 XI11_0/XI0/XI0_56/d__1_ xsel_56_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_56/MN1_0 XI11_0/XI0/XI0_56/d__0_ xsel_56_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN0_15 XI11_0/net21_0_ xsel_55_ XI11_0/XI0/XI0_55/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN0_14 XI11_0/net21_1_ xsel_55_ XI11_0/XI0/XI0_55/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN0_13 XI11_0/net21_2_ xsel_55_ XI11_0/XI0/XI0_55/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN0_12 XI11_0/net21_3_ xsel_55_ XI11_0/XI0/XI0_55/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN0_11 XI11_0/net21_4_ xsel_55_ XI11_0/XI0/XI0_55/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN0_10 XI11_0/net21_5_ xsel_55_ XI11_0/XI0/XI0_55/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN0_9 XI11_0/net21_6_ xsel_55_ XI11_0/XI0/XI0_55/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN0_8 XI11_0/net21_7_ xsel_55_ XI11_0/XI0/XI0_55/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN0_7 XI11_0/net21_8_ xsel_55_ XI11_0/XI0/XI0_55/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN0_6 XI11_0/net21_9_ xsel_55_ XI11_0/XI0/XI0_55/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN0_5 XI11_0/net21_10_ xsel_55_ XI11_0/XI0/XI0_55/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN0_4 XI11_0/net21_11_ xsel_55_ XI11_0/XI0/XI0_55/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN0_3 XI11_0/net21_12_ xsel_55_ XI11_0/XI0/XI0_55/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN0_2 XI11_0/net21_13_ xsel_55_ XI11_0/XI0/XI0_55/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN0_1 XI11_0/net21_14_ xsel_55_ XI11_0/XI0/XI0_55/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN0_0 XI11_0/net21_15_ xsel_55_ XI11_0/XI0/XI0_55/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN1_15 XI11_0/XI0/XI0_55/d__15_ xsel_55_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN1_14 XI11_0/XI0/XI0_55/d__14_ xsel_55_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN1_13 XI11_0/XI0/XI0_55/d__13_ xsel_55_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN1_12 XI11_0/XI0/XI0_55/d__12_ xsel_55_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN1_11 XI11_0/XI0/XI0_55/d__11_ xsel_55_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN1_10 XI11_0/XI0/XI0_55/d__10_ xsel_55_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN1_9 XI11_0/XI0/XI0_55/d__9_ xsel_55_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN1_8 XI11_0/XI0/XI0_55/d__8_ xsel_55_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN1_7 XI11_0/XI0/XI0_55/d__7_ xsel_55_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN1_6 XI11_0/XI0/XI0_55/d__6_ xsel_55_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN1_5 XI11_0/XI0/XI0_55/d__5_ xsel_55_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN1_4 XI11_0/XI0/XI0_55/d__4_ xsel_55_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN1_3 XI11_0/XI0/XI0_55/d__3_ xsel_55_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN1_2 XI11_0/XI0/XI0_55/d__2_ xsel_55_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN1_1 XI11_0/XI0/XI0_55/d__1_ xsel_55_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_55/MN1_0 XI11_0/XI0/XI0_55/d__0_ xsel_55_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN0_15 XI11_0/net21_0_ xsel_54_ XI11_0/XI0/XI0_54/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN0_14 XI11_0/net21_1_ xsel_54_ XI11_0/XI0/XI0_54/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN0_13 XI11_0/net21_2_ xsel_54_ XI11_0/XI0/XI0_54/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN0_12 XI11_0/net21_3_ xsel_54_ XI11_0/XI0/XI0_54/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN0_11 XI11_0/net21_4_ xsel_54_ XI11_0/XI0/XI0_54/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN0_10 XI11_0/net21_5_ xsel_54_ XI11_0/XI0/XI0_54/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN0_9 XI11_0/net21_6_ xsel_54_ XI11_0/XI0/XI0_54/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN0_8 XI11_0/net21_7_ xsel_54_ XI11_0/XI0/XI0_54/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN0_7 XI11_0/net21_8_ xsel_54_ XI11_0/XI0/XI0_54/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN0_6 XI11_0/net21_9_ xsel_54_ XI11_0/XI0/XI0_54/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN0_5 XI11_0/net21_10_ xsel_54_ XI11_0/XI0/XI0_54/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN0_4 XI11_0/net21_11_ xsel_54_ XI11_0/XI0/XI0_54/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN0_3 XI11_0/net21_12_ xsel_54_ XI11_0/XI0/XI0_54/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN0_2 XI11_0/net21_13_ xsel_54_ XI11_0/XI0/XI0_54/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN0_1 XI11_0/net21_14_ xsel_54_ XI11_0/XI0/XI0_54/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN0_0 XI11_0/net21_15_ xsel_54_ XI11_0/XI0/XI0_54/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN1_15 XI11_0/XI0/XI0_54/d__15_ xsel_54_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN1_14 XI11_0/XI0/XI0_54/d__14_ xsel_54_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN1_13 XI11_0/XI0/XI0_54/d__13_ xsel_54_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN1_12 XI11_0/XI0/XI0_54/d__12_ xsel_54_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN1_11 XI11_0/XI0/XI0_54/d__11_ xsel_54_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN1_10 XI11_0/XI0/XI0_54/d__10_ xsel_54_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN1_9 XI11_0/XI0/XI0_54/d__9_ xsel_54_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN1_8 XI11_0/XI0/XI0_54/d__8_ xsel_54_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN1_7 XI11_0/XI0/XI0_54/d__7_ xsel_54_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN1_6 XI11_0/XI0/XI0_54/d__6_ xsel_54_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN1_5 XI11_0/XI0/XI0_54/d__5_ xsel_54_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN1_4 XI11_0/XI0/XI0_54/d__4_ xsel_54_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN1_3 XI11_0/XI0/XI0_54/d__3_ xsel_54_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN1_2 XI11_0/XI0/XI0_54/d__2_ xsel_54_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN1_1 XI11_0/XI0/XI0_54/d__1_ xsel_54_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_54/MN1_0 XI11_0/XI0/XI0_54/d__0_ xsel_54_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN0_15 XI11_0/net21_0_ xsel_53_ XI11_0/XI0/XI0_53/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN0_14 XI11_0/net21_1_ xsel_53_ XI11_0/XI0/XI0_53/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN0_13 XI11_0/net21_2_ xsel_53_ XI11_0/XI0/XI0_53/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN0_12 XI11_0/net21_3_ xsel_53_ XI11_0/XI0/XI0_53/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN0_11 XI11_0/net21_4_ xsel_53_ XI11_0/XI0/XI0_53/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN0_10 XI11_0/net21_5_ xsel_53_ XI11_0/XI0/XI0_53/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN0_9 XI11_0/net21_6_ xsel_53_ XI11_0/XI0/XI0_53/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN0_8 XI11_0/net21_7_ xsel_53_ XI11_0/XI0/XI0_53/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN0_7 XI11_0/net21_8_ xsel_53_ XI11_0/XI0/XI0_53/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN0_6 XI11_0/net21_9_ xsel_53_ XI11_0/XI0/XI0_53/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN0_5 XI11_0/net21_10_ xsel_53_ XI11_0/XI0/XI0_53/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN0_4 XI11_0/net21_11_ xsel_53_ XI11_0/XI0/XI0_53/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN0_3 XI11_0/net21_12_ xsel_53_ XI11_0/XI0/XI0_53/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN0_2 XI11_0/net21_13_ xsel_53_ XI11_0/XI0/XI0_53/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN0_1 XI11_0/net21_14_ xsel_53_ XI11_0/XI0/XI0_53/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN0_0 XI11_0/net21_15_ xsel_53_ XI11_0/XI0/XI0_53/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN1_15 XI11_0/XI0/XI0_53/d__15_ xsel_53_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN1_14 XI11_0/XI0/XI0_53/d__14_ xsel_53_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN1_13 XI11_0/XI0/XI0_53/d__13_ xsel_53_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN1_12 XI11_0/XI0/XI0_53/d__12_ xsel_53_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN1_11 XI11_0/XI0/XI0_53/d__11_ xsel_53_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN1_10 XI11_0/XI0/XI0_53/d__10_ xsel_53_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN1_9 XI11_0/XI0/XI0_53/d__9_ xsel_53_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN1_8 XI11_0/XI0/XI0_53/d__8_ xsel_53_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN1_7 XI11_0/XI0/XI0_53/d__7_ xsel_53_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN1_6 XI11_0/XI0/XI0_53/d__6_ xsel_53_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN1_5 XI11_0/XI0/XI0_53/d__5_ xsel_53_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN1_4 XI11_0/XI0/XI0_53/d__4_ xsel_53_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN1_3 XI11_0/XI0/XI0_53/d__3_ xsel_53_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN1_2 XI11_0/XI0/XI0_53/d__2_ xsel_53_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN1_1 XI11_0/XI0/XI0_53/d__1_ xsel_53_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_53/MN1_0 XI11_0/XI0/XI0_53/d__0_ xsel_53_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN0_15 XI11_0/net21_0_ xsel_52_ XI11_0/XI0/XI0_52/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN0_14 XI11_0/net21_1_ xsel_52_ XI11_0/XI0/XI0_52/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN0_13 XI11_0/net21_2_ xsel_52_ XI11_0/XI0/XI0_52/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN0_12 XI11_0/net21_3_ xsel_52_ XI11_0/XI0/XI0_52/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN0_11 XI11_0/net21_4_ xsel_52_ XI11_0/XI0/XI0_52/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN0_10 XI11_0/net21_5_ xsel_52_ XI11_0/XI0/XI0_52/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN0_9 XI11_0/net21_6_ xsel_52_ XI11_0/XI0/XI0_52/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN0_8 XI11_0/net21_7_ xsel_52_ XI11_0/XI0/XI0_52/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN0_7 XI11_0/net21_8_ xsel_52_ XI11_0/XI0/XI0_52/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN0_6 XI11_0/net21_9_ xsel_52_ XI11_0/XI0/XI0_52/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN0_5 XI11_0/net21_10_ xsel_52_ XI11_0/XI0/XI0_52/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN0_4 XI11_0/net21_11_ xsel_52_ XI11_0/XI0/XI0_52/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN0_3 XI11_0/net21_12_ xsel_52_ XI11_0/XI0/XI0_52/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN0_2 XI11_0/net21_13_ xsel_52_ XI11_0/XI0/XI0_52/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN0_1 XI11_0/net21_14_ xsel_52_ XI11_0/XI0/XI0_52/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN0_0 XI11_0/net21_15_ xsel_52_ XI11_0/XI0/XI0_52/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN1_15 XI11_0/XI0/XI0_52/d__15_ xsel_52_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN1_14 XI11_0/XI0/XI0_52/d__14_ xsel_52_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN1_13 XI11_0/XI0/XI0_52/d__13_ xsel_52_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN1_12 XI11_0/XI0/XI0_52/d__12_ xsel_52_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN1_11 XI11_0/XI0/XI0_52/d__11_ xsel_52_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN1_10 XI11_0/XI0/XI0_52/d__10_ xsel_52_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN1_9 XI11_0/XI0/XI0_52/d__9_ xsel_52_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN1_8 XI11_0/XI0/XI0_52/d__8_ xsel_52_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN1_7 XI11_0/XI0/XI0_52/d__7_ xsel_52_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN1_6 XI11_0/XI0/XI0_52/d__6_ xsel_52_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN1_5 XI11_0/XI0/XI0_52/d__5_ xsel_52_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN1_4 XI11_0/XI0/XI0_52/d__4_ xsel_52_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN1_3 XI11_0/XI0/XI0_52/d__3_ xsel_52_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN1_2 XI11_0/XI0/XI0_52/d__2_ xsel_52_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN1_1 XI11_0/XI0/XI0_52/d__1_ xsel_52_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_52/MN1_0 XI11_0/XI0/XI0_52/d__0_ xsel_52_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN0_15 XI11_0/net21_0_ xsel_51_ XI11_0/XI0/XI0_51/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN0_14 XI11_0/net21_1_ xsel_51_ XI11_0/XI0/XI0_51/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN0_13 XI11_0/net21_2_ xsel_51_ XI11_0/XI0/XI0_51/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN0_12 XI11_0/net21_3_ xsel_51_ XI11_0/XI0/XI0_51/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN0_11 XI11_0/net21_4_ xsel_51_ XI11_0/XI0/XI0_51/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN0_10 XI11_0/net21_5_ xsel_51_ XI11_0/XI0/XI0_51/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN0_9 XI11_0/net21_6_ xsel_51_ XI11_0/XI0/XI0_51/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN0_8 XI11_0/net21_7_ xsel_51_ XI11_0/XI0/XI0_51/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN0_7 XI11_0/net21_8_ xsel_51_ XI11_0/XI0/XI0_51/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN0_6 XI11_0/net21_9_ xsel_51_ XI11_0/XI0/XI0_51/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN0_5 XI11_0/net21_10_ xsel_51_ XI11_0/XI0/XI0_51/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN0_4 XI11_0/net21_11_ xsel_51_ XI11_0/XI0/XI0_51/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN0_3 XI11_0/net21_12_ xsel_51_ XI11_0/XI0/XI0_51/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN0_2 XI11_0/net21_13_ xsel_51_ XI11_0/XI0/XI0_51/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN0_1 XI11_0/net21_14_ xsel_51_ XI11_0/XI0/XI0_51/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN0_0 XI11_0/net21_15_ xsel_51_ XI11_0/XI0/XI0_51/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN1_15 XI11_0/XI0/XI0_51/d__15_ xsel_51_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN1_14 XI11_0/XI0/XI0_51/d__14_ xsel_51_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN1_13 XI11_0/XI0/XI0_51/d__13_ xsel_51_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN1_12 XI11_0/XI0/XI0_51/d__12_ xsel_51_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN1_11 XI11_0/XI0/XI0_51/d__11_ xsel_51_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN1_10 XI11_0/XI0/XI0_51/d__10_ xsel_51_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN1_9 XI11_0/XI0/XI0_51/d__9_ xsel_51_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN1_8 XI11_0/XI0/XI0_51/d__8_ xsel_51_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN1_7 XI11_0/XI0/XI0_51/d__7_ xsel_51_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN1_6 XI11_0/XI0/XI0_51/d__6_ xsel_51_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN1_5 XI11_0/XI0/XI0_51/d__5_ xsel_51_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN1_4 XI11_0/XI0/XI0_51/d__4_ xsel_51_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN1_3 XI11_0/XI0/XI0_51/d__3_ xsel_51_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN1_2 XI11_0/XI0/XI0_51/d__2_ xsel_51_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN1_1 XI11_0/XI0/XI0_51/d__1_ xsel_51_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_51/MN1_0 XI11_0/XI0/XI0_51/d__0_ xsel_51_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN0_15 XI11_0/net21_0_ xsel_50_ XI11_0/XI0/XI0_50/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN0_14 XI11_0/net21_1_ xsel_50_ XI11_0/XI0/XI0_50/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN0_13 XI11_0/net21_2_ xsel_50_ XI11_0/XI0/XI0_50/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN0_12 XI11_0/net21_3_ xsel_50_ XI11_0/XI0/XI0_50/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN0_11 XI11_0/net21_4_ xsel_50_ XI11_0/XI0/XI0_50/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN0_10 XI11_0/net21_5_ xsel_50_ XI11_0/XI0/XI0_50/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN0_9 XI11_0/net21_6_ xsel_50_ XI11_0/XI0/XI0_50/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN0_8 XI11_0/net21_7_ xsel_50_ XI11_0/XI0/XI0_50/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN0_7 XI11_0/net21_8_ xsel_50_ XI11_0/XI0/XI0_50/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN0_6 XI11_0/net21_9_ xsel_50_ XI11_0/XI0/XI0_50/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN0_5 XI11_0/net21_10_ xsel_50_ XI11_0/XI0/XI0_50/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN0_4 XI11_0/net21_11_ xsel_50_ XI11_0/XI0/XI0_50/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN0_3 XI11_0/net21_12_ xsel_50_ XI11_0/XI0/XI0_50/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN0_2 XI11_0/net21_13_ xsel_50_ XI11_0/XI0/XI0_50/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN0_1 XI11_0/net21_14_ xsel_50_ XI11_0/XI0/XI0_50/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN0_0 XI11_0/net21_15_ xsel_50_ XI11_0/XI0/XI0_50/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN1_15 XI11_0/XI0/XI0_50/d__15_ xsel_50_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN1_14 XI11_0/XI0/XI0_50/d__14_ xsel_50_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN1_13 XI11_0/XI0/XI0_50/d__13_ xsel_50_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN1_12 XI11_0/XI0/XI0_50/d__12_ xsel_50_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN1_11 XI11_0/XI0/XI0_50/d__11_ xsel_50_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN1_10 XI11_0/XI0/XI0_50/d__10_ xsel_50_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN1_9 XI11_0/XI0/XI0_50/d__9_ xsel_50_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN1_8 XI11_0/XI0/XI0_50/d__8_ xsel_50_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN1_7 XI11_0/XI0/XI0_50/d__7_ xsel_50_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN1_6 XI11_0/XI0/XI0_50/d__6_ xsel_50_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN1_5 XI11_0/XI0/XI0_50/d__5_ xsel_50_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN1_4 XI11_0/XI0/XI0_50/d__4_ xsel_50_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN1_3 XI11_0/XI0/XI0_50/d__3_ xsel_50_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN1_2 XI11_0/XI0/XI0_50/d__2_ xsel_50_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN1_1 XI11_0/XI0/XI0_50/d__1_ xsel_50_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_50/MN1_0 XI11_0/XI0/XI0_50/d__0_ xsel_50_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN0_15 XI11_0/net21_0_ xsel_49_ XI11_0/XI0/XI0_49/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN0_14 XI11_0/net21_1_ xsel_49_ XI11_0/XI0/XI0_49/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN0_13 XI11_0/net21_2_ xsel_49_ XI11_0/XI0/XI0_49/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN0_12 XI11_0/net21_3_ xsel_49_ XI11_0/XI0/XI0_49/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN0_11 XI11_0/net21_4_ xsel_49_ XI11_0/XI0/XI0_49/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN0_10 XI11_0/net21_5_ xsel_49_ XI11_0/XI0/XI0_49/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN0_9 XI11_0/net21_6_ xsel_49_ XI11_0/XI0/XI0_49/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN0_8 XI11_0/net21_7_ xsel_49_ XI11_0/XI0/XI0_49/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN0_7 XI11_0/net21_8_ xsel_49_ XI11_0/XI0/XI0_49/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN0_6 XI11_0/net21_9_ xsel_49_ XI11_0/XI0/XI0_49/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN0_5 XI11_0/net21_10_ xsel_49_ XI11_0/XI0/XI0_49/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN0_4 XI11_0/net21_11_ xsel_49_ XI11_0/XI0/XI0_49/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN0_3 XI11_0/net21_12_ xsel_49_ XI11_0/XI0/XI0_49/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN0_2 XI11_0/net21_13_ xsel_49_ XI11_0/XI0/XI0_49/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN0_1 XI11_0/net21_14_ xsel_49_ XI11_0/XI0/XI0_49/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN0_0 XI11_0/net21_15_ xsel_49_ XI11_0/XI0/XI0_49/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN1_15 XI11_0/XI0/XI0_49/d__15_ xsel_49_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN1_14 XI11_0/XI0/XI0_49/d__14_ xsel_49_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN1_13 XI11_0/XI0/XI0_49/d__13_ xsel_49_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN1_12 XI11_0/XI0/XI0_49/d__12_ xsel_49_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN1_11 XI11_0/XI0/XI0_49/d__11_ xsel_49_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN1_10 XI11_0/XI0/XI0_49/d__10_ xsel_49_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN1_9 XI11_0/XI0/XI0_49/d__9_ xsel_49_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN1_8 XI11_0/XI0/XI0_49/d__8_ xsel_49_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN1_7 XI11_0/XI0/XI0_49/d__7_ xsel_49_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN1_6 XI11_0/XI0/XI0_49/d__6_ xsel_49_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN1_5 XI11_0/XI0/XI0_49/d__5_ xsel_49_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN1_4 XI11_0/XI0/XI0_49/d__4_ xsel_49_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN1_3 XI11_0/XI0/XI0_49/d__3_ xsel_49_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN1_2 XI11_0/XI0/XI0_49/d__2_ xsel_49_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN1_1 XI11_0/XI0/XI0_49/d__1_ xsel_49_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_49/MN1_0 XI11_0/XI0/XI0_49/d__0_ xsel_49_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN0_15 XI11_0/net21_0_ xsel_48_ XI11_0/XI0/XI0_48/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN0_14 XI11_0/net21_1_ xsel_48_ XI11_0/XI0/XI0_48/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN0_13 XI11_0/net21_2_ xsel_48_ XI11_0/XI0/XI0_48/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN0_12 XI11_0/net21_3_ xsel_48_ XI11_0/XI0/XI0_48/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN0_11 XI11_0/net21_4_ xsel_48_ XI11_0/XI0/XI0_48/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN0_10 XI11_0/net21_5_ xsel_48_ XI11_0/XI0/XI0_48/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN0_9 XI11_0/net21_6_ xsel_48_ XI11_0/XI0/XI0_48/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN0_8 XI11_0/net21_7_ xsel_48_ XI11_0/XI0/XI0_48/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN0_7 XI11_0/net21_8_ xsel_48_ XI11_0/XI0/XI0_48/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN0_6 XI11_0/net21_9_ xsel_48_ XI11_0/XI0/XI0_48/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN0_5 XI11_0/net21_10_ xsel_48_ XI11_0/XI0/XI0_48/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN0_4 XI11_0/net21_11_ xsel_48_ XI11_0/XI0/XI0_48/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN0_3 XI11_0/net21_12_ xsel_48_ XI11_0/XI0/XI0_48/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN0_2 XI11_0/net21_13_ xsel_48_ XI11_0/XI0/XI0_48/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN0_1 XI11_0/net21_14_ xsel_48_ XI11_0/XI0/XI0_48/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN0_0 XI11_0/net21_15_ xsel_48_ XI11_0/XI0/XI0_48/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN1_15 XI11_0/XI0/XI0_48/d__15_ xsel_48_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN1_14 XI11_0/XI0/XI0_48/d__14_ xsel_48_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN1_13 XI11_0/XI0/XI0_48/d__13_ xsel_48_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN1_12 XI11_0/XI0/XI0_48/d__12_ xsel_48_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN1_11 XI11_0/XI0/XI0_48/d__11_ xsel_48_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN1_10 XI11_0/XI0/XI0_48/d__10_ xsel_48_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN1_9 XI11_0/XI0/XI0_48/d__9_ xsel_48_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN1_8 XI11_0/XI0/XI0_48/d__8_ xsel_48_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN1_7 XI11_0/XI0/XI0_48/d__7_ xsel_48_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN1_6 XI11_0/XI0/XI0_48/d__6_ xsel_48_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN1_5 XI11_0/XI0/XI0_48/d__5_ xsel_48_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN1_4 XI11_0/XI0/XI0_48/d__4_ xsel_48_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN1_3 XI11_0/XI0/XI0_48/d__3_ xsel_48_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN1_2 XI11_0/XI0/XI0_48/d__2_ xsel_48_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN1_1 XI11_0/XI0/XI0_48/d__1_ xsel_48_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_48/MN1_0 XI11_0/XI0/XI0_48/d__0_ xsel_48_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN0_15 XI11_0/net21_0_ xsel_47_ XI11_0/XI0/XI0_47/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN0_14 XI11_0/net21_1_ xsel_47_ XI11_0/XI0/XI0_47/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN0_13 XI11_0/net21_2_ xsel_47_ XI11_0/XI0/XI0_47/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN0_12 XI11_0/net21_3_ xsel_47_ XI11_0/XI0/XI0_47/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN0_11 XI11_0/net21_4_ xsel_47_ XI11_0/XI0/XI0_47/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN0_10 XI11_0/net21_5_ xsel_47_ XI11_0/XI0/XI0_47/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN0_9 XI11_0/net21_6_ xsel_47_ XI11_0/XI0/XI0_47/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN0_8 XI11_0/net21_7_ xsel_47_ XI11_0/XI0/XI0_47/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN0_7 XI11_0/net21_8_ xsel_47_ XI11_0/XI0/XI0_47/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN0_6 XI11_0/net21_9_ xsel_47_ XI11_0/XI0/XI0_47/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN0_5 XI11_0/net21_10_ xsel_47_ XI11_0/XI0/XI0_47/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN0_4 XI11_0/net21_11_ xsel_47_ XI11_0/XI0/XI0_47/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN0_3 XI11_0/net21_12_ xsel_47_ XI11_0/XI0/XI0_47/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN0_2 XI11_0/net21_13_ xsel_47_ XI11_0/XI0/XI0_47/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN0_1 XI11_0/net21_14_ xsel_47_ XI11_0/XI0/XI0_47/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN0_0 XI11_0/net21_15_ xsel_47_ XI11_0/XI0/XI0_47/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN1_15 XI11_0/XI0/XI0_47/d__15_ xsel_47_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN1_14 XI11_0/XI0/XI0_47/d__14_ xsel_47_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN1_13 XI11_0/XI0/XI0_47/d__13_ xsel_47_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN1_12 XI11_0/XI0/XI0_47/d__12_ xsel_47_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN1_11 XI11_0/XI0/XI0_47/d__11_ xsel_47_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN1_10 XI11_0/XI0/XI0_47/d__10_ xsel_47_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN1_9 XI11_0/XI0/XI0_47/d__9_ xsel_47_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN1_8 XI11_0/XI0/XI0_47/d__8_ xsel_47_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN1_7 XI11_0/XI0/XI0_47/d__7_ xsel_47_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN1_6 XI11_0/XI0/XI0_47/d__6_ xsel_47_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN1_5 XI11_0/XI0/XI0_47/d__5_ xsel_47_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN1_4 XI11_0/XI0/XI0_47/d__4_ xsel_47_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN1_3 XI11_0/XI0/XI0_47/d__3_ xsel_47_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN1_2 XI11_0/XI0/XI0_47/d__2_ xsel_47_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN1_1 XI11_0/XI0/XI0_47/d__1_ xsel_47_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_47/MN1_0 XI11_0/XI0/XI0_47/d__0_ xsel_47_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN0_15 XI11_0/net21_0_ xsel_46_ XI11_0/XI0/XI0_46/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN0_14 XI11_0/net21_1_ xsel_46_ XI11_0/XI0/XI0_46/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN0_13 XI11_0/net21_2_ xsel_46_ XI11_0/XI0/XI0_46/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN0_12 XI11_0/net21_3_ xsel_46_ XI11_0/XI0/XI0_46/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN0_11 XI11_0/net21_4_ xsel_46_ XI11_0/XI0/XI0_46/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN0_10 XI11_0/net21_5_ xsel_46_ XI11_0/XI0/XI0_46/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN0_9 XI11_0/net21_6_ xsel_46_ XI11_0/XI0/XI0_46/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN0_8 XI11_0/net21_7_ xsel_46_ XI11_0/XI0/XI0_46/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN0_7 XI11_0/net21_8_ xsel_46_ XI11_0/XI0/XI0_46/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN0_6 XI11_0/net21_9_ xsel_46_ XI11_0/XI0/XI0_46/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN0_5 XI11_0/net21_10_ xsel_46_ XI11_0/XI0/XI0_46/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN0_4 XI11_0/net21_11_ xsel_46_ XI11_0/XI0/XI0_46/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN0_3 XI11_0/net21_12_ xsel_46_ XI11_0/XI0/XI0_46/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN0_2 XI11_0/net21_13_ xsel_46_ XI11_0/XI0/XI0_46/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN0_1 XI11_0/net21_14_ xsel_46_ XI11_0/XI0/XI0_46/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN0_0 XI11_0/net21_15_ xsel_46_ XI11_0/XI0/XI0_46/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN1_15 XI11_0/XI0/XI0_46/d__15_ xsel_46_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN1_14 XI11_0/XI0/XI0_46/d__14_ xsel_46_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN1_13 XI11_0/XI0/XI0_46/d__13_ xsel_46_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN1_12 XI11_0/XI0/XI0_46/d__12_ xsel_46_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN1_11 XI11_0/XI0/XI0_46/d__11_ xsel_46_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN1_10 XI11_0/XI0/XI0_46/d__10_ xsel_46_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN1_9 XI11_0/XI0/XI0_46/d__9_ xsel_46_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN1_8 XI11_0/XI0/XI0_46/d__8_ xsel_46_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN1_7 XI11_0/XI0/XI0_46/d__7_ xsel_46_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN1_6 XI11_0/XI0/XI0_46/d__6_ xsel_46_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN1_5 XI11_0/XI0/XI0_46/d__5_ xsel_46_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN1_4 XI11_0/XI0/XI0_46/d__4_ xsel_46_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN1_3 XI11_0/XI0/XI0_46/d__3_ xsel_46_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN1_2 XI11_0/XI0/XI0_46/d__2_ xsel_46_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN1_1 XI11_0/XI0/XI0_46/d__1_ xsel_46_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_46/MN1_0 XI11_0/XI0/XI0_46/d__0_ xsel_46_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN0_15 XI11_0/net21_0_ xsel_45_ XI11_0/XI0/XI0_45/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN0_14 XI11_0/net21_1_ xsel_45_ XI11_0/XI0/XI0_45/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN0_13 XI11_0/net21_2_ xsel_45_ XI11_0/XI0/XI0_45/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN0_12 XI11_0/net21_3_ xsel_45_ XI11_0/XI0/XI0_45/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN0_11 XI11_0/net21_4_ xsel_45_ XI11_0/XI0/XI0_45/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN0_10 XI11_0/net21_5_ xsel_45_ XI11_0/XI0/XI0_45/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN0_9 XI11_0/net21_6_ xsel_45_ XI11_0/XI0/XI0_45/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN0_8 XI11_0/net21_7_ xsel_45_ XI11_0/XI0/XI0_45/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN0_7 XI11_0/net21_8_ xsel_45_ XI11_0/XI0/XI0_45/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN0_6 XI11_0/net21_9_ xsel_45_ XI11_0/XI0/XI0_45/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN0_5 XI11_0/net21_10_ xsel_45_ XI11_0/XI0/XI0_45/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN0_4 XI11_0/net21_11_ xsel_45_ XI11_0/XI0/XI0_45/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN0_3 XI11_0/net21_12_ xsel_45_ XI11_0/XI0/XI0_45/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN0_2 XI11_0/net21_13_ xsel_45_ XI11_0/XI0/XI0_45/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN0_1 XI11_0/net21_14_ xsel_45_ XI11_0/XI0/XI0_45/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN0_0 XI11_0/net21_15_ xsel_45_ XI11_0/XI0/XI0_45/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN1_15 XI11_0/XI0/XI0_45/d__15_ xsel_45_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN1_14 XI11_0/XI0/XI0_45/d__14_ xsel_45_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN1_13 XI11_0/XI0/XI0_45/d__13_ xsel_45_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN1_12 XI11_0/XI0/XI0_45/d__12_ xsel_45_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN1_11 XI11_0/XI0/XI0_45/d__11_ xsel_45_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN1_10 XI11_0/XI0/XI0_45/d__10_ xsel_45_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN1_9 XI11_0/XI0/XI0_45/d__9_ xsel_45_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN1_8 XI11_0/XI0/XI0_45/d__8_ xsel_45_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN1_7 XI11_0/XI0/XI0_45/d__7_ xsel_45_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN1_6 XI11_0/XI0/XI0_45/d__6_ xsel_45_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN1_5 XI11_0/XI0/XI0_45/d__5_ xsel_45_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN1_4 XI11_0/XI0/XI0_45/d__4_ xsel_45_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN1_3 XI11_0/XI0/XI0_45/d__3_ xsel_45_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN1_2 XI11_0/XI0/XI0_45/d__2_ xsel_45_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN1_1 XI11_0/XI0/XI0_45/d__1_ xsel_45_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_45/MN1_0 XI11_0/XI0/XI0_45/d__0_ xsel_45_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN0_15 XI11_0/net21_0_ xsel_44_ XI11_0/XI0/XI0_44/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN0_14 XI11_0/net21_1_ xsel_44_ XI11_0/XI0/XI0_44/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN0_13 XI11_0/net21_2_ xsel_44_ XI11_0/XI0/XI0_44/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN0_12 XI11_0/net21_3_ xsel_44_ XI11_0/XI0/XI0_44/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN0_11 XI11_0/net21_4_ xsel_44_ XI11_0/XI0/XI0_44/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN0_10 XI11_0/net21_5_ xsel_44_ XI11_0/XI0/XI0_44/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN0_9 XI11_0/net21_6_ xsel_44_ XI11_0/XI0/XI0_44/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN0_8 XI11_0/net21_7_ xsel_44_ XI11_0/XI0/XI0_44/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN0_7 XI11_0/net21_8_ xsel_44_ XI11_0/XI0/XI0_44/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN0_6 XI11_0/net21_9_ xsel_44_ XI11_0/XI0/XI0_44/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN0_5 XI11_0/net21_10_ xsel_44_ XI11_0/XI0/XI0_44/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN0_4 XI11_0/net21_11_ xsel_44_ XI11_0/XI0/XI0_44/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN0_3 XI11_0/net21_12_ xsel_44_ XI11_0/XI0/XI0_44/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN0_2 XI11_0/net21_13_ xsel_44_ XI11_0/XI0/XI0_44/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN0_1 XI11_0/net21_14_ xsel_44_ XI11_0/XI0/XI0_44/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN0_0 XI11_0/net21_15_ xsel_44_ XI11_0/XI0/XI0_44/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN1_15 XI11_0/XI0/XI0_44/d__15_ xsel_44_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN1_14 XI11_0/XI0/XI0_44/d__14_ xsel_44_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN1_13 XI11_0/XI0/XI0_44/d__13_ xsel_44_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN1_12 XI11_0/XI0/XI0_44/d__12_ xsel_44_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN1_11 XI11_0/XI0/XI0_44/d__11_ xsel_44_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN1_10 XI11_0/XI0/XI0_44/d__10_ xsel_44_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN1_9 XI11_0/XI0/XI0_44/d__9_ xsel_44_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN1_8 XI11_0/XI0/XI0_44/d__8_ xsel_44_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN1_7 XI11_0/XI0/XI0_44/d__7_ xsel_44_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN1_6 XI11_0/XI0/XI0_44/d__6_ xsel_44_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN1_5 XI11_0/XI0/XI0_44/d__5_ xsel_44_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN1_4 XI11_0/XI0/XI0_44/d__4_ xsel_44_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN1_3 XI11_0/XI0/XI0_44/d__3_ xsel_44_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN1_2 XI11_0/XI0/XI0_44/d__2_ xsel_44_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN1_1 XI11_0/XI0/XI0_44/d__1_ xsel_44_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_44/MN1_0 XI11_0/XI0/XI0_44/d__0_ xsel_44_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN0_15 XI11_0/net21_0_ xsel_43_ XI11_0/XI0/XI0_43/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN0_14 XI11_0/net21_1_ xsel_43_ XI11_0/XI0/XI0_43/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN0_13 XI11_0/net21_2_ xsel_43_ XI11_0/XI0/XI0_43/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN0_12 XI11_0/net21_3_ xsel_43_ XI11_0/XI0/XI0_43/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN0_11 XI11_0/net21_4_ xsel_43_ XI11_0/XI0/XI0_43/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN0_10 XI11_0/net21_5_ xsel_43_ XI11_0/XI0/XI0_43/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN0_9 XI11_0/net21_6_ xsel_43_ XI11_0/XI0/XI0_43/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN0_8 XI11_0/net21_7_ xsel_43_ XI11_0/XI0/XI0_43/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN0_7 XI11_0/net21_8_ xsel_43_ XI11_0/XI0/XI0_43/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN0_6 XI11_0/net21_9_ xsel_43_ XI11_0/XI0/XI0_43/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN0_5 XI11_0/net21_10_ xsel_43_ XI11_0/XI0/XI0_43/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN0_4 XI11_0/net21_11_ xsel_43_ XI11_0/XI0/XI0_43/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN0_3 XI11_0/net21_12_ xsel_43_ XI11_0/XI0/XI0_43/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN0_2 XI11_0/net21_13_ xsel_43_ XI11_0/XI0/XI0_43/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN0_1 XI11_0/net21_14_ xsel_43_ XI11_0/XI0/XI0_43/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN0_0 XI11_0/net21_15_ xsel_43_ XI11_0/XI0/XI0_43/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN1_15 XI11_0/XI0/XI0_43/d__15_ xsel_43_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN1_14 XI11_0/XI0/XI0_43/d__14_ xsel_43_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN1_13 XI11_0/XI0/XI0_43/d__13_ xsel_43_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN1_12 XI11_0/XI0/XI0_43/d__12_ xsel_43_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN1_11 XI11_0/XI0/XI0_43/d__11_ xsel_43_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN1_10 XI11_0/XI0/XI0_43/d__10_ xsel_43_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN1_9 XI11_0/XI0/XI0_43/d__9_ xsel_43_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN1_8 XI11_0/XI0/XI0_43/d__8_ xsel_43_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN1_7 XI11_0/XI0/XI0_43/d__7_ xsel_43_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN1_6 XI11_0/XI0/XI0_43/d__6_ xsel_43_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN1_5 XI11_0/XI0/XI0_43/d__5_ xsel_43_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN1_4 XI11_0/XI0/XI0_43/d__4_ xsel_43_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN1_3 XI11_0/XI0/XI0_43/d__3_ xsel_43_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN1_2 XI11_0/XI0/XI0_43/d__2_ xsel_43_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN1_1 XI11_0/XI0/XI0_43/d__1_ xsel_43_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_43/MN1_0 XI11_0/XI0/XI0_43/d__0_ xsel_43_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN0_15 XI11_0/net21_0_ xsel_42_ XI11_0/XI0/XI0_42/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN0_14 XI11_0/net21_1_ xsel_42_ XI11_0/XI0/XI0_42/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN0_13 XI11_0/net21_2_ xsel_42_ XI11_0/XI0/XI0_42/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN0_12 XI11_0/net21_3_ xsel_42_ XI11_0/XI0/XI0_42/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN0_11 XI11_0/net21_4_ xsel_42_ XI11_0/XI0/XI0_42/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN0_10 XI11_0/net21_5_ xsel_42_ XI11_0/XI0/XI0_42/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN0_9 XI11_0/net21_6_ xsel_42_ XI11_0/XI0/XI0_42/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN0_8 XI11_0/net21_7_ xsel_42_ XI11_0/XI0/XI0_42/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN0_7 XI11_0/net21_8_ xsel_42_ XI11_0/XI0/XI0_42/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN0_6 XI11_0/net21_9_ xsel_42_ XI11_0/XI0/XI0_42/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN0_5 XI11_0/net21_10_ xsel_42_ XI11_0/XI0/XI0_42/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN0_4 XI11_0/net21_11_ xsel_42_ XI11_0/XI0/XI0_42/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN0_3 XI11_0/net21_12_ xsel_42_ XI11_0/XI0/XI0_42/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN0_2 XI11_0/net21_13_ xsel_42_ XI11_0/XI0/XI0_42/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN0_1 XI11_0/net21_14_ xsel_42_ XI11_0/XI0/XI0_42/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN0_0 XI11_0/net21_15_ xsel_42_ XI11_0/XI0/XI0_42/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN1_15 XI11_0/XI0/XI0_42/d__15_ xsel_42_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN1_14 XI11_0/XI0/XI0_42/d__14_ xsel_42_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN1_13 XI11_0/XI0/XI0_42/d__13_ xsel_42_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN1_12 XI11_0/XI0/XI0_42/d__12_ xsel_42_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN1_11 XI11_0/XI0/XI0_42/d__11_ xsel_42_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN1_10 XI11_0/XI0/XI0_42/d__10_ xsel_42_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN1_9 XI11_0/XI0/XI0_42/d__9_ xsel_42_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN1_8 XI11_0/XI0/XI0_42/d__8_ xsel_42_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN1_7 XI11_0/XI0/XI0_42/d__7_ xsel_42_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN1_6 XI11_0/XI0/XI0_42/d__6_ xsel_42_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN1_5 XI11_0/XI0/XI0_42/d__5_ xsel_42_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN1_4 XI11_0/XI0/XI0_42/d__4_ xsel_42_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN1_3 XI11_0/XI0/XI0_42/d__3_ xsel_42_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN1_2 XI11_0/XI0/XI0_42/d__2_ xsel_42_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN1_1 XI11_0/XI0/XI0_42/d__1_ xsel_42_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_42/MN1_0 XI11_0/XI0/XI0_42/d__0_ xsel_42_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN0_15 XI11_0/net21_0_ xsel_41_ XI11_0/XI0/XI0_41/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN0_14 XI11_0/net21_1_ xsel_41_ XI11_0/XI0/XI0_41/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN0_13 XI11_0/net21_2_ xsel_41_ XI11_0/XI0/XI0_41/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN0_12 XI11_0/net21_3_ xsel_41_ XI11_0/XI0/XI0_41/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN0_11 XI11_0/net21_4_ xsel_41_ XI11_0/XI0/XI0_41/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN0_10 XI11_0/net21_5_ xsel_41_ XI11_0/XI0/XI0_41/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN0_9 XI11_0/net21_6_ xsel_41_ XI11_0/XI0/XI0_41/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN0_8 XI11_0/net21_7_ xsel_41_ XI11_0/XI0/XI0_41/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN0_7 XI11_0/net21_8_ xsel_41_ XI11_0/XI0/XI0_41/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN0_6 XI11_0/net21_9_ xsel_41_ XI11_0/XI0/XI0_41/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN0_5 XI11_0/net21_10_ xsel_41_ XI11_0/XI0/XI0_41/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN0_4 XI11_0/net21_11_ xsel_41_ XI11_0/XI0/XI0_41/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN0_3 XI11_0/net21_12_ xsel_41_ XI11_0/XI0/XI0_41/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN0_2 XI11_0/net21_13_ xsel_41_ XI11_0/XI0/XI0_41/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN0_1 XI11_0/net21_14_ xsel_41_ XI11_0/XI0/XI0_41/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN0_0 XI11_0/net21_15_ xsel_41_ XI11_0/XI0/XI0_41/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN1_15 XI11_0/XI0/XI0_41/d__15_ xsel_41_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN1_14 XI11_0/XI0/XI0_41/d__14_ xsel_41_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN1_13 XI11_0/XI0/XI0_41/d__13_ xsel_41_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN1_12 XI11_0/XI0/XI0_41/d__12_ xsel_41_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN1_11 XI11_0/XI0/XI0_41/d__11_ xsel_41_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN1_10 XI11_0/XI0/XI0_41/d__10_ xsel_41_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN1_9 XI11_0/XI0/XI0_41/d__9_ xsel_41_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN1_8 XI11_0/XI0/XI0_41/d__8_ xsel_41_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN1_7 XI11_0/XI0/XI0_41/d__7_ xsel_41_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN1_6 XI11_0/XI0/XI0_41/d__6_ xsel_41_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN1_5 XI11_0/XI0/XI0_41/d__5_ xsel_41_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN1_4 XI11_0/XI0/XI0_41/d__4_ xsel_41_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN1_3 XI11_0/XI0/XI0_41/d__3_ xsel_41_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN1_2 XI11_0/XI0/XI0_41/d__2_ xsel_41_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN1_1 XI11_0/XI0/XI0_41/d__1_ xsel_41_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_41/MN1_0 XI11_0/XI0/XI0_41/d__0_ xsel_41_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN0_15 XI11_0/net21_0_ xsel_40_ XI11_0/XI0/XI0_40/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN0_14 XI11_0/net21_1_ xsel_40_ XI11_0/XI0/XI0_40/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN0_13 XI11_0/net21_2_ xsel_40_ XI11_0/XI0/XI0_40/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN0_12 XI11_0/net21_3_ xsel_40_ XI11_0/XI0/XI0_40/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN0_11 XI11_0/net21_4_ xsel_40_ XI11_0/XI0/XI0_40/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN0_10 XI11_0/net21_5_ xsel_40_ XI11_0/XI0/XI0_40/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN0_9 XI11_0/net21_6_ xsel_40_ XI11_0/XI0/XI0_40/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN0_8 XI11_0/net21_7_ xsel_40_ XI11_0/XI0/XI0_40/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN0_7 XI11_0/net21_8_ xsel_40_ XI11_0/XI0/XI0_40/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN0_6 XI11_0/net21_9_ xsel_40_ XI11_0/XI0/XI0_40/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN0_5 XI11_0/net21_10_ xsel_40_ XI11_0/XI0/XI0_40/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN0_4 XI11_0/net21_11_ xsel_40_ XI11_0/XI0/XI0_40/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN0_3 XI11_0/net21_12_ xsel_40_ XI11_0/XI0/XI0_40/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN0_2 XI11_0/net21_13_ xsel_40_ XI11_0/XI0/XI0_40/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN0_1 XI11_0/net21_14_ xsel_40_ XI11_0/XI0/XI0_40/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN0_0 XI11_0/net21_15_ xsel_40_ XI11_0/XI0/XI0_40/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN1_15 XI11_0/XI0/XI0_40/d__15_ xsel_40_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN1_14 XI11_0/XI0/XI0_40/d__14_ xsel_40_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN1_13 XI11_0/XI0/XI0_40/d__13_ xsel_40_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN1_12 XI11_0/XI0/XI0_40/d__12_ xsel_40_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN1_11 XI11_0/XI0/XI0_40/d__11_ xsel_40_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN1_10 XI11_0/XI0/XI0_40/d__10_ xsel_40_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN1_9 XI11_0/XI0/XI0_40/d__9_ xsel_40_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN1_8 XI11_0/XI0/XI0_40/d__8_ xsel_40_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN1_7 XI11_0/XI0/XI0_40/d__7_ xsel_40_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN1_6 XI11_0/XI0/XI0_40/d__6_ xsel_40_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN1_5 XI11_0/XI0/XI0_40/d__5_ xsel_40_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN1_4 XI11_0/XI0/XI0_40/d__4_ xsel_40_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN1_3 XI11_0/XI0/XI0_40/d__3_ xsel_40_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN1_2 XI11_0/XI0/XI0_40/d__2_ xsel_40_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN1_1 XI11_0/XI0/XI0_40/d__1_ xsel_40_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_40/MN1_0 XI11_0/XI0/XI0_40/d__0_ xsel_40_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN0_15 XI11_0/net21_0_ xsel_39_ XI11_0/XI0/XI0_39/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN0_14 XI11_0/net21_1_ xsel_39_ XI11_0/XI0/XI0_39/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN0_13 XI11_0/net21_2_ xsel_39_ XI11_0/XI0/XI0_39/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN0_12 XI11_0/net21_3_ xsel_39_ XI11_0/XI0/XI0_39/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN0_11 XI11_0/net21_4_ xsel_39_ XI11_0/XI0/XI0_39/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN0_10 XI11_0/net21_5_ xsel_39_ XI11_0/XI0/XI0_39/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN0_9 XI11_0/net21_6_ xsel_39_ XI11_0/XI0/XI0_39/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN0_8 XI11_0/net21_7_ xsel_39_ XI11_0/XI0/XI0_39/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN0_7 XI11_0/net21_8_ xsel_39_ XI11_0/XI0/XI0_39/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN0_6 XI11_0/net21_9_ xsel_39_ XI11_0/XI0/XI0_39/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN0_5 XI11_0/net21_10_ xsel_39_ XI11_0/XI0/XI0_39/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN0_4 XI11_0/net21_11_ xsel_39_ XI11_0/XI0/XI0_39/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN0_3 XI11_0/net21_12_ xsel_39_ XI11_0/XI0/XI0_39/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN0_2 XI11_0/net21_13_ xsel_39_ XI11_0/XI0/XI0_39/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN0_1 XI11_0/net21_14_ xsel_39_ XI11_0/XI0/XI0_39/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN0_0 XI11_0/net21_15_ xsel_39_ XI11_0/XI0/XI0_39/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN1_15 XI11_0/XI0/XI0_39/d__15_ xsel_39_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN1_14 XI11_0/XI0/XI0_39/d__14_ xsel_39_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN1_13 XI11_0/XI0/XI0_39/d__13_ xsel_39_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN1_12 XI11_0/XI0/XI0_39/d__12_ xsel_39_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN1_11 XI11_0/XI0/XI0_39/d__11_ xsel_39_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN1_10 XI11_0/XI0/XI0_39/d__10_ xsel_39_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN1_9 XI11_0/XI0/XI0_39/d__9_ xsel_39_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN1_8 XI11_0/XI0/XI0_39/d__8_ xsel_39_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN1_7 XI11_0/XI0/XI0_39/d__7_ xsel_39_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN1_6 XI11_0/XI0/XI0_39/d__6_ xsel_39_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN1_5 XI11_0/XI0/XI0_39/d__5_ xsel_39_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN1_4 XI11_0/XI0/XI0_39/d__4_ xsel_39_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN1_3 XI11_0/XI0/XI0_39/d__3_ xsel_39_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN1_2 XI11_0/XI0/XI0_39/d__2_ xsel_39_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN1_1 XI11_0/XI0/XI0_39/d__1_ xsel_39_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_39/MN1_0 XI11_0/XI0/XI0_39/d__0_ xsel_39_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN0_15 XI11_0/net21_0_ xsel_38_ XI11_0/XI0/XI0_38/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN0_14 XI11_0/net21_1_ xsel_38_ XI11_0/XI0/XI0_38/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN0_13 XI11_0/net21_2_ xsel_38_ XI11_0/XI0/XI0_38/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN0_12 XI11_0/net21_3_ xsel_38_ XI11_0/XI0/XI0_38/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN0_11 XI11_0/net21_4_ xsel_38_ XI11_0/XI0/XI0_38/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN0_10 XI11_0/net21_5_ xsel_38_ XI11_0/XI0/XI0_38/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN0_9 XI11_0/net21_6_ xsel_38_ XI11_0/XI0/XI0_38/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN0_8 XI11_0/net21_7_ xsel_38_ XI11_0/XI0/XI0_38/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN0_7 XI11_0/net21_8_ xsel_38_ XI11_0/XI0/XI0_38/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN0_6 XI11_0/net21_9_ xsel_38_ XI11_0/XI0/XI0_38/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN0_5 XI11_0/net21_10_ xsel_38_ XI11_0/XI0/XI0_38/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN0_4 XI11_0/net21_11_ xsel_38_ XI11_0/XI0/XI0_38/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN0_3 XI11_0/net21_12_ xsel_38_ XI11_0/XI0/XI0_38/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN0_2 XI11_0/net21_13_ xsel_38_ XI11_0/XI0/XI0_38/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN0_1 XI11_0/net21_14_ xsel_38_ XI11_0/XI0/XI0_38/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN0_0 XI11_0/net21_15_ xsel_38_ XI11_0/XI0/XI0_38/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN1_15 XI11_0/XI0/XI0_38/d__15_ xsel_38_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN1_14 XI11_0/XI0/XI0_38/d__14_ xsel_38_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN1_13 XI11_0/XI0/XI0_38/d__13_ xsel_38_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN1_12 XI11_0/XI0/XI0_38/d__12_ xsel_38_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN1_11 XI11_0/XI0/XI0_38/d__11_ xsel_38_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN1_10 XI11_0/XI0/XI0_38/d__10_ xsel_38_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN1_9 XI11_0/XI0/XI0_38/d__9_ xsel_38_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN1_8 XI11_0/XI0/XI0_38/d__8_ xsel_38_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN1_7 XI11_0/XI0/XI0_38/d__7_ xsel_38_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN1_6 XI11_0/XI0/XI0_38/d__6_ xsel_38_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN1_5 XI11_0/XI0/XI0_38/d__5_ xsel_38_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN1_4 XI11_0/XI0/XI0_38/d__4_ xsel_38_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN1_3 XI11_0/XI0/XI0_38/d__3_ xsel_38_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN1_2 XI11_0/XI0/XI0_38/d__2_ xsel_38_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN1_1 XI11_0/XI0/XI0_38/d__1_ xsel_38_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_38/MN1_0 XI11_0/XI0/XI0_38/d__0_ xsel_38_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN0_15 XI11_0/net21_0_ xsel_37_ XI11_0/XI0/XI0_37/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN0_14 XI11_0/net21_1_ xsel_37_ XI11_0/XI0/XI0_37/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN0_13 XI11_0/net21_2_ xsel_37_ XI11_0/XI0/XI0_37/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN0_12 XI11_0/net21_3_ xsel_37_ XI11_0/XI0/XI0_37/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN0_11 XI11_0/net21_4_ xsel_37_ XI11_0/XI0/XI0_37/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN0_10 XI11_0/net21_5_ xsel_37_ XI11_0/XI0/XI0_37/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN0_9 XI11_0/net21_6_ xsel_37_ XI11_0/XI0/XI0_37/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN0_8 XI11_0/net21_7_ xsel_37_ XI11_0/XI0/XI0_37/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN0_7 XI11_0/net21_8_ xsel_37_ XI11_0/XI0/XI0_37/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN0_6 XI11_0/net21_9_ xsel_37_ XI11_0/XI0/XI0_37/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN0_5 XI11_0/net21_10_ xsel_37_ XI11_0/XI0/XI0_37/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN0_4 XI11_0/net21_11_ xsel_37_ XI11_0/XI0/XI0_37/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN0_3 XI11_0/net21_12_ xsel_37_ XI11_0/XI0/XI0_37/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN0_2 XI11_0/net21_13_ xsel_37_ XI11_0/XI0/XI0_37/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN0_1 XI11_0/net21_14_ xsel_37_ XI11_0/XI0/XI0_37/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN0_0 XI11_0/net21_15_ xsel_37_ XI11_0/XI0/XI0_37/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN1_15 XI11_0/XI0/XI0_37/d__15_ xsel_37_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN1_14 XI11_0/XI0/XI0_37/d__14_ xsel_37_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN1_13 XI11_0/XI0/XI0_37/d__13_ xsel_37_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN1_12 XI11_0/XI0/XI0_37/d__12_ xsel_37_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN1_11 XI11_0/XI0/XI0_37/d__11_ xsel_37_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN1_10 XI11_0/XI0/XI0_37/d__10_ xsel_37_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN1_9 XI11_0/XI0/XI0_37/d__9_ xsel_37_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN1_8 XI11_0/XI0/XI0_37/d__8_ xsel_37_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN1_7 XI11_0/XI0/XI0_37/d__7_ xsel_37_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN1_6 XI11_0/XI0/XI0_37/d__6_ xsel_37_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN1_5 XI11_0/XI0/XI0_37/d__5_ xsel_37_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN1_4 XI11_0/XI0/XI0_37/d__4_ xsel_37_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN1_3 XI11_0/XI0/XI0_37/d__3_ xsel_37_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN1_2 XI11_0/XI0/XI0_37/d__2_ xsel_37_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN1_1 XI11_0/XI0/XI0_37/d__1_ xsel_37_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_37/MN1_0 XI11_0/XI0/XI0_37/d__0_ xsel_37_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN0_15 XI11_0/net21_0_ xsel_36_ XI11_0/XI0/XI0_36/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN0_14 XI11_0/net21_1_ xsel_36_ XI11_0/XI0/XI0_36/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN0_13 XI11_0/net21_2_ xsel_36_ XI11_0/XI0/XI0_36/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN0_12 XI11_0/net21_3_ xsel_36_ XI11_0/XI0/XI0_36/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN0_11 XI11_0/net21_4_ xsel_36_ XI11_0/XI0/XI0_36/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN0_10 XI11_0/net21_5_ xsel_36_ XI11_0/XI0/XI0_36/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN0_9 XI11_0/net21_6_ xsel_36_ XI11_0/XI0/XI0_36/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN0_8 XI11_0/net21_7_ xsel_36_ XI11_0/XI0/XI0_36/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN0_7 XI11_0/net21_8_ xsel_36_ XI11_0/XI0/XI0_36/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN0_6 XI11_0/net21_9_ xsel_36_ XI11_0/XI0/XI0_36/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN0_5 XI11_0/net21_10_ xsel_36_ XI11_0/XI0/XI0_36/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN0_4 XI11_0/net21_11_ xsel_36_ XI11_0/XI0/XI0_36/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN0_3 XI11_0/net21_12_ xsel_36_ XI11_0/XI0/XI0_36/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN0_2 XI11_0/net21_13_ xsel_36_ XI11_0/XI0/XI0_36/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN0_1 XI11_0/net21_14_ xsel_36_ XI11_0/XI0/XI0_36/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN0_0 XI11_0/net21_15_ xsel_36_ XI11_0/XI0/XI0_36/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN1_15 XI11_0/XI0/XI0_36/d__15_ xsel_36_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN1_14 XI11_0/XI0/XI0_36/d__14_ xsel_36_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN1_13 XI11_0/XI0/XI0_36/d__13_ xsel_36_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN1_12 XI11_0/XI0/XI0_36/d__12_ xsel_36_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN1_11 XI11_0/XI0/XI0_36/d__11_ xsel_36_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN1_10 XI11_0/XI0/XI0_36/d__10_ xsel_36_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN1_9 XI11_0/XI0/XI0_36/d__9_ xsel_36_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN1_8 XI11_0/XI0/XI0_36/d__8_ xsel_36_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN1_7 XI11_0/XI0/XI0_36/d__7_ xsel_36_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN1_6 XI11_0/XI0/XI0_36/d__6_ xsel_36_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN1_5 XI11_0/XI0/XI0_36/d__5_ xsel_36_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN1_4 XI11_0/XI0/XI0_36/d__4_ xsel_36_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN1_3 XI11_0/XI0/XI0_36/d__3_ xsel_36_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN1_2 XI11_0/XI0/XI0_36/d__2_ xsel_36_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN1_1 XI11_0/XI0/XI0_36/d__1_ xsel_36_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_36/MN1_0 XI11_0/XI0/XI0_36/d__0_ xsel_36_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN0_15 XI11_0/net21_0_ xsel_35_ XI11_0/XI0/XI0_35/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN0_14 XI11_0/net21_1_ xsel_35_ XI11_0/XI0/XI0_35/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN0_13 XI11_0/net21_2_ xsel_35_ XI11_0/XI0/XI0_35/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN0_12 XI11_0/net21_3_ xsel_35_ XI11_0/XI0/XI0_35/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN0_11 XI11_0/net21_4_ xsel_35_ XI11_0/XI0/XI0_35/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN0_10 XI11_0/net21_5_ xsel_35_ XI11_0/XI0/XI0_35/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN0_9 XI11_0/net21_6_ xsel_35_ XI11_0/XI0/XI0_35/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN0_8 XI11_0/net21_7_ xsel_35_ XI11_0/XI0/XI0_35/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN0_7 XI11_0/net21_8_ xsel_35_ XI11_0/XI0/XI0_35/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN0_6 XI11_0/net21_9_ xsel_35_ XI11_0/XI0/XI0_35/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN0_5 XI11_0/net21_10_ xsel_35_ XI11_0/XI0/XI0_35/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN0_4 XI11_0/net21_11_ xsel_35_ XI11_0/XI0/XI0_35/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN0_3 XI11_0/net21_12_ xsel_35_ XI11_0/XI0/XI0_35/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN0_2 XI11_0/net21_13_ xsel_35_ XI11_0/XI0/XI0_35/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN0_1 XI11_0/net21_14_ xsel_35_ XI11_0/XI0/XI0_35/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN0_0 XI11_0/net21_15_ xsel_35_ XI11_0/XI0/XI0_35/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN1_15 XI11_0/XI0/XI0_35/d__15_ xsel_35_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN1_14 XI11_0/XI0/XI0_35/d__14_ xsel_35_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN1_13 XI11_0/XI0/XI0_35/d__13_ xsel_35_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN1_12 XI11_0/XI0/XI0_35/d__12_ xsel_35_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN1_11 XI11_0/XI0/XI0_35/d__11_ xsel_35_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN1_10 XI11_0/XI0/XI0_35/d__10_ xsel_35_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN1_9 XI11_0/XI0/XI0_35/d__9_ xsel_35_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN1_8 XI11_0/XI0/XI0_35/d__8_ xsel_35_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN1_7 XI11_0/XI0/XI0_35/d__7_ xsel_35_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN1_6 XI11_0/XI0/XI0_35/d__6_ xsel_35_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN1_5 XI11_0/XI0/XI0_35/d__5_ xsel_35_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN1_4 XI11_0/XI0/XI0_35/d__4_ xsel_35_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN1_3 XI11_0/XI0/XI0_35/d__3_ xsel_35_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN1_2 XI11_0/XI0/XI0_35/d__2_ xsel_35_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN1_1 XI11_0/XI0/XI0_35/d__1_ xsel_35_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_35/MN1_0 XI11_0/XI0/XI0_35/d__0_ xsel_35_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN0_15 XI11_0/net21_0_ xsel_34_ XI11_0/XI0/XI0_34/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN0_14 XI11_0/net21_1_ xsel_34_ XI11_0/XI0/XI0_34/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN0_13 XI11_0/net21_2_ xsel_34_ XI11_0/XI0/XI0_34/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN0_12 XI11_0/net21_3_ xsel_34_ XI11_0/XI0/XI0_34/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN0_11 XI11_0/net21_4_ xsel_34_ XI11_0/XI0/XI0_34/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN0_10 XI11_0/net21_5_ xsel_34_ XI11_0/XI0/XI0_34/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN0_9 XI11_0/net21_6_ xsel_34_ XI11_0/XI0/XI0_34/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN0_8 XI11_0/net21_7_ xsel_34_ XI11_0/XI0/XI0_34/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN0_7 XI11_0/net21_8_ xsel_34_ XI11_0/XI0/XI0_34/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN0_6 XI11_0/net21_9_ xsel_34_ XI11_0/XI0/XI0_34/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN0_5 XI11_0/net21_10_ xsel_34_ XI11_0/XI0/XI0_34/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN0_4 XI11_0/net21_11_ xsel_34_ XI11_0/XI0/XI0_34/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN0_3 XI11_0/net21_12_ xsel_34_ XI11_0/XI0/XI0_34/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN0_2 XI11_0/net21_13_ xsel_34_ XI11_0/XI0/XI0_34/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN0_1 XI11_0/net21_14_ xsel_34_ XI11_0/XI0/XI0_34/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN0_0 XI11_0/net21_15_ xsel_34_ XI11_0/XI0/XI0_34/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN1_15 XI11_0/XI0/XI0_34/d__15_ xsel_34_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN1_14 XI11_0/XI0/XI0_34/d__14_ xsel_34_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN1_13 XI11_0/XI0/XI0_34/d__13_ xsel_34_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN1_12 XI11_0/XI0/XI0_34/d__12_ xsel_34_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN1_11 XI11_0/XI0/XI0_34/d__11_ xsel_34_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN1_10 XI11_0/XI0/XI0_34/d__10_ xsel_34_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN1_9 XI11_0/XI0/XI0_34/d__9_ xsel_34_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN1_8 XI11_0/XI0/XI0_34/d__8_ xsel_34_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN1_7 XI11_0/XI0/XI0_34/d__7_ xsel_34_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN1_6 XI11_0/XI0/XI0_34/d__6_ xsel_34_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN1_5 XI11_0/XI0/XI0_34/d__5_ xsel_34_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN1_4 XI11_0/XI0/XI0_34/d__4_ xsel_34_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN1_3 XI11_0/XI0/XI0_34/d__3_ xsel_34_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN1_2 XI11_0/XI0/XI0_34/d__2_ xsel_34_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN1_1 XI11_0/XI0/XI0_34/d__1_ xsel_34_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_34/MN1_0 XI11_0/XI0/XI0_34/d__0_ xsel_34_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN0_15 XI11_0/net21_0_ xsel_33_ XI11_0/XI0/XI0_33/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN0_14 XI11_0/net21_1_ xsel_33_ XI11_0/XI0/XI0_33/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN0_13 XI11_0/net21_2_ xsel_33_ XI11_0/XI0/XI0_33/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN0_12 XI11_0/net21_3_ xsel_33_ XI11_0/XI0/XI0_33/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN0_11 XI11_0/net21_4_ xsel_33_ XI11_0/XI0/XI0_33/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN0_10 XI11_0/net21_5_ xsel_33_ XI11_0/XI0/XI0_33/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN0_9 XI11_0/net21_6_ xsel_33_ XI11_0/XI0/XI0_33/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN0_8 XI11_0/net21_7_ xsel_33_ XI11_0/XI0/XI0_33/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN0_7 XI11_0/net21_8_ xsel_33_ XI11_0/XI0/XI0_33/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN0_6 XI11_0/net21_9_ xsel_33_ XI11_0/XI0/XI0_33/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN0_5 XI11_0/net21_10_ xsel_33_ XI11_0/XI0/XI0_33/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN0_4 XI11_0/net21_11_ xsel_33_ XI11_0/XI0/XI0_33/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN0_3 XI11_0/net21_12_ xsel_33_ XI11_0/XI0/XI0_33/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN0_2 XI11_0/net21_13_ xsel_33_ XI11_0/XI0/XI0_33/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN0_1 XI11_0/net21_14_ xsel_33_ XI11_0/XI0/XI0_33/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN0_0 XI11_0/net21_15_ xsel_33_ XI11_0/XI0/XI0_33/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN1_15 XI11_0/XI0/XI0_33/d__15_ xsel_33_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN1_14 XI11_0/XI0/XI0_33/d__14_ xsel_33_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN1_13 XI11_0/XI0/XI0_33/d__13_ xsel_33_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN1_12 XI11_0/XI0/XI0_33/d__12_ xsel_33_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN1_11 XI11_0/XI0/XI0_33/d__11_ xsel_33_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN1_10 XI11_0/XI0/XI0_33/d__10_ xsel_33_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN1_9 XI11_0/XI0/XI0_33/d__9_ xsel_33_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN1_8 XI11_0/XI0/XI0_33/d__8_ xsel_33_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN1_7 XI11_0/XI0/XI0_33/d__7_ xsel_33_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN1_6 XI11_0/XI0/XI0_33/d__6_ xsel_33_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN1_5 XI11_0/XI0/XI0_33/d__5_ xsel_33_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN1_4 XI11_0/XI0/XI0_33/d__4_ xsel_33_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN1_3 XI11_0/XI0/XI0_33/d__3_ xsel_33_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN1_2 XI11_0/XI0/XI0_33/d__2_ xsel_33_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN1_1 XI11_0/XI0/XI0_33/d__1_ xsel_33_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_33/MN1_0 XI11_0/XI0/XI0_33/d__0_ xsel_33_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN0_15 XI11_0/net21_0_ xsel_32_ XI11_0/XI0/XI0_32/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN0_14 XI11_0/net21_1_ xsel_32_ XI11_0/XI0/XI0_32/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN0_13 XI11_0/net21_2_ xsel_32_ XI11_0/XI0/XI0_32/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN0_12 XI11_0/net21_3_ xsel_32_ XI11_0/XI0/XI0_32/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN0_11 XI11_0/net21_4_ xsel_32_ XI11_0/XI0/XI0_32/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN0_10 XI11_0/net21_5_ xsel_32_ XI11_0/XI0/XI0_32/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN0_9 XI11_0/net21_6_ xsel_32_ XI11_0/XI0/XI0_32/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN0_8 XI11_0/net21_7_ xsel_32_ XI11_0/XI0/XI0_32/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN0_7 XI11_0/net21_8_ xsel_32_ XI11_0/XI0/XI0_32/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN0_6 XI11_0/net21_9_ xsel_32_ XI11_0/XI0/XI0_32/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN0_5 XI11_0/net21_10_ xsel_32_ XI11_0/XI0/XI0_32/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN0_4 XI11_0/net21_11_ xsel_32_ XI11_0/XI0/XI0_32/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN0_3 XI11_0/net21_12_ xsel_32_ XI11_0/XI0/XI0_32/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN0_2 XI11_0/net21_13_ xsel_32_ XI11_0/XI0/XI0_32/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN0_1 XI11_0/net21_14_ xsel_32_ XI11_0/XI0/XI0_32/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN0_0 XI11_0/net21_15_ xsel_32_ XI11_0/XI0/XI0_32/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN1_15 XI11_0/XI0/XI0_32/d__15_ xsel_32_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN1_14 XI11_0/XI0/XI0_32/d__14_ xsel_32_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN1_13 XI11_0/XI0/XI0_32/d__13_ xsel_32_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN1_12 XI11_0/XI0/XI0_32/d__12_ xsel_32_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN1_11 XI11_0/XI0/XI0_32/d__11_ xsel_32_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN1_10 XI11_0/XI0/XI0_32/d__10_ xsel_32_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN1_9 XI11_0/XI0/XI0_32/d__9_ xsel_32_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN1_8 XI11_0/XI0/XI0_32/d__8_ xsel_32_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN1_7 XI11_0/XI0/XI0_32/d__7_ xsel_32_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN1_6 XI11_0/XI0/XI0_32/d__6_ xsel_32_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN1_5 XI11_0/XI0/XI0_32/d__5_ xsel_32_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN1_4 XI11_0/XI0/XI0_32/d__4_ xsel_32_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN1_3 XI11_0/XI0/XI0_32/d__3_ xsel_32_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN1_2 XI11_0/XI0/XI0_32/d__2_ xsel_32_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN1_1 XI11_0/XI0/XI0_32/d__1_ xsel_32_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_32/MN1_0 XI11_0/XI0/XI0_32/d__0_ xsel_32_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN0_15 XI11_0/net21_0_ xsel_31_ XI11_0/XI0/XI0_31/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN0_14 XI11_0/net21_1_ xsel_31_ XI11_0/XI0/XI0_31/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN0_13 XI11_0/net21_2_ xsel_31_ XI11_0/XI0/XI0_31/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN0_12 XI11_0/net21_3_ xsel_31_ XI11_0/XI0/XI0_31/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN0_11 XI11_0/net21_4_ xsel_31_ XI11_0/XI0/XI0_31/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN0_10 XI11_0/net21_5_ xsel_31_ XI11_0/XI0/XI0_31/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN0_9 XI11_0/net21_6_ xsel_31_ XI11_0/XI0/XI0_31/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN0_8 XI11_0/net21_7_ xsel_31_ XI11_0/XI0/XI0_31/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN0_7 XI11_0/net21_8_ xsel_31_ XI11_0/XI0/XI0_31/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN0_6 XI11_0/net21_9_ xsel_31_ XI11_0/XI0/XI0_31/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN0_5 XI11_0/net21_10_ xsel_31_ XI11_0/XI0/XI0_31/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN0_4 XI11_0/net21_11_ xsel_31_ XI11_0/XI0/XI0_31/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN0_3 XI11_0/net21_12_ xsel_31_ XI11_0/XI0/XI0_31/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN0_2 XI11_0/net21_13_ xsel_31_ XI11_0/XI0/XI0_31/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN0_1 XI11_0/net21_14_ xsel_31_ XI11_0/XI0/XI0_31/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN0_0 XI11_0/net21_15_ xsel_31_ XI11_0/XI0/XI0_31/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN1_15 XI11_0/XI0/XI0_31/d__15_ xsel_31_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN1_14 XI11_0/XI0/XI0_31/d__14_ xsel_31_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN1_13 XI11_0/XI0/XI0_31/d__13_ xsel_31_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN1_12 XI11_0/XI0/XI0_31/d__12_ xsel_31_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN1_11 XI11_0/XI0/XI0_31/d__11_ xsel_31_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN1_10 XI11_0/XI0/XI0_31/d__10_ xsel_31_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN1_9 XI11_0/XI0/XI0_31/d__9_ xsel_31_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN1_8 XI11_0/XI0/XI0_31/d__8_ xsel_31_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN1_7 XI11_0/XI0/XI0_31/d__7_ xsel_31_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN1_6 XI11_0/XI0/XI0_31/d__6_ xsel_31_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN1_5 XI11_0/XI0/XI0_31/d__5_ xsel_31_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN1_4 XI11_0/XI0/XI0_31/d__4_ xsel_31_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN1_3 XI11_0/XI0/XI0_31/d__3_ xsel_31_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN1_2 XI11_0/XI0/XI0_31/d__2_ xsel_31_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN1_1 XI11_0/XI0/XI0_31/d__1_ xsel_31_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_31/MN1_0 XI11_0/XI0/XI0_31/d__0_ xsel_31_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN0_15 XI11_0/net21_0_ xsel_30_ XI11_0/XI0/XI0_30/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN0_14 XI11_0/net21_1_ xsel_30_ XI11_0/XI0/XI0_30/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN0_13 XI11_0/net21_2_ xsel_30_ XI11_0/XI0/XI0_30/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN0_12 XI11_0/net21_3_ xsel_30_ XI11_0/XI0/XI0_30/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN0_11 XI11_0/net21_4_ xsel_30_ XI11_0/XI0/XI0_30/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN0_10 XI11_0/net21_5_ xsel_30_ XI11_0/XI0/XI0_30/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN0_9 XI11_0/net21_6_ xsel_30_ XI11_0/XI0/XI0_30/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN0_8 XI11_0/net21_7_ xsel_30_ XI11_0/XI0/XI0_30/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN0_7 XI11_0/net21_8_ xsel_30_ XI11_0/XI0/XI0_30/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN0_6 XI11_0/net21_9_ xsel_30_ XI11_0/XI0/XI0_30/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN0_5 XI11_0/net21_10_ xsel_30_ XI11_0/XI0/XI0_30/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN0_4 XI11_0/net21_11_ xsel_30_ XI11_0/XI0/XI0_30/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN0_3 XI11_0/net21_12_ xsel_30_ XI11_0/XI0/XI0_30/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN0_2 XI11_0/net21_13_ xsel_30_ XI11_0/XI0/XI0_30/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN0_1 XI11_0/net21_14_ xsel_30_ XI11_0/XI0/XI0_30/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN0_0 XI11_0/net21_15_ xsel_30_ XI11_0/XI0/XI0_30/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN1_15 XI11_0/XI0/XI0_30/d__15_ xsel_30_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN1_14 XI11_0/XI0/XI0_30/d__14_ xsel_30_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN1_13 XI11_0/XI0/XI0_30/d__13_ xsel_30_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN1_12 XI11_0/XI0/XI0_30/d__12_ xsel_30_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN1_11 XI11_0/XI0/XI0_30/d__11_ xsel_30_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN1_10 XI11_0/XI0/XI0_30/d__10_ xsel_30_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN1_9 XI11_0/XI0/XI0_30/d__9_ xsel_30_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN1_8 XI11_0/XI0/XI0_30/d__8_ xsel_30_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN1_7 XI11_0/XI0/XI0_30/d__7_ xsel_30_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN1_6 XI11_0/XI0/XI0_30/d__6_ xsel_30_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN1_5 XI11_0/XI0/XI0_30/d__5_ xsel_30_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN1_4 XI11_0/XI0/XI0_30/d__4_ xsel_30_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN1_3 XI11_0/XI0/XI0_30/d__3_ xsel_30_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN1_2 XI11_0/XI0/XI0_30/d__2_ xsel_30_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN1_1 XI11_0/XI0/XI0_30/d__1_ xsel_30_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_30/MN1_0 XI11_0/XI0/XI0_30/d__0_ xsel_30_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN0_15 XI11_0/net21_0_ xsel_29_ XI11_0/XI0/XI0_29/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN0_14 XI11_0/net21_1_ xsel_29_ XI11_0/XI0/XI0_29/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN0_13 XI11_0/net21_2_ xsel_29_ XI11_0/XI0/XI0_29/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN0_12 XI11_0/net21_3_ xsel_29_ XI11_0/XI0/XI0_29/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN0_11 XI11_0/net21_4_ xsel_29_ XI11_0/XI0/XI0_29/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN0_10 XI11_0/net21_5_ xsel_29_ XI11_0/XI0/XI0_29/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN0_9 XI11_0/net21_6_ xsel_29_ XI11_0/XI0/XI0_29/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN0_8 XI11_0/net21_7_ xsel_29_ XI11_0/XI0/XI0_29/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN0_7 XI11_0/net21_8_ xsel_29_ XI11_0/XI0/XI0_29/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN0_6 XI11_0/net21_9_ xsel_29_ XI11_0/XI0/XI0_29/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN0_5 XI11_0/net21_10_ xsel_29_ XI11_0/XI0/XI0_29/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN0_4 XI11_0/net21_11_ xsel_29_ XI11_0/XI0/XI0_29/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN0_3 XI11_0/net21_12_ xsel_29_ XI11_0/XI0/XI0_29/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN0_2 XI11_0/net21_13_ xsel_29_ XI11_0/XI0/XI0_29/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN0_1 XI11_0/net21_14_ xsel_29_ XI11_0/XI0/XI0_29/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN0_0 XI11_0/net21_15_ xsel_29_ XI11_0/XI0/XI0_29/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN1_15 XI11_0/XI0/XI0_29/d__15_ xsel_29_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN1_14 XI11_0/XI0/XI0_29/d__14_ xsel_29_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN1_13 XI11_0/XI0/XI0_29/d__13_ xsel_29_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN1_12 XI11_0/XI0/XI0_29/d__12_ xsel_29_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN1_11 XI11_0/XI0/XI0_29/d__11_ xsel_29_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN1_10 XI11_0/XI0/XI0_29/d__10_ xsel_29_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN1_9 XI11_0/XI0/XI0_29/d__9_ xsel_29_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN1_8 XI11_0/XI0/XI0_29/d__8_ xsel_29_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN1_7 XI11_0/XI0/XI0_29/d__7_ xsel_29_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN1_6 XI11_0/XI0/XI0_29/d__6_ xsel_29_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN1_5 XI11_0/XI0/XI0_29/d__5_ xsel_29_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN1_4 XI11_0/XI0/XI0_29/d__4_ xsel_29_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN1_3 XI11_0/XI0/XI0_29/d__3_ xsel_29_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN1_2 XI11_0/XI0/XI0_29/d__2_ xsel_29_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN1_1 XI11_0/XI0/XI0_29/d__1_ xsel_29_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_29/MN1_0 XI11_0/XI0/XI0_29/d__0_ xsel_29_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN0_15 XI11_0/net21_0_ xsel_28_ XI11_0/XI0/XI0_28/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN0_14 XI11_0/net21_1_ xsel_28_ XI11_0/XI0/XI0_28/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN0_13 XI11_0/net21_2_ xsel_28_ XI11_0/XI0/XI0_28/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN0_12 XI11_0/net21_3_ xsel_28_ XI11_0/XI0/XI0_28/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN0_11 XI11_0/net21_4_ xsel_28_ XI11_0/XI0/XI0_28/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN0_10 XI11_0/net21_5_ xsel_28_ XI11_0/XI0/XI0_28/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN0_9 XI11_0/net21_6_ xsel_28_ XI11_0/XI0/XI0_28/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN0_8 XI11_0/net21_7_ xsel_28_ XI11_0/XI0/XI0_28/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN0_7 XI11_0/net21_8_ xsel_28_ XI11_0/XI0/XI0_28/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN0_6 XI11_0/net21_9_ xsel_28_ XI11_0/XI0/XI0_28/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN0_5 XI11_0/net21_10_ xsel_28_ XI11_0/XI0/XI0_28/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN0_4 XI11_0/net21_11_ xsel_28_ XI11_0/XI0/XI0_28/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN0_3 XI11_0/net21_12_ xsel_28_ XI11_0/XI0/XI0_28/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN0_2 XI11_0/net21_13_ xsel_28_ XI11_0/XI0/XI0_28/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN0_1 XI11_0/net21_14_ xsel_28_ XI11_0/XI0/XI0_28/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN0_0 XI11_0/net21_15_ xsel_28_ XI11_0/XI0/XI0_28/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN1_15 XI11_0/XI0/XI0_28/d__15_ xsel_28_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN1_14 XI11_0/XI0/XI0_28/d__14_ xsel_28_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN1_13 XI11_0/XI0/XI0_28/d__13_ xsel_28_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN1_12 XI11_0/XI0/XI0_28/d__12_ xsel_28_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN1_11 XI11_0/XI0/XI0_28/d__11_ xsel_28_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN1_10 XI11_0/XI0/XI0_28/d__10_ xsel_28_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN1_9 XI11_0/XI0/XI0_28/d__9_ xsel_28_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN1_8 XI11_0/XI0/XI0_28/d__8_ xsel_28_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN1_7 XI11_0/XI0/XI0_28/d__7_ xsel_28_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN1_6 XI11_0/XI0/XI0_28/d__6_ xsel_28_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN1_5 XI11_0/XI0/XI0_28/d__5_ xsel_28_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN1_4 XI11_0/XI0/XI0_28/d__4_ xsel_28_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN1_3 XI11_0/XI0/XI0_28/d__3_ xsel_28_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN1_2 XI11_0/XI0/XI0_28/d__2_ xsel_28_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN1_1 XI11_0/XI0/XI0_28/d__1_ xsel_28_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_28/MN1_0 XI11_0/XI0/XI0_28/d__0_ xsel_28_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN0_15 XI11_0/net21_0_ xsel_27_ XI11_0/XI0/XI0_27/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN0_14 XI11_0/net21_1_ xsel_27_ XI11_0/XI0/XI0_27/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN0_13 XI11_0/net21_2_ xsel_27_ XI11_0/XI0/XI0_27/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN0_12 XI11_0/net21_3_ xsel_27_ XI11_0/XI0/XI0_27/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN0_11 XI11_0/net21_4_ xsel_27_ XI11_0/XI0/XI0_27/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN0_10 XI11_0/net21_5_ xsel_27_ XI11_0/XI0/XI0_27/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN0_9 XI11_0/net21_6_ xsel_27_ XI11_0/XI0/XI0_27/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN0_8 XI11_0/net21_7_ xsel_27_ XI11_0/XI0/XI0_27/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN0_7 XI11_0/net21_8_ xsel_27_ XI11_0/XI0/XI0_27/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN0_6 XI11_0/net21_9_ xsel_27_ XI11_0/XI0/XI0_27/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN0_5 XI11_0/net21_10_ xsel_27_ XI11_0/XI0/XI0_27/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN0_4 XI11_0/net21_11_ xsel_27_ XI11_0/XI0/XI0_27/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN0_3 XI11_0/net21_12_ xsel_27_ XI11_0/XI0/XI0_27/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN0_2 XI11_0/net21_13_ xsel_27_ XI11_0/XI0/XI0_27/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN0_1 XI11_0/net21_14_ xsel_27_ XI11_0/XI0/XI0_27/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN0_0 XI11_0/net21_15_ xsel_27_ XI11_0/XI0/XI0_27/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN1_15 XI11_0/XI0/XI0_27/d__15_ xsel_27_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN1_14 XI11_0/XI0/XI0_27/d__14_ xsel_27_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN1_13 XI11_0/XI0/XI0_27/d__13_ xsel_27_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN1_12 XI11_0/XI0/XI0_27/d__12_ xsel_27_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN1_11 XI11_0/XI0/XI0_27/d__11_ xsel_27_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN1_10 XI11_0/XI0/XI0_27/d__10_ xsel_27_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN1_9 XI11_0/XI0/XI0_27/d__9_ xsel_27_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN1_8 XI11_0/XI0/XI0_27/d__8_ xsel_27_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN1_7 XI11_0/XI0/XI0_27/d__7_ xsel_27_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN1_6 XI11_0/XI0/XI0_27/d__6_ xsel_27_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN1_5 XI11_0/XI0/XI0_27/d__5_ xsel_27_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN1_4 XI11_0/XI0/XI0_27/d__4_ xsel_27_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN1_3 XI11_0/XI0/XI0_27/d__3_ xsel_27_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN1_2 XI11_0/XI0/XI0_27/d__2_ xsel_27_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN1_1 XI11_0/XI0/XI0_27/d__1_ xsel_27_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_27/MN1_0 XI11_0/XI0/XI0_27/d__0_ xsel_27_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN0_15 XI11_0/net21_0_ xsel_26_ XI11_0/XI0/XI0_26/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN0_14 XI11_0/net21_1_ xsel_26_ XI11_0/XI0/XI0_26/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN0_13 XI11_0/net21_2_ xsel_26_ XI11_0/XI0/XI0_26/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN0_12 XI11_0/net21_3_ xsel_26_ XI11_0/XI0/XI0_26/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN0_11 XI11_0/net21_4_ xsel_26_ XI11_0/XI0/XI0_26/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN0_10 XI11_0/net21_5_ xsel_26_ XI11_0/XI0/XI0_26/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN0_9 XI11_0/net21_6_ xsel_26_ XI11_0/XI0/XI0_26/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN0_8 XI11_0/net21_7_ xsel_26_ XI11_0/XI0/XI0_26/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN0_7 XI11_0/net21_8_ xsel_26_ XI11_0/XI0/XI0_26/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN0_6 XI11_0/net21_9_ xsel_26_ XI11_0/XI0/XI0_26/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN0_5 XI11_0/net21_10_ xsel_26_ XI11_0/XI0/XI0_26/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN0_4 XI11_0/net21_11_ xsel_26_ XI11_0/XI0/XI0_26/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN0_3 XI11_0/net21_12_ xsel_26_ XI11_0/XI0/XI0_26/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN0_2 XI11_0/net21_13_ xsel_26_ XI11_0/XI0/XI0_26/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN0_1 XI11_0/net21_14_ xsel_26_ XI11_0/XI0/XI0_26/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN0_0 XI11_0/net21_15_ xsel_26_ XI11_0/XI0/XI0_26/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN1_15 XI11_0/XI0/XI0_26/d__15_ xsel_26_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN1_14 XI11_0/XI0/XI0_26/d__14_ xsel_26_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN1_13 XI11_0/XI0/XI0_26/d__13_ xsel_26_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN1_12 XI11_0/XI0/XI0_26/d__12_ xsel_26_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN1_11 XI11_0/XI0/XI0_26/d__11_ xsel_26_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN1_10 XI11_0/XI0/XI0_26/d__10_ xsel_26_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN1_9 XI11_0/XI0/XI0_26/d__9_ xsel_26_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN1_8 XI11_0/XI0/XI0_26/d__8_ xsel_26_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN1_7 XI11_0/XI0/XI0_26/d__7_ xsel_26_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN1_6 XI11_0/XI0/XI0_26/d__6_ xsel_26_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN1_5 XI11_0/XI0/XI0_26/d__5_ xsel_26_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN1_4 XI11_0/XI0/XI0_26/d__4_ xsel_26_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN1_3 XI11_0/XI0/XI0_26/d__3_ xsel_26_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN1_2 XI11_0/XI0/XI0_26/d__2_ xsel_26_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN1_1 XI11_0/XI0/XI0_26/d__1_ xsel_26_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_26/MN1_0 XI11_0/XI0/XI0_26/d__0_ xsel_26_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN0_15 XI11_0/net21_0_ xsel_25_ XI11_0/XI0/XI0_25/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN0_14 XI11_0/net21_1_ xsel_25_ XI11_0/XI0/XI0_25/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN0_13 XI11_0/net21_2_ xsel_25_ XI11_0/XI0/XI0_25/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN0_12 XI11_0/net21_3_ xsel_25_ XI11_0/XI0/XI0_25/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN0_11 XI11_0/net21_4_ xsel_25_ XI11_0/XI0/XI0_25/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN0_10 XI11_0/net21_5_ xsel_25_ XI11_0/XI0/XI0_25/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN0_9 XI11_0/net21_6_ xsel_25_ XI11_0/XI0/XI0_25/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN0_8 XI11_0/net21_7_ xsel_25_ XI11_0/XI0/XI0_25/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN0_7 XI11_0/net21_8_ xsel_25_ XI11_0/XI0/XI0_25/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN0_6 XI11_0/net21_9_ xsel_25_ XI11_0/XI0/XI0_25/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN0_5 XI11_0/net21_10_ xsel_25_ XI11_0/XI0/XI0_25/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN0_4 XI11_0/net21_11_ xsel_25_ XI11_0/XI0/XI0_25/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN0_3 XI11_0/net21_12_ xsel_25_ XI11_0/XI0/XI0_25/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN0_2 XI11_0/net21_13_ xsel_25_ XI11_0/XI0/XI0_25/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN0_1 XI11_0/net21_14_ xsel_25_ XI11_0/XI0/XI0_25/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN0_0 XI11_0/net21_15_ xsel_25_ XI11_0/XI0/XI0_25/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN1_15 XI11_0/XI0/XI0_25/d__15_ xsel_25_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN1_14 XI11_0/XI0/XI0_25/d__14_ xsel_25_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN1_13 XI11_0/XI0/XI0_25/d__13_ xsel_25_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN1_12 XI11_0/XI0/XI0_25/d__12_ xsel_25_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN1_11 XI11_0/XI0/XI0_25/d__11_ xsel_25_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN1_10 XI11_0/XI0/XI0_25/d__10_ xsel_25_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN1_9 XI11_0/XI0/XI0_25/d__9_ xsel_25_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN1_8 XI11_0/XI0/XI0_25/d__8_ xsel_25_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN1_7 XI11_0/XI0/XI0_25/d__7_ xsel_25_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN1_6 XI11_0/XI0/XI0_25/d__6_ xsel_25_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN1_5 XI11_0/XI0/XI0_25/d__5_ xsel_25_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN1_4 XI11_0/XI0/XI0_25/d__4_ xsel_25_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN1_3 XI11_0/XI0/XI0_25/d__3_ xsel_25_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN1_2 XI11_0/XI0/XI0_25/d__2_ xsel_25_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN1_1 XI11_0/XI0/XI0_25/d__1_ xsel_25_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_25/MN1_0 XI11_0/XI0/XI0_25/d__0_ xsel_25_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN0_15 XI11_0/net21_0_ xsel_24_ XI11_0/XI0/XI0_24/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN0_14 XI11_0/net21_1_ xsel_24_ XI11_0/XI0/XI0_24/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN0_13 XI11_0/net21_2_ xsel_24_ XI11_0/XI0/XI0_24/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN0_12 XI11_0/net21_3_ xsel_24_ XI11_0/XI0/XI0_24/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN0_11 XI11_0/net21_4_ xsel_24_ XI11_0/XI0/XI0_24/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN0_10 XI11_0/net21_5_ xsel_24_ XI11_0/XI0/XI0_24/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN0_9 XI11_0/net21_6_ xsel_24_ XI11_0/XI0/XI0_24/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN0_8 XI11_0/net21_7_ xsel_24_ XI11_0/XI0/XI0_24/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN0_7 XI11_0/net21_8_ xsel_24_ XI11_0/XI0/XI0_24/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN0_6 XI11_0/net21_9_ xsel_24_ XI11_0/XI0/XI0_24/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN0_5 XI11_0/net21_10_ xsel_24_ XI11_0/XI0/XI0_24/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN0_4 XI11_0/net21_11_ xsel_24_ XI11_0/XI0/XI0_24/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN0_3 XI11_0/net21_12_ xsel_24_ XI11_0/XI0/XI0_24/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN0_2 XI11_0/net21_13_ xsel_24_ XI11_0/XI0/XI0_24/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN0_1 XI11_0/net21_14_ xsel_24_ XI11_0/XI0/XI0_24/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN0_0 XI11_0/net21_15_ xsel_24_ XI11_0/XI0/XI0_24/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN1_15 XI11_0/XI0/XI0_24/d__15_ xsel_24_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN1_14 XI11_0/XI0/XI0_24/d__14_ xsel_24_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN1_13 XI11_0/XI0/XI0_24/d__13_ xsel_24_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN1_12 XI11_0/XI0/XI0_24/d__12_ xsel_24_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN1_11 XI11_0/XI0/XI0_24/d__11_ xsel_24_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN1_10 XI11_0/XI0/XI0_24/d__10_ xsel_24_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN1_9 XI11_0/XI0/XI0_24/d__9_ xsel_24_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN1_8 XI11_0/XI0/XI0_24/d__8_ xsel_24_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN1_7 XI11_0/XI0/XI0_24/d__7_ xsel_24_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN1_6 XI11_0/XI0/XI0_24/d__6_ xsel_24_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN1_5 XI11_0/XI0/XI0_24/d__5_ xsel_24_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN1_4 XI11_0/XI0/XI0_24/d__4_ xsel_24_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN1_3 XI11_0/XI0/XI0_24/d__3_ xsel_24_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN1_2 XI11_0/XI0/XI0_24/d__2_ xsel_24_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN1_1 XI11_0/XI0/XI0_24/d__1_ xsel_24_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_24/MN1_0 XI11_0/XI0/XI0_24/d__0_ xsel_24_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN0_15 XI11_0/net21_0_ xsel_23_ XI11_0/XI0/XI0_23/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN0_14 XI11_0/net21_1_ xsel_23_ XI11_0/XI0/XI0_23/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN0_13 XI11_0/net21_2_ xsel_23_ XI11_0/XI0/XI0_23/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN0_12 XI11_0/net21_3_ xsel_23_ XI11_0/XI0/XI0_23/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN0_11 XI11_0/net21_4_ xsel_23_ XI11_0/XI0/XI0_23/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN0_10 XI11_0/net21_5_ xsel_23_ XI11_0/XI0/XI0_23/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN0_9 XI11_0/net21_6_ xsel_23_ XI11_0/XI0/XI0_23/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN0_8 XI11_0/net21_7_ xsel_23_ XI11_0/XI0/XI0_23/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN0_7 XI11_0/net21_8_ xsel_23_ XI11_0/XI0/XI0_23/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN0_6 XI11_0/net21_9_ xsel_23_ XI11_0/XI0/XI0_23/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN0_5 XI11_0/net21_10_ xsel_23_ XI11_0/XI0/XI0_23/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN0_4 XI11_0/net21_11_ xsel_23_ XI11_0/XI0/XI0_23/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN0_3 XI11_0/net21_12_ xsel_23_ XI11_0/XI0/XI0_23/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN0_2 XI11_0/net21_13_ xsel_23_ XI11_0/XI0/XI0_23/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN0_1 XI11_0/net21_14_ xsel_23_ XI11_0/XI0/XI0_23/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN0_0 XI11_0/net21_15_ xsel_23_ XI11_0/XI0/XI0_23/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN1_15 XI11_0/XI0/XI0_23/d__15_ xsel_23_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN1_14 XI11_0/XI0/XI0_23/d__14_ xsel_23_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN1_13 XI11_0/XI0/XI0_23/d__13_ xsel_23_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN1_12 XI11_0/XI0/XI0_23/d__12_ xsel_23_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN1_11 XI11_0/XI0/XI0_23/d__11_ xsel_23_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN1_10 XI11_0/XI0/XI0_23/d__10_ xsel_23_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN1_9 XI11_0/XI0/XI0_23/d__9_ xsel_23_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN1_8 XI11_0/XI0/XI0_23/d__8_ xsel_23_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN1_7 XI11_0/XI0/XI0_23/d__7_ xsel_23_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN1_6 XI11_0/XI0/XI0_23/d__6_ xsel_23_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN1_5 XI11_0/XI0/XI0_23/d__5_ xsel_23_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN1_4 XI11_0/XI0/XI0_23/d__4_ xsel_23_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN1_3 XI11_0/XI0/XI0_23/d__3_ xsel_23_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN1_2 XI11_0/XI0/XI0_23/d__2_ xsel_23_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN1_1 XI11_0/XI0/XI0_23/d__1_ xsel_23_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_23/MN1_0 XI11_0/XI0/XI0_23/d__0_ xsel_23_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN0_15 XI11_0/net21_0_ xsel_22_ XI11_0/XI0/XI0_22/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN0_14 XI11_0/net21_1_ xsel_22_ XI11_0/XI0/XI0_22/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN0_13 XI11_0/net21_2_ xsel_22_ XI11_0/XI0/XI0_22/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN0_12 XI11_0/net21_3_ xsel_22_ XI11_0/XI0/XI0_22/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN0_11 XI11_0/net21_4_ xsel_22_ XI11_0/XI0/XI0_22/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN0_10 XI11_0/net21_5_ xsel_22_ XI11_0/XI0/XI0_22/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN0_9 XI11_0/net21_6_ xsel_22_ XI11_0/XI0/XI0_22/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN0_8 XI11_0/net21_7_ xsel_22_ XI11_0/XI0/XI0_22/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN0_7 XI11_0/net21_8_ xsel_22_ XI11_0/XI0/XI0_22/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN0_6 XI11_0/net21_9_ xsel_22_ XI11_0/XI0/XI0_22/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN0_5 XI11_0/net21_10_ xsel_22_ XI11_0/XI0/XI0_22/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN0_4 XI11_0/net21_11_ xsel_22_ XI11_0/XI0/XI0_22/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN0_3 XI11_0/net21_12_ xsel_22_ XI11_0/XI0/XI0_22/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN0_2 XI11_0/net21_13_ xsel_22_ XI11_0/XI0/XI0_22/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN0_1 XI11_0/net21_14_ xsel_22_ XI11_0/XI0/XI0_22/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN0_0 XI11_0/net21_15_ xsel_22_ XI11_0/XI0/XI0_22/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN1_15 XI11_0/XI0/XI0_22/d__15_ xsel_22_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN1_14 XI11_0/XI0/XI0_22/d__14_ xsel_22_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN1_13 XI11_0/XI0/XI0_22/d__13_ xsel_22_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN1_12 XI11_0/XI0/XI0_22/d__12_ xsel_22_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN1_11 XI11_0/XI0/XI0_22/d__11_ xsel_22_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN1_10 XI11_0/XI0/XI0_22/d__10_ xsel_22_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN1_9 XI11_0/XI0/XI0_22/d__9_ xsel_22_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN1_8 XI11_0/XI0/XI0_22/d__8_ xsel_22_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN1_7 XI11_0/XI0/XI0_22/d__7_ xsel_22_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN1_6 XI11_0/XI0/XI0_22/d__6_ xsel_22_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN1_5 XI11_0/XI0/XI0_22/d__5_ xsel_22_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN1_4 XI11_0/XI0/XI0_22/d__4_ xsel_22_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN1_3 XI11_0/XI0/XI0_22/d__3_ xsel_22_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN1_2 XI11_0/XI0/XI0_22/d__2_ xsel_22_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN1_1 XI11_0/XI0/XI0_22/d__1_ xsel_22_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_22/MN1_0 XI11_0/XI0/XI0_22/d__0_ xsel_22_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN0_15 XI11_0/net21_0_ xsel_21_ XI11_0/XI0/XI0_21/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN0_14 XI11_0/net21_1_ xsel_21_ XI11_0/XI0/XI0_21/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN0_13 XI11_0/net21_2_ xsel_21_ XI11_0/XI0/XI0_21/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN0_12 XI11_0/net21_3_ xsel_21_ XI11_0/XI0/XI0_21/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN0_11 XI11_0/net21_4_ xsel_21_ XI11_0/XI0/XI0_21/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN0_10 XI11_0/net21_5_ xsel_21_ XI11_0/XI0/XI0_21/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN0_9 XI11_0/net21_6_ xsel_21_ XI11_0/XI0/XI0_21/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN0_8 XI11_0/net21_7_ xsel_21_ XI11_0/XI0/XI0_21/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN0_7 XI11_0/net21_8_ xsel_21_ XI11_0/XI0/XI0_21/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN0_6 XI11_0/net21_9_ xsel_21_ XI11_0/XI0/XI0_21/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN0_5 XI11_0/net21_10_ xsel_21_ XI11_0/XI0/XI0_21/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN0_4 XI11_0/net21_11_ xsel_21_ XI11_0/XI0/XI0_21/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN0_3 XI11_0/net21_12_ xsel_21_ XI11_0/XI0/XI0_21/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN0_2 XI11_0/net21_13_ xsel_21_ XI11_0/XI0/XI0_21/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN0_1 XI11_0/net21_14_ xsel_21_ XI11_0/XI0/XI0_21/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN0_0 XI11_0/net21_15_ xsel_21_ XI11_0/XI0/XI0_21/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN1_15 XI11_0/XI0/XI0_21/d__15_ xsel_21_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN1_14 XI11_0/XI0/XI0_21/d__14_ xsel_21_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN1_13 XI11_0/XI0/XI0_21/d__13_ xsel_21_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN1_12 XI11_0/XI0/XI0_21/d__12_ xsel_21_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN1_11 XI11_0/XI0/XI0_21/d__11_ xsel_21_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN1_10 XI11_0/XI0/XI0_21/d__10_ xsel_21_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN1_9 XI11_0/XI0/XI0_21/d__9_ xsel_21_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN1_8 XI11_0/XI0/XI0_21/d__8_ xsel_21_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN1_7 XI11_0/XI0/XI0_21/d__7_ xsel_21_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN1_6 XI11_0/XI0/XI0_21/d__6_ xsel_21_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN1_5 XI11_0/XI0/XI0_21/d__5_ xsel_21_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN1_4 XI11_0/XI0/XI0_21/d__4_ xsel_21_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN1_3 XI11_0/XI0/XI0_21/d__3_ xsel_21_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN1_2 XI11_0/XI0/XI0_21/d__2_ xsel_21_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN1_1 XI11_0/XI0/XI0_21/d__1_ xsel_21_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_21/MN1_0 XI11_0/XI0/XI0_21/d__0_ xsel_21_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN0_15 XI11_0/net21_0_ xsel_20_ XI11_0/XI0/XI0_20/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN0_14 XI11_0/net21_1_ xsel_20_ XI11_0/XI0/XI0_20/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN0_13 XI11_0/net21_2_ xsel_20_ XI11_0/XI0/XI0_20/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN0_12 XI11_0/net21_3_ xsel_20_ XI11_0/XI0/XI0_20/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN0_11 XI11_0/net21_4_ xsel_20_ XI11_0/XI0/XI0_20/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN0_10 XI11_0/net21_5_ xsel_20_ XI11_0/XI0/XI0_20/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN0_9 XI11_0/net21_6_ xsel_20_ XI11_0/XI0/XI0_20/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN0_8 XI11_0/net21_7_ xsel_20_ XI11_0/XI0/XI0_20/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN0_7 XI11_0/net21_8_ xsel_20_ XI11_0/XI0/XI0_20/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN0_6 XI11_0/net21_9_ xsel_20_ XI11_0/XI0/XI0_20/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN0_5 XI11_0/net21_10_ xsel_20_ XI11_0/XI0/XI0_20/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN0_4 XI11_0/net21_11_ xsel_20_ XI11_0/XI0/XI0_20/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN0_3 XI11_0/net21_12_ xsel_20_ XI11_0/XI0/XI0_20/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN0_2 XI11_0/net21_13_ xsel_20_ XI11_0/XI0/XI0_20/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN0_1 XI11_0/net21_14_ xsel_20_ XI11_0/XI0/XI0_20/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN0_0 XI11_0/net21_15_ xsel_20_ XI11_0/XI0/XI0_20/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN1_15 XI11_0/XI0/XI0_20/d__15_ xsel_20_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN1_14 XI11_0/XI0/XI0_20/d__14_ xsel_20_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN1_13 XI11_0/XI0/XI0_20/d__13_ xsel_20_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN1_12 XI11_0/XI0/XI0_20/d__12_ xsel_20_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN1_11 XI11_0/XI0/XI0_20/d__11_ xsel_20_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN1_10 XI11_0/XI0/XI0_20/d__10_ xsel_20_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN1_9 XI11_0/XI0/XI0_20/d__9_ xsel_20_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN1_8 XI11_0/XI0/XI0_20/d__8_ xsel_20_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN1_7 XI11_0/XI0/XI0_20/d__7_ xsel_20_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN1_6 XI11_0/XI0/XI0_20/d__6_ xsel_20_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN1_5 XI11_0/XI0/XI0_20/d__5_ xsel_20_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN1_4 XI11_0/XI0/XI0_20/d__4_ xsel_20_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN1_3 XI11_0/XI0/XI0_20/d__3_ xsel_20_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN1_2 XI11_0/XI0/XI0_20/d__2_ xsel_20_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN1_1 XI11_0/XI0/XI0_20/d__1_ xsel_20_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_20/MN1_0 XI11_0/XI0/XI0_20/d__0_ xsel_20_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN0_15 XI11_0/net21_0_ xsel_19_ XI11_0/XI0/XI0_19/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN0_14 XI11_0/net21_1_ xsel_19_ XI11_0/XI0/XI0_19/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN0_13 XI11_0/net21_2_ xsel_19_ XI11_0/XI0/XI0_19/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN0_12 XI11_0/net21_3_ xsel_19_ XI11_0/XI0/XI0_19/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN0_11 XI11_0/net21_4_ xsel_19_ XI11_0/XI0/XI0_19/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN0_10 XI11_0/net21_5_ xsel_19_ XI11_0/XI0/XI0_19/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN0_9 XI11_0/net21_6_ xsel_19_ XI11_0/XI0/XI0_19/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN0_8 XI11_0/net21_7_ xsel_19_ XI11_0/XI0/XI0_19/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN0_7 XI11_0/net21_8_ xsel_19_ XI11_0/XI0/XI0_19/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN0_6 XI11_0/net21_9_ xsel_19_ XI11_0/XI0/XI0_19/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN0_5 XI11_0/net21_10_ xsel_19_ XI11_0/XI0/XI0_19/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN0_4 XI11_0/net21_11_ xsel_19_ XI11_0/XI0/XI0_19/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN0_3 XI11_0/net21_12_ xsel_19_ XI11_0/XI0/XI0_19/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN0_2 XI11_0/net21_13_ xsel_19_ XI11_0/XI0/XI0_19/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN0_1 XI11_0/net21_14_ xsel_19_ XI11_0/XI0/XI0_19/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN0_0 XI11_0/net21_15_ xsel_19_ XI11_0/XI0/XI0_19/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN1_15 XI11_0/XI0/XI0_19/d__15_ xsel_19_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN1_14 XI11_0/XI0/XI0_19/d__14_ xsel_19_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN1_13 XI11_0/XI0/XI0_19/d__13_ xsel_19_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN1_12 XI11_0/XI0/XI0_19/d__12_ xsel_19_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN1_11 XI11_0/XI0/XI0_19/d__11_ xsel_19_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN1_10 XI11_0/XI0/XI0_19/d__10_ xsel_19_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN1_9 XI11_0/XI0/XI0_19/d__9_ xsel_19_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN1_8 XI11_0/XI0/XI0_19/d__8_ xsel_19_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN1_7 XI11_0/XI0/XI0_19/d__7_ xsel_19_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN1_6 XI11_0/XI0/XI0_19/d__6_ xsel_19_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN1_5 XI11_0/XI0/XI0_19/d__5_ xsel_19_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN1_4 XI11_0/XI0/XI0_19/d__4_ xsel_19_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN1_3 XI11_0/XI0/XI0_19/d__3_ xsel_19_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN1_2 XI11_0/XI0/XI0_19/d__2_ xsel_19_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN1_1 XI11_0/XI0/XI0_19/d__1_ xsel_19_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_19/MN1_0 XI11_0/XI0/XI0_19/d__0_ xsel_19_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN0_15 XI11_0/net21_0_ xsel_18_ XI11_0/XI0/XI0_18/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN0_14 XI11_0/net21_1_ xsel_18_ XI11_0/XI0/XI0_18/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN0_13 XI11_0/net21_2_ xsel_18_ XI11_0/XI0/XI0_18/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN0_12 XI11_0/net21_3_ xsel_18_ XI11_0/XI0/XI0_18/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN0_11 XI11_0/net21_4_ xsel_18_ XI11_0/XI0/XI0_18/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN0_10 XI11_0/net21_5_ xsel_18_ XI11_0/XI0/XI0_18/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN0_9 XI11_0/net21_6_ xsel_18_ XI11_0/XI0/XI0_18/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN0_8 XI11_0/net21_7_ xsel_18_ XI11_0/XI0/XI0_18/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN0_7 XI11_0/net21_8_ xsel_18_ XI11_0/XI0/XI0_18/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN0_6 XI11_0/net21_9_ xsel_18_ XI11_0/XI0/XI0_18/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN0_5 XI11_0/net21_10_ xsel_18_ XI11_0/XI0/XI0_18/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN0_4 XI11_0/net21_11_ xsel_18_ XI11_0/XI0/XI0_18/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN0_3 XI11_0/net21_12_ xsel_18_ XI11_0/XI0/XI0_18/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN0_2 XI11_0/net21_13_ xsel_18_ XI11_0/XI0/XI0_18/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN0_1 XI11_0/net21_14_ xsel_18_ XI11_0/XI0/XI0_18/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN0_0 XI11_0/net21_15_ xsel_18_ XI11_0/XI0/XI0_18/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN1_15 XI11_0/XI0/XI0_18/d__15_ xsel_18_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN1_14 XI11_0/XI0/XI0_18/d__14_ xsel_18_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN1_13 XI11_0/XI0/XI0_18/d__13_ xsel_18_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN1_12 XI11_0/XI0/XI0_18/d__12_ xsel_18_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN1_11 XI11_0/XI0/XI0_18/d__11_ xsel_18_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN1_10 XI11_0/XI0/XI0_18/d__10_ xsel_18_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN1_9 XI11_0/XI0/XI0_18/d__9_ xsel_18_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN1_8 XI11_0/XI0/XI0_18/d__8_ xsel_18_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN1_7 XI11_0/XI0/XI0_18/d__7_ xsel_18_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN1_6 XI11_0/XI0/XI0_18/d__6_ xsel_18_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN1_5 XI11_0/XI0/XI0_18/d__5_ xsel_18_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN1_4 XI11_0/XI0/XI0_18/d__4_ xsel_18_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN1_3 XI11_0/XI0/XI0_18/d__3_ xsel_18_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN1_2 XI11_0/XI0/XI0_18/d__2_ xsel_18_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN1_1 XI11_0/XI0/XI0_18/d__1_ xsel_18_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_18/MN1_0 XI11_0/XI0/XI0_18/d__0_ xsel_18_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN0_15 XI11_0/net21_0_ xsel_17_ XI11_0/XI0/XI0_17/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN0_14 XI11_0/net21_1_ xsel_17_ XI11_0/XI0/XI0_17/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN0_13 XI11_0/net21_2_ xsel_17_ XI11_0/XI0/XI0_17/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN0_12 XI11_0/net21_3_ xsel_17_ XI11_0/XI0/XI0_17/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN0_11 XI11_0/net21_4_ xsel_17_ XI11_0/XI0/XI0_17/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN0_10 XI11_0/net21_5_ xsel_17_ XI11_0/XI0/XI0_17/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN0_9 XI11_0/net21_6_ xsel_17_ XI11_0/XI0/XI0_17/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN0_8 XI11_0/net21_7_ xsel_17_ XI11_0/XI0/XI0_17/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN0_7 XI11_0/net21_8_ xsel_17_ XI11_0/XI0/XI0_17/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN0_6 XI11_0/net21_9_ xsel_17_ XI11_0/XI0/XI0_17/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN0_5 XI11_0/net21_10_ xsel_17_ XI11_0/XI0/XI0_17/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN0_4 XI11_0/net21_11_ xsel_17_ XI11_0/XI0/XI0_17/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN0_3 XI11_0/net21_12_ xsel_17_ XI11_0/XI0/XI0_17/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN0_2 XI11_0/net21_13_ xsel_17_ XI11_0/XI0/XI0_17/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN0_1 XI11_0/net21_14_ xsel_17_ XI11_0/XI0/XI0_17/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN0_0 XI11_0/net21_15_ xsel_17_ XI11_0/XI0/XI0_17/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN1_15 XI11_0/XI0/XI0_17/d__15_ xsel_17_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN1_14 XI11_0/XI0/XI0_17/d__14_ xsel_17_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN1_13 XI11_0/XI0/XI0_17/d__13_ xsel_17_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN1_12 XI11_0/XI0/XI0_17/d__12_ xsel_17_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN1_11 XI11_0/XI0/XI0_17/d__11_ xsel_17_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN1_10 XI11_0/XI0/XI0_17/d__10_ xsel_17_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN1_9 XI11_0/XI0/XI0_17/d__9_ xsel_17_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN1_8 XI11_0/XI0/XI0_17/d__8_ xsel_17_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN1_7 XI11_0/XI0/XI0_17/d__7_ xsel_17_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN1_6 XI11_0/XI0/XI0_17/d__6_ xsel_17_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN1_5 XI11_0/XI0/XI0_17/d__5_ xsel_17_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN1_4 XI11_0/XI0/XI0_17/d__4_ xsel_17_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN1_3 XI11_0/XI0/XI0_17/d__3_ xsel_17_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN1_2 XI11_0/XI0/XI0_17/d__2_ xsel_17_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN1_1 XI11_0/XI0/XI0_17/d__1_ xsel_17_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_17/MN1_0 XI11_0/XI0/XI0_17/d__0_ xsel_17_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN0_15 XI11_0/net21_0_ xsel_16_ XI11_0/XI0/XI0_16/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN0_14 XI11_0/net21_1_ xsel_16_ XI11_0/XI0/XI0_16/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN0_13 XI11_0/net21_2_ xsel_16_ XI11_0/XI0/XI0_16/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN0_12 XI11_0/net21_3_ xsel_16_ XI11_0/XI0/XI0_16/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN0_11 XI11_0/net21_4_ xsel_16_ XI11_0/XI0/XI0_16/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN0_10 XI11_0/net21_5_ xsel_16_ XI11_0/XI0/XI0_16/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN0_9 XI11_0/net21_6_ xsel_16_ XI11_0/XI0/XI0_16/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN0_8 XI11_0/net21_7_ xsel_16_ XI11_0/XI0/XI0_16/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN0_7 XI11_0/net21_8_ xsel_16_ XI11_0/XI0/XI0_16/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN0_6 XI11_0/net21_9_ xsel_16_ XI11_0/XI0/XI0_16/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN0_5 XI11_0/net21_10_ xsel_16_ XI11_0/XI0/XI0_16/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN0_4 XI11_0/net21_11_ xsel_16_ XI11_0/XI0/XI0_16/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN0_3 XI11_0/net21_12_ xsel_16_ XI11_0/XI0/XI0_16/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN0_2 XI11_0/net21_13_ xsel_16_ XI11_0/XI0/XI0_16/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN0_1 XI11_0/net21_14_ xsel_16_ XI11_0/XI0/XI0_16/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN0_0 XI11_0/net21_15_ xsel_16_ XI11_0/XI0/XI0_16/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN1_15 XI11_0/XI0/XI0_16/d__15_ xsel_16_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN1_14 XI11_0/XI0/XI0_16/d__14_ xsel_16_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN1_13 XI11_0/XI0/XI0_16/d__13_ xsel_16_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN1_12 XI11_0/XI0/XI0_16/d__12_ xsel_16_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN1_11 XI11_0/XI0/XI0_16/d__11_ xsel_16_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN1_10 XI11_0/XI0/XI0_16/d__10_ xsel_16_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN1_9 XI11_0/XI0/XI0_16/d__9_ xsel_16_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN1_8 XI11_0/XI0/XI0_16/d__8_ xsel_16_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN1_7 XI11_0/XI0/XI0_16/d__7_ xsel_16_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN1_6 XI11_0/XI0/XI0_16/d__6_ xsel_16_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN1_5 XI11_0/XI0/XI0_16/d__5_ xsel_16_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN1_4 XI11_0/XI0/XI0_16/d__4_ xsel_16_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN1_3 XI11_0/XI0/XI0_16/d__3_ xsel_16_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN1_2 XI11_0/XI0/XI0_16/d__2_ xsel_16_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN1_1 XI11_0/XI0/XI0_16/d__1_ xsel_16_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_16/MN1_0 XI11_0/XI0/XI0_16/d__0_ xsel_16_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN0_15 XI11_0/net21_0_ xsel_15_ XI11_0/XI0/XI0_15/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN0_14 XI11_0/net21_1_ xsel_15_ XI11_0/XI0/XI0_15/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN0_13 XI11_0/net21_2_ xsel_15_ XI11_0/XI0/XI0_15/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN0_12 XI11_0/net21_3_ xsel_15_ XI11_0/XI0/XI0_15/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN0_11 XI11_0/net21_4_ xsel_15_ XI11_0/XI0/XI0_15/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN0_10 XI11_0/net21_5_ xsel_15_ XI11_0/XI0/XI0_15/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN0_9 XI11_0/net21_6_ xsel_15_ XI11_0/XI0/XI0_15/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN0_8 XI11_0/net21_7_ xsel_15_ XI11_0/XI0/XI0_15/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN0_7 XI11_0/net21_8_ xsel_15_ XI11_0/XI0/XI0_15/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN0_6 XI11_0/net21_9_ xsel_15_ XI11_0/XI0/XI0_15/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN0_5 XI11_0/net21_10_ xsel_15_ XI11_0/XI0/XI0_15/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN0_4 XI11_0/net21_11_ xsel_15_ XI11_0/XI0/XI0_15/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN0_3 XI11_0/net21_12_ xsel_15_ XI11_0/XI0/XI0_15/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN0_2 XI11_0/net21_13_ xsel_15_ XI11_0/XI0/XI0_15/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN0_1 XI11_0/net21_14_ xsel_15_ XI11_0/XI0/XI0_15/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN0_0 XI11_0/net21_15_ xsel_15_ XI11_0/XI0/XI0_15/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN1_15 XI11_0/XI0/XI0_15/d__15_ xsel_15_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN1_14 XI11_0/XI0/XI0_15/d__14_ xsel_15_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN1_13 XI11_0/XI0/XI0_15/d__13_ xsel_15_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN1_12 XI11_0/XI0/XI0_15/d__12_ xsel_15_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN1_11 XI11_0/XI0/XI0_15/d__11_ xsel_15_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN1_10 XI11_0/XI0/XI0_15/d__10_ xsel_15_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN1_9 XI11_0/XI0/XI0_15/d__9_ xsel_15_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN1_8 XI11_0/XI0/XI0_15/d__8_ xsel_15_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN1_7 XI11_0/XI0/XI0_15/d__7_ xsel_15_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN1_6 XI11_0/XI0/XI0_15/d__6_ xsel_15_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN1_5 XI11_0/XI0/XI0_15/d__5_ xsel_15_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN1_4 XI11_0/XI0/XI0_15/d__4_ xsel_15_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN1_3 XI11_0/XI0/XI0_15/d__3_ xsel_15_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN1_2 XI11_0/XI0/XI0_15/d__2_ xsel_15_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN1_1 XI11_0/XI0/XI0_15/d__1_ xsel_15_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_15/MN1_0 XI11_0/XI0/XI0_15/d__0_ xsel_15_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN0_15 XI11_0/net21_0_ xsel_14_ XI11_0/XI0/XI0_14/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN0_14 XI11_0/net21_1_ xsel_14_ XI11_0/XI0/XI0_14/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN0_13 XI11_0/net21_2_ xsel_14_ XI11_0/XI0/XI0_14/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN0_12 XI11_0/net21_3_ xsel_14_ XI11_0/XI0/XI0_14/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN0_11 XI11_0/net21_4_ xsel_14_ XI11_0/XI0/XI0_14/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN0_10 XI11_0/net21_5_ xsel_14_ XI11_0/XI0/XI0_14/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN0_9 XI11_0/net21_6_ xsel_14_ XI11_0/XI0/XI0_14/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN0_8 XI11_0/net21_7_ xsel_14_ XI11_0/XI0/XI0_14/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN0_7 XI11_0/net21_8_ xsel_14_ XI11_0/XI0/XI0_14/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN0_6 XI11_0/net21_9_ xsel_14_ XI11_0/XI0/XI0_14/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN0_5 XI11_0/net21_10_ xsel_14_ XI11_0/XI0/XI0_14/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN0_4 XI11_0/net21_11_ xsel_14_ XI11_0/XI0/XI0_14/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN0_3 XI11_0/net21_12_ xsel_14_ XI11_0/XI0/XI0_14/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN0_2 XI11_0/net21_13_ xsel_14_ XI11_0/XI0/XI0_14/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN0_1 XI11_0/net21_14_ xsel_14_ XI11_0/XI0/XI0_14/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN0_0 XI11_0/net21_15_ xsel_14_ XI11_0/XI0/XI0_14/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN1_15 XI11_0/XI0/XI0_14/d__15_ xsel_14_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN1_14 XI11_0/XI0/XI0_14/d__14_ xsel_14_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN1_13 XI11_0/XI0/XI0_14/d__13_ xsel_14_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN1_12 XI11_0/XI0/XI0_14/d__12_ xsel_14_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN1_11 XI11_0/XI0/XI0_14/d__11_ xsel_14_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN1_10 XI11_0/XI0/XI0_14/d__10_ xsel_14_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN1_9 XI11_0/XI0/XI0_14/d__9_ xsel_14_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN1_8 XI11_0/XI0/XI0_14/d__8_ xsel_14_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN1_7 XI11_0/XI0/XI0_14/d__7_ xsel_14_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN1_6 XI11_0/XI0/XI0_14/d__6_ xsel_14_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN1_5 XI11_0/XI0/XI0_14/d__5_ xsel_14_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN1_4 XI11_0/XI0/XI0_14/d__4_ xsel_14_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN1_3 XI11_0/XI0/XI0_14/d__3_ xsel_14_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN1_2 XI11_0/XI0/XI0_14/d__2_ xsel_14_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN1_1 XI11_0/XI0/XI0_14/d__1_ xsel_14_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_14/MN1_0 XI11_0/XI0/XI0_14/d__0_ xsel_14_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN0_15 XI11_0/net21_0_ xsel_13_ XI11_0/XI0/XI0_13/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN0_14 XI11_0/net21_1_ xsel_13_ XI11_0/XI0/XI0_13/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN0_13 XI11_0/net21_2_ xsel_13_ XI11_0/XI0/XI0_13/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN0_12 XI11_0/net21_3_ xsel_13_ XI11_0/XI0/XI0_13/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN0_11 XI11_0/net21_4_ xsel_13_ XI11_0/XI0/XI0_13/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN0_10 XI11_0/net21_5_ xsel_13_ XI11_0/XI0/XI0_13/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN0_9 XI11_0/net21_6_ xsel_13_ XI11_0/XI0/XI0_13/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN0_8 XI11_0/net21_7_ xsel_13_ XI11_0/XI0/XI0_13/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN0_7 XI11_0/net21_8_ xsel_13_ XI11_0/XI0/XI0_13/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN0_6 XI11_0/net21_9_ xsel_13_ XI11_0/XI0/XI0_13/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN0_5 XI11_0/net21_10_ xsel_13_ XI11_0/XI0/XI0_13/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN0_4 XI11_0/net21_11_ xsel_13_ XI11_0/XI0/XI0_13/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN0_3 XI11_0/net21_12_ xsel_13_ XI11_0/XI0/XI0_13/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN0_2 XI11_0/net21_13_ xsel_13_ XI11_0/XI0/XI0_13/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN0_1 XI11_0/net21_14_ xsel_13_ XI11_0/XI0/XI0_13/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN0_0 XI11_0/net21_15_ xsel_13_ XI11_0/XI0/XI0_13/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN1_15 XI11_0/XI0/XI0_13/d__15_ xsel_13_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN1_14 XI11_0/XI0/XI0_13/d__14_ xsel_13_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN1_13 XI11_0/XI0/XI0_13/d__13_ xsel_13_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN1_12 XI11_0/XI0/XI0_13/d__12_ xsel_13_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN1_11 XI11_0/XI0/XI0_13/d__11_ xsel_13_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN1_10 XI11_0/XI0/XI0_13/d__10_ xsel_13_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN1_9 XI11_0/XI0/XI0_13/d__9_ xsel_13_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN1_8 XI11_0/XI0/XI0_13/d__8_ xsel_13_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN1_7 XI11_0/XI0/XI0_13/d__7_ xsel_13_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN1_6 XI11_0/XI0/XI0_13/d__6_ xsel_13_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN1_5 XI11_0/XI0/XI0_13/d__5_ xsel_13_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN1_4 XI11_0/XI0/XI0_13/d__4_ xsel_13_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN1_3 XI11_0/XI0/XI0_13/d__3_ xsel_13_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN1_2 XI11_0/XI0/XI0_13/d__2_ xsel_13_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN1_1 XI11_0/XI0/XI0_13/d__1_ xsel_13_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_13/MN1_0 XI11_0/XI0/XI0_13/d__0_ xsel_13_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN0_15 XI11_0/net21_0_ xsel_12_ XI11_0/XI0/XI0_12/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN0_14 XI11_0/net21_1_ xsel_12_ XI11_0/XI0/XI0_12/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN0_13 XI11_0/net21_2_ xsel_12_ XI11_0/XI0/XI0_12/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN0_12 XI11_0/net21_3_ xsel_12_ XI11_0/XI0/XI0_12/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN0_11 XI11_0/net21_4_ xsel_12_ XI11_0/XI0/XI0_12/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN0_10 XI11_0/net21_5_ xsel_12_ XI11_0/XI0/XI0_12/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN0_9 XI11_0/net21_6_ xsel_12_ XI11_0/XI0/XI0_12/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN0_8 XI11_0/net21_7_ xsel_12_ XI11_0/XI0/XI0_12/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN0_7 XI11_0/net21_8_ xsel_12_ XI11_0/XI0/XI0_12/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN0_6 XI11_0/net21_9_ xsel_12_ XI11_0/XI0/XI0_12/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN0_5 XI11_0/net21_10_ xsel_12_ XI11_0/XI0/XI0_12/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN0_4 XI11_0/net21_11_ xsel_12_ XI11_0/XI0/XI0_12/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN0_3 XI11_0/net21_12_ xsel_12_ XI11_0/XI0/XI0_12/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN0_2 XI11_0/net21_13_ xsel_12_ XI11_0/XI0/XI0_12/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN0_1 XI11_0/net21_14_ xsel_12_ XI11_0/XI0/XI0_12/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN0_0 XI11_0/net21_15_ xsel_12_ XI11_0/XI0/XI0_12/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN1_15 XI11_0/XI0/XI0_12/d__15_ xsel_12_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN1_14 XI11_0/XI0/XI0_12/d__14_ xsel_12_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN1_13 XI11_0/XI0/XI0_12/d__13_ xsel_12_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN1_12 XI11_0/XI0/XI0_12/d__12_ xsel_12_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN1_11 XI11_0/XI0/XI0_12/d__11_ xsel_12_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN1_10 XI11_0/XI0/XI0_12/d__10_ xsel_12_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN1_9 XI11_0/XI0/XI0_12/d__9_ xsel_12_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN1_8 XI11_0/XI0/XI0_12/d__8_ xsel_12_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN1_7 XI11_0/XI0/XI0_12/d__7_ xsel_12_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN1_6 XI11_0/XI0/XI0_12/d__6_ xsel_12_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN1_5 XI11_0/XI0/XI0_12/d__5_ xsel_12_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN1_4 XI11_0/XI0/XI0_12/d__4_ xsel_12_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN1_3 XI11_0/XI0/XI0_12/d__3_ xsel_12_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN1_2 XI11_0/XI0/XI0_12/d__2_ xsel_12_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN1_1 XI11_0/XI0/XI0_12/d__1_ xsel_12_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_12/MN1_0 XI11_0/XI0/XI0_12/d__0_ xsel_12_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN0_15 XI11_0/net21_0_ xsel_11_ XI11_0/XI0/XI0_11/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN0_14 XI11_0/net21_1_ xsel_11_ XI11_0/XI0/XI0_11/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN0_13 XI11_0/net21_2_ xsel_11_ XI11_0/XI0/XI0_11/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN0_12 XI11_0/net21_3_ xsel_11_ XI11_0/XI0/XI0_11/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN0_11 XI11_0/net21_4_ xsel_11_ XI11_0/XI0/XI0_11/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN0_10 XI11_0/net21_5_ xsel_11_ XI11_0/XI0/XI0_11/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN0_9 XI11_0/net21_6_ xsel_11_ XI11_0/XI0/XI0_11/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN0_8 XI11_0/net21_7_ xsel_11_ XI11_0/XI0/XI0_11/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN0_7 XI11_0/net21_8_ xsel_11_ XI11_0/XI0/XI0_11/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN0_6 XI11_0/net21_9_ xsel_11_ XI11_0/XI0/XI0_11/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN0_5 XI11_0/net21_10_ xsel_11_ XI11_0/XI0/XI0_11/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN0_4 XI11_0/net21_11_ xsel_11_ XI11_0/XI0/XI0_11/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN0_3 XI11_0/net21_12_ xsel_11_ XI11_0/XI0/XI0_11/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN0_2 XI11_0/net21_13_ xsel_11_ XI11_0/XI0/XI0_11/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN0_1 XI11_0/net21_14_ xsel_11_ XI11_0/XI0/XI0_11/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN0_0 XI11_0/net21_15_ xsel_11_ XI11_0/XI0/XI0_11/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN1_15 XI11_0/XI0/XI0_11/d__15_ xsel_11_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN1_14 XI11_0/XI0/XI0_11/d__14_ xsel_11_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN1_13 XI11_0/XI0/XI0_11/d__13_ xsel_11_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN1_12 XI11_0/XI0/XI0_11/d__12_ xsel_11_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN1_11 XI11_0/XI0/XI0_11/d__11_ xsel_11_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN1_10 XI11_0/XI0/XI0_11/d__10_ xsel_11_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN1_9 XI11_0/XI0/XI0_11/d__9_ xsel_11_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN1_8 XI11_0/XI0/XI0_11/d__8_ xsel_11_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN1_7 XI11_0/XI0/XI0_11/d__7_ xsel_11_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN1_6 XI11_0/XI0/XI0_11/d__6_ xsel_11_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN1_5 XI11_0/XI0/XI0_11/d__5_ xsel_11_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN1_4 XI11_0/XI0/XI0_11/d__4_ xsel_11_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN1_3 XI11_0/XI0/XI0_11/d__3_ xsel_11_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN1_2 XI11_0/XI0/XI0_11/d__2_ xsel_11_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN1_1 XI11_0/XI0/XI0_11/d__1_ xsel_11_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_11/MN1_0 XI11_0/XI0/XI0_11/d__0_ xsel_11_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN0_15 XI11_0/net21_0_ xsel_10_ XI11_0/XI0/XI0_10/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN0_14 XI11_0/net21_1_ xsel_10_ XI11_0/XI0/XI0_10/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN0_13 XI11_0/net21_2_ xsel_10_ XI11_0/XI0/XI0_10/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN0_12 XI11_0/net21_3_ xsel_10_ XI11_0/XI0/XI0_10/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN0_11 XI11_0/net21_4_ xsel_10_ XI11_0/XI0/XI0_10/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN0_10 XI11_0/net21_5_ xsel_10_ XI11_0/XI0/XI0_10/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN0_9 XI11_0/net21_6_ xsel_10_ XI11_0/XI0/XI0_10/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN0_8 XI11_0/net21_7_ xsel_10_ XI11_0/XI0/XI0_10/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN0_7 XI11_0/net21_8_ xsel_10_ XI11_0/XI0/XI0_10/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN0_6 XI11_0/net21_9_ xsel_10_ XI11_0/XI0/XI0_10/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN0_5 XI11_0/net21_10_ xsel_10_ XI11_0/XI0/XI0_10/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN0_4 XI11_0/net21_11_ xsel_10_ XI11_0/XI0/XI0_10/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN0_3 XI11_0/net21_12_ xsel_10_ XI11_0/XI0/XI0_10/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN0_2 XI11_0/net21_13_ xsel_10_ XI11_0/XI0/XI0_10/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN0_1 XI11_0/net21_14_ xsel_10_ XI11_0/XI0/XI0_10/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN0_0 XI11_0/net21_15_ xsel_10_ XI11_0/XI0/XI0_10/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN1_15 XI11_0/XI0/XI0_10/d__15_ xsel_10_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN1_14 XI11_0/XI0/XI0_10/d__14_ xsel_10_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN1_13 XI11_0/XI0/XI0_10/d__13_ xsel_10_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN1_12 XI11_0/XI0/XI0_10/d__12_ xsel_10_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN1_11 XI11_0/XI0/XI0_10/d__11_ xsel_10_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN1_10 XI11_0/XI0/XI0_10/d__10_ xsel_10_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN1_9 XI11_0/XI0/XI0_10/d__9_ xsel_10_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN1_8 XI11_0/XI0/XI0_10/d__8_ xsel_10_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN1_7 XI11_0/XI0/XI0_10/d__7_ xsel_10_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN1_6 XI11_0/XI0/XI0_10/d__6_ xsel_10_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN1_5 XI11_0/XI0/XI0_10/d__5_ xsel_10_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN1_4 XI11_0/XI0/XI0_10/d__4_ xsel_10_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN1_3 XI11_0/XI0/XI0_10/d__3_ xsel_10_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN1_2 XI11_0/XI0/XI0_10/d__2_ xsel_10_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN1_1 XI11_0/XI0/XI0_10/d__1_ xsel_10_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_10/MN1_0 XI11_0/XI0/XI0_10/d__0_ xsel_10_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN0_15 XI11_0/net21_0_ xsel_9_ XI11_0/XI0/XI0_9/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN0_14 XI11_0/net21_1_ xsel_9_ XI11_0/XI0/XI0_9/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN0_13 XI11_0/net21_2_ xsel_9_ XI11_0/XI0/XI0_9/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN0_12 XI11_0/net21_3_ xsel_9_ XI11_0/XI0/XI0_9/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN0_11 XI11_0/net21_4_ xsel_9_ XI11_0/XI0/XI0_9/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN0_10 XI11_0/net21_5_ xsel_9_ XI11_0/XI0/XI0_9/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN0_9 XI11_0/net21_6_ xsel_9_ XI11_0/XI0/XI0_9/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN0_8 XI11_0/net21_7_ xsel_9_ XI11_0/XI0/XI0_9/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN0_7 XI11_0/net21_8_ xsel_9_ XI11_0/XI0/XI0_9/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN0_6 XI11_0/net21_9_ xsel_9_ XI11_0/XI0/XI0_9/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN0_5 XI11_0/net21_10_ xsel_9_ XI11_0/XI0/XI0_9/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN0_4 XI11_0/net21_11_ xsel_9_ XI11_0/XI0/XI0_9/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN0_3 XI11_0/net21_12_ xsel_9_ XI11_0/XI0/XI0_9/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN0_2 XI11_0/net21_13_ xsel_9_ XI11_0/XI0/XI0_9/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN0_1 XI11_0/net21_14_ xsel_9_ XI11_0/XI0/XI0_9/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN0_0 XI11_0/net21_15_ xsel_9_ XI11_0/XI0/XI0_9/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN1_15 XI11_0/XI0/XI0_9/d__15_ xsel_9_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN1_14 XI11_0/XI0/XI0_9/d__14_ xsel_9_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN1_13 XI11_0/XI0/XI0_9/d__13_ xsel_9_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN1_12 XI11_0/XI0/XI0_9/d__12_ xsel_9_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN1_11 XI11_0/XI0/XI0_9/d__11_ xsel_9_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN1_10 XI11_0/XI0/XI0_9/d__10_ xsel_9_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN1_9 XI11_0/XI0/XI0_9/d__9_ xsel_9_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN1_8 XI11_0/XI0/XI0_9/d__8_ xsel_9_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN1_7 XI11_0/XI0/XI0_9/d__7_ xsel_9_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN1_6 XI11_0/XI0/XI0_9/d__6_ xsel_9_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN1_5 XI11_0/XI0/XI0_9/d__5_ xsel_9_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN1_4 XI11_0/XI0/XI0_9/d__4_ xsel_9_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN1_3 XI11_0/XI0/XI0_9/d__3_ xsel_9_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN1_2 XI11_0/XI0/XI0_9/d__2_ xsel_9_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN1_1 XI11_0/XI0/XI0_9/d__1_ xsel_9_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_9/MN1_0 XI11_0/XI0/XI0_9/d__0_ xsel_9_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN0_15 XI11_0/net21_0_ xsel_8_ XI11_0/XI0/XI0_8/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN0_14 XI11_0/net21_1_ xsel_8_ XI11_0/XI0/XI0_8/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN0_13 XI11_0/net21_2_ xsel_8_ XI11_0/XI0/XI0_8/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN0_12 XI11_0/net21_3_ xsel_8_ XI11_0/XI0/XI0_8/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN0_11 XI11_0/net21_4_ xsel_8_ XI11_0/XI0/XI0_8/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN0_10 XI11_0/net21_5_ xsel_8_ XI11_0/XI0/XI0_8/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN0_9 XI11_0/net21_6_ xsel_8_ XI11_0/XI0/XI0_8/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN0_8 XI11_0/net21_7_ xsel_8_ XI11_0/XI0/XI0_8/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN0_7 XI11_0/net21_8_ xsel_8_ XI11_0/XI0/XI0_8/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN0_6 XI11_0/net21_9_ xsel_8_ XI11_0/XI0/XI0_8/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN0_5 XI11_0/net21_10_ xsel_8_ XI11_0/XI0/XI0_8/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN0_4 XI11_0/net21_11_ xsel_8_ XI11_0/XI0/XI0_8/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN0_3 XI11_0/net21_12_ xsel_8_ XI11_0/XI0/XI0_8/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN0_2 XI11_0/net21_13_ xsel_8_ XI11_0/XI0/XI0_8/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN0_1 XI11_0/net21_14_ xsel_8_ XI11_0/XI0/XI0_8/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN0_0 XI11_0/net21_15_ xsel_8_ XI11_0/XI0/XI0_8/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN1_15 XI11_0/XI0/XI0_8/d__15_ xsel_8_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN1_14 XI11_0/XI0/XI0_8/d__14_ xsel_8_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN1_13 XI11_0/XI0/XI0_8/d__13_ xsel_8_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN1_12 XI11_0/XI0/XI0_8/d__12_ xsel_8_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN1_11 XI11_0/XI0/XI0_8/d__11_ xsel_8_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN1_10 XI11_0/XI0/XI0_8/d__10_ xsel_8_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN1_9 XI11_0/XI0/XI0_8/d__9_ xsel_8_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN1_8 XI11_0/XI0/XI0_8/d__8_ xsel_8_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN1_7 XI11_0/XI0/XI0_8/d__7_ xsel_8_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN1_6 XI11_0/XI0/XI0_8/d__6_ xsel_8_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN1_5 XI11_0/XI0/XI0_8/d__5_ xsel_8_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN1_4 XI11_0/XI0/XI0_8/d__4_ xsel_8_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN1_3 XI11_0/XI0/XI0_8/d__3_ xsel_8_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN1_2 XI11_0/XI0/XI0_8/d__2_ xsel_8_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN1_1 XI11_0/XI0/XI0_8/d__1_ xsel_8_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_8/MN1_0 XI11_0/XI0/XI0_8/d__0_ xsel_8_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN0_15 XI11_0/net21_0_ xsel_7_ XI11_0/XI0/XI0_7/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN0_14 XI11_0/net21_1_ xsel_7_ XI11_0/XI0/XI0_7/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN0_13 XI11_0/net21_2_ xsel_7_ XI11_0/XI0/XI0_7/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN0_12 XI11_0/net21_3_ xsel_7_ XI11_0/XI0/XI0_7/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN0_11 XI11_0/net21_4_ xsel_7_ XI11_0/XI0/XI0_7/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN0_10 XI11_0/net21_5_ xsel_7_ XI11_0/XI0/XI0_7/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN0_9 XI11_0/net21_6_ xsel_7_ XI11_0/XI0/XI0_7/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN0_8 XI11_0/net21_7_ xsel_7_ XI11_0/XI0/XI0_7/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN0_7 XI11_0/net21_8_ xsel_7_ XI11_0/XI0/XI0_7/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN0_6 XI11_0/net21_9_ xsel_7_ XI11_0/XI0/XI0_7/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN0_5 XI11_0/net21_10_ xsel_7_ XI11_0/XI0/XI0_7/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN0_4 XI11_0/net21_11_ xsel_7_ XI11_0/XI0/XI0_7/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN0_3 XI11_0/net21_12_ xsel_7_ XI11_0/XI0/XI0_7/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN0_2 XI11_0/net21_13_ xsel_7_ XI11_0/XI0/XI0_7/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN0_1 XI11_0/net21_14_ xsel_7_ XI11_0/XI0/XI0_7/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN0_0 XI11_0/net21_15_ xsel_7_ XI11_0/XI0/XI0_7/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN1_15 XI11_0/XI0/XI0_7/d__15_ xsel_7_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN1_14 XI11_0/XI0/XI0_7/d__14_ xsel_7_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN1_13 XI11_0/XI0/XI0_7/d__13_ xsel_7_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN1_12 XI11_0/XI0/XI0_7/d__12_ xsel_7_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN1_11 XI11_0/XI0/XI0_7/d__11_ xsel_7_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN1_10 XI11_0/XI0/XI0_7/d__10_ xsel_7_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN1_9 XI11_0/XI0/XI0_7/d__9_ xsel_7_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN1_8 XI11_0/XI0/XI0_7/d__8_ xsel_7_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN1_7 XI11_0/XI0/XI0_7/d__7_ xsel_7_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN1_6 XI11_0/XI0/XI0_7/d__6_ xsel_7_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN1_5 XI11_0/XI0/XI0_7/d__5_ xsel_7_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN1_4 XI11_0/XI0/XI0_7/d__4_ xsel_7_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN1_3 XI11_0/XI0/XI0_7/d__3_ xsel_7_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN1_2 XI11_0/XI0/XI0_7/d__2_ xsel_7_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN1_1 XI11_0/XI0/XI0_7/d__1_ xsel_7_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_7/MN1_0 XI11_0/XI0/XI0_7/d__0_ xsel_7_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN0_15 XI11_0/net21_0_ xsel_6_ XI11_0/XI0/XI0_6/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN0_14 XI11_0/net21_1_ xsel_6_ XI11_0/XI0/XI0_6/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN0_13 XI11_0/net21_2_ xsel_6_ XI11_0/XI0/XI0_6/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN0_12 XI11_0/net21_3_ xsel_6_ XI11_0/XI0/XI0_6/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN0_11 XI11_0/net21_4_ xsel_6_ XI11_0/XI0/XI0_6/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN0_10 XI11_0/net21_5_ xsel_6_ XI11_0/XI0/XI0_6/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN0_9 XI11_0/net21_6_ xsel_6_ XI11_0/XI0/XI0_6/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN0_8 XI11_0/net21_7_ xsel_6_ XI11_0/XI0/XI0_6/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN0_7 XI11_0/net21_8_ xsel_6_ XI11_0/XI0/XI0_6/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN0_6 XI11_0/net21_9_ xsel_6_ XI11_0/XI0/XI0_6/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN0_5 XI11_0/net21_10_ xsel_6_ XI11_0/XI0/XI0_6/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN0_4 XI11_0/net21_11_ xsel_6_ XI11_0/XI0/XI0_6/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN0_3 XI11_0/net21_12_ xsel_6_ XI11_0/XI0/XI0_6/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN0_2 XI11_0/net21_13_ xsel_6_ XI11_0/XI0/XI0_6/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN0_1 XI11_0/net21_14_ xsel_6_ XI11_0/XI0/XI0_6/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN0_0 XI11_0/net21_15_ xsel_6_ XI11_0/XI0/XI0_6/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN1_15 XI11_0/XI0/XI0_6/d__15_ xsel_6_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN1_14 XI11_0/XI0/XI0_6/d__14_ xsel_6_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN1_13 XI11_0/XI0/XI0_6/d__13_ xsel_6_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN1_12 XI11_0/XI0/XI0_6/d__12_ xsel_6_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN1_11 XI11_0/XI0/XI0_6/d__11_ xsel_6_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN1_10 XI11_0/XI0/XI0_6/d__10_ xsel_6_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN1_9 XI11_0/XI0/XI0_6/d__9_ xsel_6_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN1_8 XI11_0/XI0/XI0_6/d__8_ xsel_6_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN1_7 XI11_0/XI0/XI0_6/d__7_ xsel_6_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN1_6 XI11_0/XI0/XI0_6/d__6_ xsel_6_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN1_5 XI11_0/XI0/XI0_6/d__5_ xsel_6_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN1_4 XI11_0/XI0/XI0_6/d__4_ xsel_6_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN1_3 XI11_0/XI0/XI0_6/d__3_ xsel_6_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN1_2 XI11_0/XI0/XI0_6/d__2_ xsel_6_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN1_1 XI11_0/XI0/XI0_6/d__1_ xsel_6_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_6/MN1_0 XI11_0/XI0/XI0_6/d__0_ xsel_6_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN0_15 XI11_0/net21_0_ xsel_5_ XI11_0/XI0/XI0_5/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN0_14 XI11_0/net21_1_ xsel_5_ XI11_0/XI0/XI0_5/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN0_13 XI11_0/net21_2_ xsel_5_ XI11_0/XI0/XI0_5/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN0_12 XI11_0/net21_3_ xsel_5_ XI11_0/XI0/XI0_5/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN0_11 XI11_0/net21_4_ xsel_5_ XI11_0/XI0/XI0_5/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN0_10 XI11_0/net21_5_ xsel_5_ XI11_0/XI0/XI0_5/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN0_9 XI11_0/net21_6_ xsel_5_ XI11_0/XI0/XI0_5/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN0_8 XI11_0/net21_7_ xsel_5_ XI11_0/XI0/XI0_5/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN0_7 XI11_0/net21_8_ xsel_5_ XI11_0/XI0/XI0_5/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN0_6 XI11_0/net21_9_ xsel_5_ XI11_0/XI0/XI0_5/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN0_5 XI11_0/net21_10_ xsel_5_ XI11_0/XI0/XI0_5/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN0_4 XI11_0/net21_11_ xsel_5_ XI11_0/XI0/XI0_5/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN0_3 XI11_0/net21_12_ xsel_5_ XI11_0/XI0/XI0_5/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN0_2 XI11_0/net21_13_ xsel_5_ XI11_0/XI0/XI0_5/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN0_1 XI11_0/net21_14_ xsel_5_ XI11_0/XI0/XI0_5/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN0_0 XI11_0/net21_15_ xsel_5_ XI11_0/XI0/XI0_5/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN1_15 XI11_0/XI0/XI0_5/d__15_ xsel_5_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN1_14 XI11_0/XI0/XI0_5/d__14_ xsel_5_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN1_13 XI11_0/XI0/XI0_5/d__13_ xsel_5_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN1_12 XI11_0/XI0/XI0_5/d__12_ xsel_5_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN1_11 XI11_0/XI0/XI0_5/d__11_ xsel_5_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN1_10 XI11_0/XI0/XI0_5/d__10_ xsel_5_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN1_9 XI11_0/XI0/XI0_5/d__9_ xsel_5_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN1_8 XI11_0/XI0/XI0_5/d__8_ xsel_5_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN1_7 XI11_0/XI0/XI0_5/d__7_ xsel_5_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN1_6 XI11_0/XI0/XI0_5/d__6_ xsel_5_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN1_5 XI11_0/XI0/XI0_5/d__5_ xsel_5_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN1_4 XI11_0/XI0/XI0_5/d__4_ xsel_5_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN1_3 XI11_0/XI0/XI0_5/d__3_ xsel_5_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN1_2 XI11_0/XI0/XI0_5/d__2_ xsel_5_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN1_1 XI11_0/XI0/XI0_5/d__1_ xsel_5_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_5/MN1_0 XI11_0/XI0/XI0_5/d__0_ xsel_5_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN0_15 XI11_0/net21_0_ xsel_4_ XI11_0/XI0/XI0_4/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN0_14 XI11_0/net21_1_ xsel_4_ XI11_0/XI0/XI0_4/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN0_13 XI11_0/net21_2_ xsel_4_ XI11_0/XI0/XI0_4/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN0_12 XI11_0/net21_3_ xsel_4_ XI11_0/XI0/XI0_4/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN0_11 XI11_0/net21_4_ xsel_4_ XI11_0/XI0/XI0_4/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN0_10 XI11_0/net21_5_ xsel_4_ XI11_0/XI0/XI0_4/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN0_9 XI11_0/net21_6_ xsel_4_ XI11_0/XI0/XI0_4/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN0_8 XI11_0/net21_7_ xsel_4_ XI11_0/XI0/XI0_4/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN0_7 XI11_0/net21_8_ xsel_4_ XI11_0/XI0/XI0_4/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN0_6 XI11_0/net21_9_ xsel_4_ XI11_0/XI0/XI0_4/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN0_5 XI11_0/net21_10_ xsel_4_ XI11_0/XI0/XI0_4/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN0_4 XI11_0/net21_11_ xsel_4_ XI11_0/XI0/XI0_4/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN0_3 XI11_0/net21_12_ xsel_4_ XI11_0/XI0/XI0_4/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN0_2 XI11_0/net21_13_ xsel_4_ XI11_0/XI0/XI0_4/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN0_1 XI11_0/net21_14_ xsel_4_ XI11_0/XI0/XI0_4/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN0_0 XI11_0/net21_15_ xsel_4_ XI11_0/XI0/XI0_4/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN1_15 XI11_0/XI0/XI0_4/d__15_ xsel_4_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN1_14 XI11_0/XI0/XI0_4/d__14_ xsel_4_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN1_13 XI11_0/XI0/XI0_4/d__13_ xsel_4_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN1_12 XI11_0/XI0/XI0_4/d__12_ xsel_4_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN1_11 XI11_0/XI0/XI0_4/d__11_ xsel_4_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN1_10 XI11_0/XI0/XI0_4/d__10_ xsel_4_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN1_9 XI11_0/XI0/XI0_4/d__9_ xsel_4_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN1_8 XI11_0/XI0/XI0_4/d__8_ xsel_4_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN1_7 XI11_0/XI0/XI0_4/d__7_ xsel_4_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN1_6 XI11_0/XI0/XI0_4/d__6_ xsel_4_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN1_5 XI11_0/XI0/XI0_4/d__5_ xsel_4_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN1_4 XI11_0/XI0/XI0_4/d__4_ xsel_4_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN1_3 XI11_0/XI0/XI0_4/d__3_ xsel_4_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN1_2 XI11_0/XI0/XI0_4/d__2_ xsel_4_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN1_1 XI11_0/XI0/XI0_4/d__1_ xsel_4_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_4/MN1_0 XI11_0/XI0/XI0_4/d__0_ xsel_4_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN0_15 XI11_0/net21_0_ xsel_3_ XI11_0/XI0/XI0_3/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN0_14 XI11_0/net21_1_ xsel_3_ XI11_0/XI0/XI0_3/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN0_13 XI11_0/net21_2_ xsel_3_ XI11_0/XI0/XI0_3/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN0_12 XI11_0/net21_3_ xsel_3_ XI11_0/XI0/XI0_3/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN0_11 XI11_0/net21_4_ xsel_3_ XI11_0/XI0/XI0_3/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN0_10 XI11_0/net21_5_ xsel_3_ XI11_0/XI0/XI0_3/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN0_9 XI11_0/net21_6_ xsel_3_ XI11_0/XI0/XI0_3/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN0_8 XI11_0/net21_7_ xsel_3_ XI11_0/XI0/XI0_3/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN0_7 XI11_0/net21_8_ xsel_3_ XI11_0/XI0/XI0_3/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN0_6 XI11_0/net21_9_ xsel_3_ XI11_0/XI0/XI0_3/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN0_5 XI11_0/net21_10_ xsel_3_ XI11_0/XI0/XI0_3/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN0_4 XI11_0/net21_11_ xsel_3_ XI11_0/XI0/XI0_3/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN0_3 XI11_0/net21_12_ xsel_3_ XI11_0/XI0/XI0_3/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN0_2 XI11_0/net21_13_ xsel_3_ XI11_0/XI0/XI0_3/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN0_1 XI11_0/net21_14_ xsel_3_ XI11_0/XI0/XI0_3/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN0_0 XI11_0/net21_15_ xsel_3_ XI11_0/XI0/XI0_3/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN1_15 XI11_0/XI0/XI0_3/d__15_ xsel_3_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN1_14 XI11_0/XI0/XI0_3/d__14_ xsel_3_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN1_13 XI11_0/XI0/XI0_3/d__13_ xsel_3_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN1_12 XI11_0/XI0/XI0_3/d__12_ xsel_3_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN1_11 XI11_0/XI0/XI0_3/d__11_ xsel_3_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN1_10 XI11_0/XI0/XI0_3/d__10_ xsel_3_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN1_9 XI11_0/XI0/XI0_3/d__9_ xsel_3_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN1_8 XI11_0/XI0/XI0_3/d__8_ xsel_3_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN1_7 XI11_0/XI0/XI0_3/d__7_ xsel_3_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN1_6 XI11_0/XI0/XI0_3/d__6_ xsel_3_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN1_5 XI11_0/XI0/XI0_3/d__5_ xsel_3_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN1_4 XI11_0/XI0/XI0_3/d__4_ xsel_3_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN1_3 XI11_0/XI0/XI0_3/d__3_ xsel_3_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN1_2 XI11_0/XI0/XI0_3/d__2_ xsel_3_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN1_1 XI11_0/XI0/XI0_3/d__1_ xsel_3_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_3/MN1_0 XI11_0/XI0/XI0_3/d__0_ xsel_3_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN0_15 XI11_0/net21_0_ xsel_2_ XI11_0/XI0/XI0_2/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN0_14 XI11_0/net21_1_ xsel_2_ XI11_0/XI0/XI0_2/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN0_13 XI11_0/net21_2_ xsel_2_ XI11_0/XI0/XI0_2/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN0_12 XI11_0/net21_3_ xsel_2_ XI11_0/XI0/XI0_2/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN0_11 XI11_0/net21_4_ xsel_2_ XI11_0/XI0/XI0_2/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN0_10 XI11_0/net21_5_ xsel_2_ XI11_0/XI0/XI0_2/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN0_9 XI11_0/net21_6_ xsel_2_ XI11_0/XI0/XI0_2/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN0_8 XI11_0/net21_7_ xsel_2_ XI11_0/XI0/XI0_2/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN0_7 XI11_0/net21_8_ xsel_2_ XI11_0/XI0/XI0_2/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN0_6 XI11_0/net21_9_ xsel_2_ XI11_0/XI0/XI0_2/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN0_5 XI11_0/net21_10_ xsel_2_ XI11_0/XI0/XI0_2/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN0_4 XI11_0/net21_11_ xsel_2_ XI11_0/XI0/XI0_2/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN0_3 XI11_0/net21_12_ xsel_2_ XI11_0/XI0/XI0_2/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN0_2 XI11_0/net21_13_ xsel_2_ XI11_0/XI0/XI0_2/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN0_1 XI11_0/net21_14_ xsel_2_ XI11_0/XI0/XI0_2/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN0_0 XI11_0/net21_15_ xsel_2_ XI11_0/XI0/XI0_2/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN1_15 XI11_0/XI0/XI0_2/d__15_ xsel_2_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN1_14 XI11_0/XI0/XI0_2/d__14_ xsel_2_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN1_13 XI11_0/XI0/XI0_2/d__13_ xsel_2_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN1_12 XI11_0/XI0/XI0_2/d__12_ xsel_2_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN1_11 XI11_0/XI0/XI0_2/d__11_ xsel_2_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN1_10 XI11_0/XI0/XI0_2/d__10_ xsel_2_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN1_9 XI11_0/XI0/XI0_2/d__9_ xsel_2_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN1_8 XI11_0/XI0/XI0_2/d__8_ xsel_2_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN1_7 XI11_0/XI0/XI0_2/d__7_ xsel_2_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN1_6 XI11_0/XI0/XI0_2/d__6_ xsel_2_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN1_5 XI11_0/XI0/XI0_2/d__5_ xsel_2_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN1_4 XI11_0/XI0/XI0_2/d__4_ xsel_2_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN1_3 XI11_0/XI0/XI0_2/d__3_ xsel_2_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN1_2 XI11_0/XI0/XI0_2/d__2_ xsel_2_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN1_1 XI11_0/XI0/XI0_2/d__1_ xsel_2_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_2/MN1_0 XI11_0/XI0/XI0_2/d__0_ xsel_2_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN0_15 XI11_0/net21_0_ xsel_1_ XI11_0/XI0/XI0_1/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN0_14 XI11_0/net21_1_ xsel_1_ XI11_0/XI0/XI0_1/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN0_13 XI11_0/net21_2_ xsel_1_ XI11_0/XI0/XI0_1/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN0_12 XI11_0/net21_3_ xsel_1_ XI11_0/XI0/XI0_1/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN0_11 XI11_0/net21_4_ xsel_1_ XI11_0/XI0/XI0_1/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN0_10 XI11_0/net21_5_ xsel_1_ XI11_0/XI0/XI0_1/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN0_9 XI11_0/net21_6_ xsel_1_ XI11_0/XI0/XI0_1/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN0_8 XI11_0/net21_7_ xsel_1_ XI11_0/XI0/XI0_1/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN0_7 XI11_0/net21_8_ xsel_1_ XI11_0/XI0/XI0_1/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN0_6 XI11_0/net21_9_ xsel_1_ XI11_0/XI0/XI0_1/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN0_5 XI11_0/net21_10_ xsel_1_ XI11_0/XI0/XI0_1/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN0_4 XI11_0/net21_11_ xsel_1_ XI11_0/XI0/XI0_1/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN0_3 XI11_0/net21_12_ xsel_1_ XI11_0/XI0/XI0_1/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN0_2 XI11_0/net21_13_ xsel_1_ XI11_0/XI0/XI0_1/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN0_1 XI11_0/net21_14_ xsel_1_ XI11_0/XI0/XI0_1/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN0_0 XI11_0/net21_15_ xsel_1_ XI11_0/XI0/XI0_1/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN1_15 XI11_0/XI0/XI0_1/d__15_ xsel_1_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN1_14 XI11_0/XI0/XI0_1/d__14_ xsel_1_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN1_13 XI11_0/XI0/XI0_1/d__13_ xsel_1_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN1_12 XI11_0/XI0/XI0_1/d__12_ xsel_1_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN1_11 XI11_0/XI0/XI0_1/d__11_ xsel_1_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN1_10 XI11_0/XI0/XI0_1/d__10_ xsel_1_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN1_9 XI11_0/XI0/XI0_1/d__9_ xsel_1_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN1_8 XI11_0/XI0/XI0_1/d__8_ xsel_1_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN1_7 XI11_0/XI0/XI0_1/d__7_ xsel_1_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN1_6 XI11_0/XI0/XI0_1/d__6_ xsel_1_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN1_5 XI11_0/XI0/XI0_1/d__5_ xsel_1_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN1_4 XI11_0/XI0/XI0_1/d__4_ xsel_1_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN1_3 XI11_0/XI0/XI0_1/d__3_ xsel_1_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN1_2 XI11_0/XI0/XI0_1/d__2_ xsel_1_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN1_1 XI11_0/XI0/XI0_1/d__1_ xsel_1_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_1/MN1_0 XI11_0/XI0/XI0_1/d__0_ xsel_1_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN0_15 XI11_0/net21_0_ xsel_0_ XI11_0/XI0/XI0_0/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN0_14 XI11_0/net21_1_ xsel_0_ XI11_0/XI0/XI0_0/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN0_13 XI11_0/net21_2_ xsel_0_ XI11_0/XI0/XI0_0/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN0_12 XI11_0/net21_3_ xsel_0_ XI11_0/XI0/XI0_0/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN0_11 XI11_0/net21_4_ xsel_0_ XI11_0/XI0/XI0_0/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN0_10 XI11_0/net21_5_ xsel_0_ XI11_0/XI0/XI0_0/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN0_9 XI11_0/net21_6_ xsel_0_ XI11_0/XI0/XI0_0/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN0_8 XI11_0/net21_7_ xsel_0_ XI11_0/XI0/XI0_0/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN0_7 XI11_0/net21_8_ xsel_0_ XI11_0/XI0/XI0_0/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN0_6 XI11_0/net21_9_ xsel_0_ XI11_0/XI0/XI0_0/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN0_5 XI11_0/net21_10_ xsel_0_ XI11_0/XI0/XI0_0/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN0_4 XI11_0/net21_11_ xsel_0_ XI11_0/XI0/XI0_0/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN0_3 XI11_0/net21_12_ xsel_0_ XI11_0/XI0/XI0_0/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN0_2 XI11_0/net21_13_ xsel_0_ XI11_0/XI0/XI0_0/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN0_1 XI11_0/net21_14_ xsel_0_ XI11_0/XI0/XI0_0/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN0_0 XI11_0/net21_15_ xsel_0_ XI11_0/XI0/XI0_0/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN1_15 XI11_0/XI0/XI0_0/d__15_ xsel_0_ XI11_0/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN1_14 XI11_0/XI0/XI0_0/d__14_ xsel_0_ XI11_0/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN1_13 XI11_0/XI0/XI0_0/d__13_ xsel_0_ XI11_0/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN1_12 XI11_0/XI0/XI0_0/d__12_ xsel_0_ XI11_0/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN1_11 XI11_0/XI0/XI0_0/d__11_ xsel_0_ XI11_0/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN1_10 XI11_0/XI0/XI0_0/d__10_ xsel_0_ XI11_0/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN1_9 XI11_0/XI0/XI0_0/d__9_ xsel_0_ XI11_0/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN1_8 XI11_0/XI0/XI0_0/d__8_ xsel_0_ XI11_0/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN1_7 XI11_0/XI0/XI0_0/d__7_ xsel_0_ XI11_0/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN1_6 XI11_0/XI0/XI0_0/d__6_ xsel_0_ XI11_0/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN1_5 XI11_0/XI0/XI0_0/d__5_ xsel_0_ XI11_0/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN1_4 XI11_0/XI0/XI0_0/d__4_ xsel_0_ XI11_0/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN1_3 XI11_0/XI0/XI0_0/d__3_ xsel_0_ XI11_0/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN1_2 XI11_0/XI0/XI0_0/d__2_ xsel_0_ XI11_0/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN1_1 XI11_0/XI0/XI0_0/d__1_ xsel_0_ XI11_0/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_0/XI0/XI0_0/MN1_0 XI11_0/XI0/XI0_0/d__0_ xsel_0_ XI11_0/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI10/XI0/MN14 XI10/XI0/net30 vdd XI10/XI0/net81 gnd MN l=6e-07 w=5e-07 $[n18ll] 
XI10/XI0/MN5 XI10/XI0/net090 XI10/XI0/net095 XI10/XI0/net81 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI10/XI0/MN10 XI10/XI0/net81 CS XI10/XI0/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI10/XI0/MN12 XI10/XI0/net30 XI10/XI0/net044 XI10/XI0/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI10/XI0/MN11 XI10/XI0/net095 XI10/XI0/net090 XI10/XI0/net30 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI10/XI0/MN13 XI10/XI0/net78 CLK gnd gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI10/XI0/MP25 XI10/XI0/net090 CLK vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI10/XI0/MP27 XI10/XI0/net095 CLK vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI10/XI0/MP24 XI10/XI0/net090 XI10/XI0/net095 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI10/XI0/MP26 XI10/XI0/net095 XI10/XI0/net090 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI4_7/MN13 gnd XI5/XI4_7/m XI5/XI4_7/net15 gnd MN l=1.8e-07 w=7.4e-07 $[n18ll] 
XI5/XI4_7/MN14 XI5/XI4_7/net20 XI5/XI4_7/s gnd gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_7/MN12 XI5/XI4_7/net20 XI5/XI4_7/cn XI5/XI4_7/net24 gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_7/MN10 XI5/XI4_7/net15 XI5/XI4_7/c XI5/XI4_7/net24 gnd MN l=1.8e-07 w=7.4e-07 $[n18ll] 
XI5/XI4_7/MN8 XI5/XI4_7/net26 XI5/XI4_7/m gnd gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_7/MN6 XI5/XI4_7/net26 XI5/XI4_7/c XI5/XI4_7/pm gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_7/MN3 gnd DIN_7_ XI5/XI4_7/net36 gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_7/MN2 XI5/XI4_7/net36 XI5/XI4_7/cn XI5/XI4_7/pm gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_7/MP15 vdd XI5/XI4_7/s XI5/XI4_7/net60 vdd MP l=1.8e-07 w=3e-07 $[p18ll] 
XI5/XI4_7/MP11 XI5/XI4_7/net66 XI5/XI4_7/m vdd vdd MP l=1.8e-07 w=1.12e-06 $[p18ll] 
XI5/XI4_7/MP8 XI5/XI4_7/net66 XI5/XI4_7/cn XI5/XI4_7/net24 vdd MP l=1.8e-07 w=1.12e-06 $[p18ll] 
XI5/XI4_7/MP7 XI5/XI4_7/net60 XI5/XI4_7/c XI5/XI4_7/net24 vdd MP l=1.8e-07 w=3e-07 $[p18ll] 
XI5/XI4_7/MP4 XI5/XI4_7/net75 XI5/XI4_7/m vdd vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_7/MP2 XI5/XI4_7/net75 XI5/XI4_7/cn XI5/XI4_7/pm vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_7/MP100 XI5/XI4_7/net77 XI5/XI4_7/c XI5/XI4_7/pm vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_7/MP1 vdd DIN_7_ XI5/XI4_7/net77 vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_6/MN13 gnd XI5/XI4_6/m XI5/XI4_6/net15 gnd MN l=1.8e-07 w=7.4e-07 $[n18ll] 
XI5/XI4_6/MN14 XI5/XI4_6/net20 XI5/XI4_6/s gnd gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_6/MN12 XI5/XI4_6/net20 XI5/XI4_6/cn XI5/XI4_6/net24 gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_6/MN10 XI5/XI4_6/net15 XI5/XI4_6/c XI5/XI4_6/net24 gnd MN l=1.8e-07 w=7.4e-07 $[n18ll] 
XI5/XI4_6/MN8 XI5/XI4_6/net26 XI5/XI4_6/m gnd gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_6/MN6 XI5/XI4_6/net26 XI5/XI4_6/c XI5/XI4_6/pm gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_6/MN3 gnd DIN_6_ XI5/XI4_6/net36 gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_6/MN2 XI5/XI4_6/net36 XI5/XI4_6/cn XI5/XI4_6/pm gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_6/MP15 vdd XI5/XI4_6/s XI5/XI4_6/net60 vdd MP l=1.8e-07 w=3e-07 $[p18ll] 
XI5/XI4_6/MP11 XI5/XI4_6/net66 XI5/XI4_6/m vdd vdd MP l=1.8e-07 w=1.12e-06 $[p18ll] 
XI5/XI4_6/MP8 XI5/XI4_6/net66 XI5/XI4_6/cn XI5/XI4_6/net24 vdd MP l=1.8e-07 w=1.12e-06 $[p18ll] 
XI5/XI4_6/MP7 XI5/XI4_6/net60 XI5/XI4_6/c XI5/XI4_6/net24 vdd MP l=1.8e-07 w=3e-07 $[p18ll] 
XI5/XI4_6/MP4 XI5/XI4_6/net75 XI5/XI4_6/m vdd vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_6/MP2 XI5/XI4_6/net75 XI5/XI4_6/cn XI5/XI4_6/pm vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_6/MP100 XI5/XI4_6/net77 XI5/XI4_6/c XI5/XI4_6/pm vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_6/MP1 vdd DIN_6_ XI5/XI4_6/net77 vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_5/MN13 gnd XI5/XI4_5/m XI5/XI4_5/net15 gnd MN l=1.8e-07 w=7.4e-07 $[n18ll] 
XI5/XI4_5/MN14 XI5/XI4_5/net20 XI5/XI4_5/s gnd gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_5/MN12 XI5/XI4_5/net20 XI5/XI4_5/cn XI5/XI4_5/net24 gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_5/MN10 XI5/XI4_5/net15 XI5/XI4_5/c XI5/XI4_5/net24 gnd MN l=1.8e-07 w=7.4e-07 $[n18ll] 
XI5/XI4_5/MN8 XI5/XI4_5/net26 XI5/XI4_5/m gnd gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_5/MN6 XI5/XI4_5/net26 XI5/XI4_5/c XI5/XI4_5/pm gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_5/MN3 gnd DIN_5_ XI5/XI4_5/net36 gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_5/MN2 XI5/XI4_5/net36 XI5/XI4_5/cn XI5/XI4_5/pm gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_5/MP15 vdd XI5/XI4_5/s XI5/XI4_5/net60 vdd MP l=1.8e-07 w=3e-07 $[p18ll] 
XI5/XI4_5/MP11 XI5/XI4_5/net66 XI5/XI4_5/m vdd vdd MP l=1.8e-07 w=1.12e-06 $[p18ll] 
XI5/XI4_5/MP8 XI5/XI4_5/net66 XI5/XI4_5/cn XI5/XI4_5/net24 vdd MP l=1.8e-07 w=1.12e-06 $[p18ll] 
XI5/XI4_5/MP7 XI5/XI4_5/net60 XI5/XI4_5/c XI5/XI4_5/net24 vdd MP l=1.8e-07 w=3e-07 $[p18ll] 
XI5/XI4_5/MP4 XI5/XI4_5/net75 XI5/XI4_5/m vdd vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_5/MP2 XI5/XI4_5/net75 XI5/XI4_5/cn XI5/XI4_5/pm vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_5/MP100 XI5/XI4_5/net77 XI5/XI4_5/c XI5/XI4_5/pm vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_5/MP1 vdd DIN_5_ XI5/XI4_5/net77 vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_4/MN13 gnd XI5/XI4_4/m XI5/XI4_4/net15 gnd MN l=1.8e-07 w=7.4e-07 $[n18ll] 
XI5/XI4_4/MN14 XI5/XI4_4/net20 XI5/XI4_4/s gnd gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_4/MN12 XI5/XI4_4/net20 XI5/XI4_4/cn XI5/XI4_4/net24 gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_4/MN10 XI5/XI4_4/net15 XI5/XI4_4/c XI5/XI4_4/net24 gnd MN l=1.8e-07 w=7.4e-07 $[n18ll] 
XI5/XI4_4/MN8 XI5/XI4_4/net26 XI5/XI4_4/m gnd gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_4/MN6 XI5/XI4_4/net26 XI5/XI4_4/c XI5/XI4_4/pm gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_4/MN3 gnd DIN_4_ XI5/XI4_4/net36 gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_4/MN2 XI5/XI4_4/net36 XI5/XI4_4/cn XI5/XI4_4/pm gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_4/MP15 vdd XI5/XI4_4/s XI5/XI4_4/net60 vdd MP l=1.8e-07 w=3e-07 $[p18ll] 
XI5/XI4_4/MP11 XI5/XI4_4/net66 XI5/XI4_4/m vdd vdd MP l=1.8e-07 w=1.12e-06 $[p18ll] 
XI5/XI4_4/MP8 XI5/XI4_4/net66 XI5/XI4_4/cn XI5/XI4_4/net24 vdd MP l=1.8e-07 w=1.12e-06 $[p18ll] 
XI5/XI4_4/MP7 XI5/XI4_4/net60 XI5/XI4_4/c XI5/XI4_4/net24 vdd MP l=1.8e-07 w=3e-07 $[p18ll] 
XI5/XI4_4/MP4 XI5/XI4_4/net75 XI5/XI4_4/m vdd vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_4/MP2 XI5/XI4_4/net75 XI5/XI4_4/cn XI5/XI4_4/pm vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_4/MP100 XI5/XI4_4/net77 XI5/XI4_4/c XI5/XI4_4/pm vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_4/MP1 vdd DIN_4_ XI5/XI4_4/net77 vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_3/MN13 gnd XI5/XI4_3/m XI5/XI4_3/net15 gnd MN l=1.8e-07 w=7.4e-07 $[n18ll] 
XI5/XI4_3/MN14 XI5/XI4_3/net20 XI5/XI4_3/s gnd gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_3/MN12 XI5/XI4_3/net20 XI5/XI4_3/cn XI5/XI4_3/net24 gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_3/MN10 XI5/XI4_3/net15 XI5/XI4_3/c XI5/XI4_3/net24 gnd MN l=1.8e-07 w=7.4e-07 $[n18ll] 
XI5/XI4_3/MN8 XI5/XI4_3/net26 XI5/XI4_3/m gnd gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_3/MN6 XI5/XI4_3/net26 XI5/XI4_3/c XI5/XI4_3/pm gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_3/MN3 gnd DIN_3_ XI5/XI4_3/net36 gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_3/MN2 XI5/XI4_3/net36 XI5/XI4_3/cn XI5/XI4_3/pm gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_3/MP15 vdd XI5/XI4_3/s XI5/XI4_3/net60 vdd MP l=1.8e-07 w=3e-07 $[p18ll] 
XI5/XI4_3/MP11 XI5/XI4_3/net66 XI5/XI4_3/m vdd vdd MP l=1.8e-07 w=1.12e-06 $[p18ll] 
XI5/XI4_3/MP8 XI5/XI4_3/net66 XI5/XI4_3/cn XI5/XI4_3/net24 vdd MP l=1.8e-07 w=1.12e-06 $[p18ll] 
XI5/XI4_3/MP7 XI5/XI4_3/net60 XI5/XI4_3/c XI5/XI4_3/net24 vdd MP l=1.8e-07 w=3e-07 $[p18ll] 
XI5/XI4_3/MP4 XI5/XI4_3/net75 XI5/XI4_3/m vdd vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_3/MP2 XI5/XI4_3/net75 XI5/XI4_3/cn XI5/XI4_3/pm vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_3/MP100 XI5/XI4_3/net77 XI5/XI4_3/c XI5/XI4_3/pm vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_3/MP1 vdd DIN_3_ XI5/XI4_3/net77 vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_2/MN13 gnd XI5/XI4_2/m XI5/XI4_2/net15 gnd MN l=1.8e-07 w=7.4e-07 $[n18ll] 
XI5/XI4_2/MN14 XI5/XI4_2/net20 XI5/XI4_2/s gnd gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_2/MN12 XI5/XI4_2/net20 XI5/XI4_2/cn XI5/XI4_2/net24 gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_2/MN10 XI5/XI4_2/net15 XI5/XI4_2/c XI5/XI4_2/net24 gnd MN l=1.8e-07 w=7.4e-07 $[n18ll] 
XI5/XI4_2/MN8 XI5/XI4_2/net26 XI5/XI4_2/m gnd gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_2/MN6 XI5/XI4_2/net26 XI5/XI4_2/c XI5/XI4_2/pm gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_2/MN3 gnd DIN_2_ XI5/XI4_2/net36 gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_2/MN2 XI5/XI4_2/net36 XI5/XI4_2/cn XI5/XI4_2/pm gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_2/MP15 vdd XI5/XI4_2/s XI5/XI4_2/net60 vdd MP l=1.8e-07 w=3e-07 $[p18ll] 
XI5/XI4_2/MP11 XI5/XI4_2/net66 XI5/XI4_2/m vdd vdd MP l=1.8e-07 w=1.12e-06 $[p18ll] 
XI5/XI4_2/MP8 XI5/XI4_2/net66 XI5/XI4_2/cn XI5/XI4_2/net24 vdd MP l=1.8e-07 w=1.12e-06 $[p18ll] 
XI5/XI4_2/MP7 XI5/XI4_2/net60 XI5/XI4_2/c XI5/XI4_2/net24 vdd MP l=1.8e-07 w=3e-07 $[p18ll] 
XI5/XI4_2/MP4 XI5/XI4_2/net75 XI5/XI4_2/m vdd vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_2/MP2 XI5/XI4_2/net75 XI5/XI4_2/cn XI5/XI4_2/pm vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_2/MP100 XI5/XI4_2/net77 XI5/XI4_2/c XI5/XI4_2/pm vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_2/MP1 vdd DIN_2_ XI5/XI4_2/net77 vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_1/MN13 gnd XI5/XI4_1/m XI5/XI4_1/net15 gnd MN l=1.8e-07 w=7.4e-07 $[n18ll] 
XI5/XI4_1/MN14 XI5/XI4_1/net20 XI5/XI4_1/s gnd gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_1/MN12 XI5/XI4_1/net20 XI5/XI4_1/cn XI5/XI4_1/net24 gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_1/MN10 XI5/XI4_1/net15 XI5/XI4_1/c XI5/XI4_1/net24 gnd MN l=1.8e-07 w=7.4e-07 $[n18ll] 
XI5/XI4_1/MN8 XI5/XI4_1/net26 XI5/XI4_1/m gnd gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_1/MN6 XI5/XI4_1/net26 XI5/XI4_1/c XI5/XI4_1/pm gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_1/MN3 gnd DIN_1_ XI5/XI4_1/net36 gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_1/MN2 XI5/XI4_1/net36 XI5/XI4_1/cn XI5/XI4_1/pm gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_1/MP15 vdd XI5/XI4_1/s XI5/XI4_1/net60 vdd MP l=1.8e-07 w=3e-07 $[p18ll] 
XI5/XI4_1/MP11 XI5/XI4_1/net66 XI5/XI4_1/m vdd vdd MP l=1.8e-07 w=1.12e-06 $[p18ll] 
XI5/XI4_1/MP8 XI5/XI4_1/net66 XI5/XI4_1/cn XI5/XI4_1/net24 vdd MP l=1.8e-07 w=1.12e-06 $[p18ll] 
XI5/XI4_1/MP7 XI5/XI4_1/net60 XI5/XI4_1/c XI5/XI4_1/net24 vdd MP l=1.8e-07 w=3e-07 $[p18ll] 
XI5/XI4_1/MP4 XI5/XI4_1/net75 XI5/XI4_1/m vdd vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_1/MP2 XI5/XI4_1/net75 XI5/XI4_1/cn XI5/XI4_1/pm vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_1/MP100 XI5/XI4_1/net77 XI5/XI4_1/c XI5/XI4_1/pm vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_1/MP1 vdd DIN_1_ XI5/XI4_1/net77 vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_0/MN13 gnd XI5/XI4_0/m XI5/XI4_0/net15 gnd MN l=1.8e-07 w=7.4e-07 $[n18ll] 
XI5/XI4_0/MN14 XI5/XI4_0/net20 XI5/XI4_0/s gnd gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_0/MN12 XI5/XI4_0/net20 XI5/XI4_0/cn XI5/XI4_0/net24 gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_0/MN10 XI5/XI4_0/net15 XI5/XI4_0/c XI5/XI4_0/net24 gnd MN l=1.8e-07 w=7.4e-07 $[n18ll] 
XI5/XI4_0/MN8 XI5/XI4_0/net26 XI5/XI4_0/m gnd gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_0/MN6 XI5/XI4_0/net26 XI5/XI4_0/c XI5/XI4_0/pm gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_0/MN3 gnd DIN_0_ XI5/XI4_0/net36 gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_0/MN2 XI5/XI4_0/net36 XI5/XI4_0/cn XI5/XI4_0/pm gnd MN l=1.8e-07 w=3e-07 $[n18ll] 
XI5/XI4_0/MP15 vdd XI5/XI4_0/s XI5/XI4_0/net60 vdd MP l=1.8e-07 w=3e-07 $[p18ll] 
XI5/XI4_0/MP11 XI5/XI4_0/net66 XI5/XI4_0/m vdd vdd MP l=1.8e-07 w=1.12e-06 $[p18ll] 
XI5/XI4_0/MP8 XI5/XI4_0/net66 XI5/XI4_0/cn XI5/XI4_0/net24 vdd MP l=1.8e-07 w=1.12e-06 $[p18ll] 
XI5/XI4_0/MP7 XI5/XI4_0/net60 XI5/XI4_0/c XI5/XI4_0/net24 vdd MP l=1.8e-07 w=3e-07 $[p18ll] 
XI5/XI4_0/MP4 XI5/XI4_0/net75 XI5/XI4_0/m vdd vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_0/MP2 XI5/XI4_0/net75 XI5/XI4_0/cn XI5/XI4_0/pm vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_0/MP100 XI5/XI4_0/net77 XI5/XI4_0/c XI5/XI4_0/pm vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI4_0/MP1 vdd DIN_0_ XI5/XI4_0/net77 vdd MP l=1.8e-07 w=4.2e-07 $[p18ll] 
XI5/XI2/MN14 XI5/XI2/net30 vdd XI5/XI2/net81 gnd MN l=6e-07 w=5e-07 $[n18ll] 
XI5/XI2/MN5 XI5/XI2/net090 XI5/XI2/net095 XI5/XI2/net81 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI2/MN10 XI5/XI2/net81 RD XI5/XI2/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI2/MN12 XI5/XI2/net30 XI5/XI2/net044 XI5/XI2/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI2/MN11 XI5/XI2/net095 XI5/XI2/net090 XI5/XI2/net30 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI2/MN13 XI5/XI2/net78 XI5/ck gnd gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI2/MP25 XI5/XI2/net090 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI2/MP27 XI5/XI2/net095 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI2/MP24 XI5/XI2/net090 XI5/XI2/net095 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI2/MP26 XI5/XI2/net095 XI5/XI2/net090 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI1/MN14 XI5/XI1/net30 vdd XI5/XI1/net81 gnd MN l=6e-07 w=5e-07 $[n18ll] 
XI5/XI1/MN5 XI5/XI1/net090 XI5/XI1/net095 XI5/XI1/net81 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI1/MN10 XI5/XI1/net81 WR XI5/XI1/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI1/MN12 XI5/XI1/net30 XI5/XI1/net044 XI5/XI1/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI1/MN11 XI5/XI1/net095 XI5/XI1/net090 XI5/XI1/net30 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI1/MN13 XI5/XI1/net78 XI5/ck gnd gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI1/MP25 XI5/XI1/net090 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI1/MP27 XI5/XI1/net095 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI1/MP24 XI5/XI1/net090 XI5/XI1/net095 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI1/MP26 XI5/XI1/net095 XI5/XI1/net090 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_9/MN14 XI5/XI0_9/net30 vdd XI5/XI0_9/net81 gnd MN l=6e-07 w=5e-07 $[n18ll] 
XI5/XI0_9/MN5 XI5/XI0_9/net090 XI5/XI0_9/net095 XI5/XI0_9/net81 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_9/MN10 XI5/XI0_9/net81 A_9_ XI5/XI0_9/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_9/MN12 XI5/XI0_9/net30 XI5/XI0_9/net044 XI5/XI0_9/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_9/MN11 XI5/XI0_9/net095 XI5/XI0_9/net090 XI5/XI0_9/net30 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_9/MN13 XI5/XI0_9/net78 XI5/ck gnd gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_9/MP25 XI5/XI0_9/net090 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_9/MP27 XI5/XI0_9/net095 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_9/MP24 XI5/XI0_9/net090 XI5/XI0_9/net095 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_9/MP26 XI5/XI0_9/net095 XI5/XI0_9/net090 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_8/MN14 XI5/XI0_8/net30 vdd XI5/XI0_8/net81 gnd MN l=6e-07 w=5e-07 $[n18ll] 
XI5/XI0_8/MN5 XI5/XI0_8/net090 XI5/XI0_8/net095 XI5/XI0_8/net81 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_8/MN10 XI5/XI0_8/net81 A_8_ XI5/XI0_8/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_8/MN12 XI5/XI0_8/net30 XI5/XI0_8/net044 XI5/XI0_8/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_8/MN11 XI5/XI0_8/net095 XI5/XI0_8/net090 XI5/XI0_8/net30 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_8/MN13 XI5/XI0_8/net78 XI5/ck gnd gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_8/MP25 XI5/XI0_8/net090 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_8/MP27 XI5/XI0_8/net095 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_8/MP24 XI5/XI0_8/net090 XI5/XI0_8/net095 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_8/MP26 XI5/XI0_8/net095 XI5/XI0_8/net090 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_7/MN14 XI5/XI0_7/net30 vdd XI5/XI0_7/net81 gnd MN l=6e-07 w=5e-07 $[n18ll] 
XI5/XI0_7/MN5 XI5/XI0_7/net090 XI5/XI0_7/net095 XI5/XI0_7/net81 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_7/MN10 XI5/XI0_7/net81 A_7_ XI5/XI0_7/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_7/MN12 XI5/XI0_7/net30 XI5/XI0_7/net044 XI5/XI0_7/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_7/MN11 XI5/XI0_7/net095 XI5/XI0_7/net090 XI5/XI0_7/net30 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_7/MN13 XI5/XI0_7/net78 XI5/ck gnd gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_7/MP25 XI5/XI0_7/net090 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_7/MP27 XI5/XI0_7/net095 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_7/MP24 XI5/XI0_7/net090 XI5/XI0_7/net095 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_7/MP26 XI5/XI0_7/net095 XI5/XI0_7/net090 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_6/MN14 XI5/XI0_6/net30 vdd XI5/XI0_6/net81 gnd MN l=6e-07 w=5e-07 $[n18ll] 
XI5/XI0_6/MN5 XI5/XI0_6/net090 XI5/XI0_6/net095 XI5/XI0_6/net81 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_6/MN10 XI5/XI0_6/net81 A_6_ XI5/XI0_6/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_6/MN12 XI5/XI0_6/net30 XI5/XI0_6/net044 XI5/XI0_6/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_6/MN11 XI5/XI0_6/net095 XI5/XI0_6/net090 XI5/XI0_6/net30 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_6/MN13 XI5/XI0_6/net78 XI5/ck gnd gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_6/MP25 XI5/XI0_6/net090 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_6/MP27 XI5/XI0_6/net095 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_6/MP24 XI5/XI0_6/net090 XI5/XI0_6/net095 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_6/MP26 XI5/XI0_6/net095 XI5/XI0_6/net090 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_5/MN14 XI5/XI0_5/net30 vdd XI5/XI0_5/net81 gnd MN l=6e-07 w=5e-07 $[n18ll] 
XI5/XI0_5/MN5 XI5/XI0_5/net090 XI5/XI0_5/net095 XI5/XI0_5/net81 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_5/MN10 XI5/XI0_5/net81 A_5_ XI5/XI0_5/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_5/MN12 XI5/XI0_5/net30 XI5/XI0_5/net044 XI5/XI0_5/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_5/MN11 XI5/XI0_5/net095 XI5/XI0_5/net090 XI5/XI0_5/net30 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_5/MN13 XI5/XI0_5/net78 XI5/ck gnd gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_5/MP25 XI5/XI0_5/net090 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_5/MP27 XI5/XI0_5/net095 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_5/MP24 XI5/XI0_5/net090 XI5/XI0_5/net095 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_5/MP26 XI5/XI0_5/net095 XI5/XI0_5/net090 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_4/MN14 XI5/XI0_4/net30 vdd XI5/XI0_4/net81 gnd MN l=6e-07 w=5e-07 $[n18ll] 
XI5/XI0_4/MN5 XI5/XI0_4/net090 XI5/XI0_4/net095 XI5/XI0_4/net81 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_4/MN10 XI5/XI0_4/net81 A_4_ XI5/XI0_4/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_4/MN12 XI5/XI0_4/net30 XI5/XI0_4/net044 XI5/XI0_4/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_4/MN11 XI5/XI0_4/net095 XI5/XI0_4/net090 XI5/XI0_4/net30 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_4/MN13 XI5/XI0_4/net78 XI5/ck gnd gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_4/MP25 XI5/XI0_4/net090 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_4/MP27 XI5/XI0_4/net095 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_4/MP24 XI5/XI0_4/net090 XI5/XI0_4/net095 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_4/MP26 XI5/XI0_4/net095 XI5/XI0_4/net090 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_3/MN14 XI5/XI0_3/net30 vdd XI5/XI0_3/net81 gnd MN l=6e-07 w=5e-07 $[n18ll] 
XI5/XI0_3/MN5 XI5/XI0_3/net090 XI5/XI0_3/net095 XI5/XI0_3/net81 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_3/MN10 XI5/XI0_3/net81 A_3_ XI5/XI0_3/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_3/MN12 XI5/XI0_3/net30 XI5/XI0_3/net044 XI5/XI0_3/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_3/MN11 XI5/XI0_3/net095 XI5/XI0_3/net090 XI5/XI0_3/net30 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_3/MN13 XI5/XI0_3/net78 XI5/ck gnd gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_3/MP25 XI5/XI0_3/net090 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_3/MP27 XI5/XI0_3/net095 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_3/MP24 XI5/XI0_3/net090 XI5/XI0_3/net095 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_3/MP26 XI5/XI0_3/net095 XI5/XI0_3/net090 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_2/MN14 XI5/XI0_2/net30 vdd XI5/XI0_2/net81 gnd MN l=6e-07 w=5e-07 $[n18ll] 
XI5/XI0_2/MN5 XI5/XI0_2/net090 XI5/XI0_2/net095 XI5/XI0_2/net81 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_2/MN10 XI5/XI0_2/net81 A_2_ XI5/XI0_2/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_2/MN12 XI5/XI0_2/net30 XI5/XI0_2/net044 XI5/XI0_2/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_2/MN11 XI5/XI0_2/net095 XI5/XI0_2/net090 XI5/XI0_2/net30 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_2/MN13 XI5/XI0_2/net78 XI5/ck gnd gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_2/MP25 XI5/XI0_2/net090 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_2/MP27 XI5/XI0_2/net095 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_2/MP24 XI5/XI0_2/net090 XI5/XI0_2/net095 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_2/MP26 XI5/XI0_2/net095 XI5/XI0_2/net090 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_1/MN14 XI5/XI0_1/net30 vdd XI5/XI0_1/net81 gnd MN l=6e-07 w=5e-07 $[n18ll] 
XI5/XI0_1/MN5 XI5/XI0_1/net090 XI5/XI0_1/net095 XI5/XI0_1/net81 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_1/MN10 XI5/XI0_1/net81 A_1_ XI5/XI0_1/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_1/MN12 XI5/XI0_1/net30 XI5/XI0_1/net044 XI5/XI0_1/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_1/MN11 XI5/XI0_1/net095 XI5/XI0_1/net090 XI5/XI0_1/net30 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_1/MN13 XI5/XI0_1/net78 XI5/ck gnd gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_1/MP25 XI5/XI0_1/net090 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_1/MP27 XI5/XI0_1/net095 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_1/MP24 XI5/XI0_1/net090 XI5/XI0_1/net095 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_1/MP26 XI5/XI0_1/net095 XI5/XI0_1/net090 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_0/MN14 XI5/XI0_0/net30 vdd XI5/XI0_0/net81 gnd MN l=6e-07 w=5e-07 $[n18ll] 
XI5/XI0_0/MN5 XI5/XI0_0/net090 XI5/XI0_0/net095 XI5/XI0_0/net81 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_0/MN10 XI5/XI0_0/net81 A_0_ XI5/XI0_0/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_0/MN12 XI5/XI0_0/net30 XI5/XI0_0/net044 XI5/XI0_0/net78 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_0/MN11 XI5/XI0_0/net095 XI5/XI0_0/net090 XI5/XI0_0/net30 gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_0/MN13 XI5/XI0_0/net78 XI5/ck gnd gnd MN l=1.8e-07 w=1.2e-06 $[n18ll] 
XI5/XI0_0/MP25 XI5/XI0_0/net090 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_0/MP27 XI5/XI0_0/net095 XI5/ck vdd vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI5/XI0_0/MP24 XI5/XI0_0/net090 XI5/XI0_0/net095 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XI5/XI0_0/MP26 XI5/XI0_0/net095 XI5/XI0_0/net090 vdd vdd MP l=1.8e-07 w=1e-06 $[p18ll] 
XG1 sck_bar XI11_7/XI3/net7 XI11_7/XI3/net17 DECAP_NAND2_G1
XG2 XI11_7/XI4/data_out_ rd_en XI11_7/XI4/net063 DECAP_NAND2_G2
XG3 wr_en wrdata_7_ XI11_7/XI4/net26 DECAP_NAND2_G2
XG4 wr_en wrdata__7_ XI11_7/XI4/net8 DECAP_NAND2_G2
XG5 wr_en wrdata__7_ XI11_7/XI4/net20 DECAP_NAND2_G2
XG6 wr_en wrdata_7_ XI11_7/XI4/net23 DECAP_NAND2_G2
XG7 rd_en XI11_7/XI4/data_out XI11_7/XI4/net090 DECAP_NAND2_G2
XG8 sck_bar XI11_6/XI3/net7 XI11_6/XI3/net17 DECAP_NAND2_G1
XG9 rd_en XI11_6/XI4/data_out_ XI11_6/XI4/net063 DECAP_NAND2_G2
XG10 wr_en wrdata_6_ XI11_6/XI4/net26 DECAP_NAND2_G2
XG11 wr_en wrdata__6_ XI11_6/XI4/net8 DECAP_NAND2_G2
XG12 wr_en wrdata__6_ XI11_6/XI4/net20 DECAP_NAND2_G2
XG13 wr_en wrdata_6_ XI11_6/XI4/net23 DECAP_NAND2_G2
XG14 rd_en XI11_6/XI4/data_out XI11_6/XI4/net090 DECAP_NAND2_G2
XG15 sck_bar XI11_5/XI3/net7 XI11_5/XI3/net17 DECAP_NAND2_G1
XG16 rd_en XI11_5/XI4/data_out_ XI11_5/XI4/net063 DECAP_NAND2_G2
XG17 wr_en wrdata_5_ XI11_5/XI4/net26 DECAP_NAND2_G2
XG18 wr_en wrdata__5_ XI11_5/XI4/net8 DECAP_NAND2_G2
XG19 wr_en wrdata__5_ XI11_5/XI4/net20 DECAP_NAND2_G2
XG20 wr_en wrdata_5_ XI11_5/XI4/net23 DECAP_NAND2_G2
XG21 rd_en XI11_5/XI4/data_out XI11_5/XI4/net090 DECAP_NAND2_G2
XG22 sck_bar XI11_4/XI3/net7 XI11_4/XI3/net17 DECAP_NAND2_G1
XG23 rd_en XI11_4/XI4/data_out_ XI11_4/XI4/net063 DECAP_NAND2_G2
XG24 wr_en wrdata_4_ XI11_4/XI4/net26 DECAP_NAND2_G2
XG25 wr_en wrdata__4_ XI11_4/XI4/net8 DECAP_NAND2_G2
XG26 wr_en wrdata__4_ XI11_4/XI4/net20 DECAP_NAND2_G2
XG27 wr_en wrdata_4_ XI11_4/XI4/net23 DECAP_NAND2_G2
XG28 rd_en XI11_4/XI4/data_out XI11_4/XI4/net090 DECAP_NAND2_G2
XG29 sck_bar XI11_3/XI3/net7 XI11_3/XI3/net17 DECAP_NAND2_G1
XG30 rd_en XI11_3/XI4/data_out_ XI11_3/XI4/net063 DECAP_NAND2_G2
XG31 wr_en wrdata_3_ XI11_3/XI4/net26 DECAP_NAND2_G2
XG32 wr_en wrdata__3_ XI11_3/XI4/net8 DECAP_NAND2_G2
XG33 wr_en wrdata__3_ XI11_3/XI4/net20 DECAP_NAND2_G2
XG34 wr_en wrdata_3_ XI11_3/XI4/net23 DECAP_NAND2_G2
XG35 rd_en XI11_3/XI4/data_out XI11_3/XI4/net090 DECAP_NAND2_G2
XG36 sck_bar XI11_2/XI3/net7 XI11_2/XI3/net17 DECAP_NAND2_G1
XG37 rd_en XI11_2/XI4/data_out_ XI11_2/XI4/net063 DECAP_NAND2_G2
XG38 wr_en wrdata_2_ XI11_2/XI4/net26 DECAP_NAND2_G2
XG39 wr_en wrdata__2_ XI11_2/XI4/net8 DECAP_NAND2_G2
XG40 wr_en wrdata__2_ XI11_2/XI4/net20 DECAP_NAND2_G2
XG41 wr_en wrdata_2_ XI11_2/XI4/net23 DECAP_NAND2_G2
XG42 rd_en XI11_2/XI4/data_out XI11_2/XI4/net090 DECAP_NAND2_G2
XG43 sck_bar XI11_1/XI3/net7 XI11_1/XI3/net17 DECAP_NAND2_G1
XG44 rd_en XI11_1/XI4/data_out_ XI11_1/XI4/net063 DECAP_NAND2_G2
XG45 wr_en wrdata_1_ XI11_1/XI4/net26 DECAP_NAND2_G2
XG46 wr_en wrdata__1_ XI11_1/XI4/net8 DECAP_NAND2_G2
XG47 wr_en wrdata__1_ XI11_1/XI4/net20 DECAP_NAND2_G2
XG48 wr_en wrdata_1_ XI11_1/XI4/net23 DECAP_NAND2_G2
XG49 rd_en XI11_1/XI4/data_out XI11_1/XI4/net090 DECAP_NAND2_G2
XG50 sck_bar XI11_0/XI3/net7 XI11_0/XI3/net17 DECAP_NAND2_G1
XG51 rd_en XI11_0/XI4/data_out_ XI11_0/XI4/net063 DECAP_NAND2_G2
XG52 wr_en wrdata_0_ XI11_0/XI4/net26 DECAP_NAND2_G2
XG53 wr_en wrdata__0_ XI11_0/XI4/net8 DECAP_NAND2_G2
XG54 wr_en wrdata__0_ XI11_0/XI4/net20 DECAP_NAND2_G2
XG55 wr_en wrdata_0_ XI11_0/XI4/net23 DECAP_NAND2_G2
XG56 rd_en XI11_0/XI4/data_out XI11_0/XI4/net090 DECAP_NAND2_G2
XG57 XI2/net029_0_ XI2/net026_0_ XI2/net024_0_ DECAP_NOR2_G3
XG58 XI2/net029_1_ XI2/net026_1_ XI2/net024_1_ DECAP_NOR2_G3
XG59 XI2/net029_2_ XI2/net026_2_ XI2/net024_2_ DECAP_NOR2_G3
XG60 XI2/net029_3_ XI2/net026_3_ XI2/net024_3_ DECAP_NOR2_G3
XG61 XI2/net029_4_ XI2/net026_4_ XI2/net024_4_ DECAP_NOR2_G3
XG62 XI2/net029_5_ XI2/net026_5_ XI2/net024_5_ DECAP_NOR2_G3
XG63 XI2/net029_6_ XI2/net026_6_ XI2/net024_6_ DECAP_NOR2_G3
XG64 XI2/net029_7_ XI2/net026_7_ XI2/net024_7_ DECAP_NOR2_G3
XG65 XI2/net029_8_ XI2/net026_8_ XI2/net024_8_ DECAP_NOR2_G3
XG66 XI2/net029_9_ XI2/net026_9_ XI2/net024_9_ DECAP_NOR2_G3
XG67 XI2/net029_10_ XI2/net026_10_ XI2/net024_10_ DECAP_NOR2_G3
XG68 XI2/net029_11_ XI2/net026_11_ XI2/net024_11_ DECAP_NOR2_G3
XG69 XI2/net029_12_ XI2/net026_12_ XI2/net024_12_ DECAP_NOR2_G3
XG70 XI2/net029_13_ XI2/net026_13_ XI2/net024_13_ DECAP_NOR2_G3
XG71 XI2/net029_14_ XI2/net026_14_ XI2/net024_14_ DECAP_NOR2_G3
XG72 XI2/net029_15_ XI2/net026_15_ XI2/net024_15_ DECAP_NOR2_G3
XG73 XI2/net029_16_ XI2/net026_16_ XI2/net024_16_ DECAP_NOR2_G3
XG74 XI2/net029_17_ XI2/net026_17_ XI2/net024_17_ DECAP_NOR2_G3
XG75 XI2/net029_18_ XI2/net026_18_ XI2/net024_18_ DECAP_NOR2_G3
XG76 XI2/net029_19_ XI2/net026_19_ XI2/net024_19_ DECAP_NOR2_G3
XG77 XI2/net029_20_ XI2/net026_20_ XI2/net024_20_ DECAP_NOR2_G3
XG78 XI2/net029_21_ XI2/net026_21_ XI2/net024_21_ DECAP_NOR2_G3
XG79 XI2/net029_22_ XI2/net026_22_ XI2/net024_22_ DECAP_NOR2_G3
XG80 XI2/net029_23_ XI2/net026_23_ XI2/net024_23_ DECAP_NOR2_G3
XG81 XI2/net029_24_ XI2/net026_24_ XI2/net024_24_ DECAP_NOR2_G3
XG82 XI2/net029_25_ XI2/net026_25_ XI2/net024_25_ DECAP_NOR2_G3
XG83 XI2/net029_26_ XI2/net026_26_ XI2/net024_26_ DECAP_NOR2_G3
XG84 XI2/net029_27_ XI2/net026_27_ XI2/net024_27_ DECAP_NOR2_G3
XG85 XI2/net029_28_ XI2/net026_28_ XI2/net024_28_ DECAP_NOR2_G3
XG86 XI2/net029_29_ XI2/net026_29_ XI2/net024_29_ DECAP_NOR2_G3
XG87 XI2/net029_30_ XI2/net026_30_ XI2/net024_30_ DECAP_NOR2_G3
XG88 XI2/net029_31_ XI2/net026_31_ XI2/net024_31_ DECAP_NOR2_G3
XG89 XI2/net029_32_ XI2/net026_32_ XI2/net024_32_ DECAP_NOR2_G3
XG90 XI2/net029_33_ XI2/net026_33_ XI2/net024_33_ DECAP_NOR2_G3
XG91 XI2/net029_34_ XI2/net026_34_ XI2/net024_34_ DECAP_NOR2_G3
XG92 XI2/net029_35_ XI2/net026_35_ XI2/net024_35_ DECAP_NOR2_G3
XG93 XI2/net029_36_ XI2/net026_36_ XI2/net024_36_ DECAP_NOR2_G3
XG94 XI2/net029_37_ XI2/net026_37_ XI2/net024_37_ DECAP_NOR2_G3
XG95 XI2/net029_38_ XI2/net026_38_ XI2/net024_38_ DECAP_NOR2_G3
XG96 XI2/net029_39_ XI2/net026_39_ XI2/net024_39_ DECAP_NOR2_G3
XG97 XI2/net029_40_ XI2/net026_40_ XI2/net024_40_ DECAP_NOR2_G3
XG98 XI2/net029_41_ XI2/net026_41_ XI2/net024_41_ DECAP_NOR2_G3
XG99 XI2/net029_42_ XI2/net026_42_ XI2/net024_42_ DECAP_NOR2_G3
XG100 XI2/net029_43_ XI2/net026_43_ XI2/net024_43_ DECAP_NOR2_G3
XG101 XI2/net029_44_ XI2/net026_44_ XI2/net024_44_ DECAP_NOR2_G3
XG102 XI2/net029_45_ XI2/net026_45_ XI2/net024_45_ DECAP_NOR2_G3
XG103 XI2/net029_46_ XI2/net026_46_ XI2/net024_46_ DECAP_NOR2_G3
XG104 XI2/net029_47_ XI2/net026_47_ XI2/net024_47_ DECAP_NOR2_G3
XG105 XI2/net029_48_ XI2/net026_48_ XI2/net024_48_ DECAP_NOR2_G3
XG106 XI2/net029_49_ XI2/net026_49_ XI2/net024_49_ DECAP_NOR2_G3
XG107 XI2/net029_50_ XI2/net026_50_ XI2/net024_50_ DECAP_NOR2_G3
XG108 XI2/net029_51_ XI2/net026_51_ XI2/net024_51_ DECAP_NOR2_G3
XG109 XI2/net029_52_ XI2/net026_52_ XI2/net024_52_ DECAP_NOR2_G3
XG110 XI2/net029_53_ XI2/net026_53_ XI2/net024_53_ DECAP_NOR2_G3
XG111 XI2/net029_54_ XI2/net026_54_ XI2/net024_54_ DECAP_NOR2_G3
XG112 XI2/net029_55_ XI2/net026_55_ XI2/net024_55_ DECAP_NOR2_G3
XG113 XI2/net029_56_ XI2/net026_56_ XI2/net024_56_ DECAP_NOR2_G3
XG114 XI2/net029_57_ XI2/net026_57_ XI2/net024_57_ DECAP_NOR2_G3
XG115 XI2/net029_58_ XI2/net026_58_ XI2/net024_58_ DECAP_NOR2_G3
XG116 XI2/net029_59_ XI2/net026_59_ XI2/net024_59_ DECAP_NOR2_G3
XG117 XI2/net029_60_ XI2/net026_60_ XI2/net024_60_ DECAP_NOR2_G3
XG118 XI2/net029_61_ XI2/net026_61_ XI2/net024_61_ DECAP_NOR2_G3
XG119 XI2/net029_62_ XI2/net026_62_ XI2/net024_62_ DECAP_NOR2_G3
XG120 XI2/net029_63_ XI2/net026_63_ XI2/net024_63_ DECAP_NOR2_G3
XG121 addr_2_ addr_1_ addr_0_ XI2/net029_0_ DECAP_NAND3_G4
XG122 addr_2_ addr_1_ addr__0_ XI2/net029_1_ DECAP_NAND3_G4
XG123 addr_2_ addr__1_ addr_0_ XI2/net029_2_ DECAP_NAND3_G4
XG124 addr_2_ addr__1_ addr__0_ XI2/net029_3_ DECAP_NAND3_G4
XG125 addr__2_ addr_1_ addr_0_ XI2/net029_4_ DECAP_NAND3_G4
XG126 addr__2_ addr_1_ addr__0_ XI2/net029_5_ DECAP_NAND3_G4
XG127 addr__2_ addr__1_ addr_0_ XI2/net029_6_ DECAP_NAND3_G4
XG128 addr__2_ addr__1_ addr__0_ XI2/net029_7_ DECAP_NAND3_G4
XG129 addr_2_ addr_1_ addr_0_ XI2/net029_8_ DECAP_NAND3_G4
XG130 addr_2_ addr_1_ addr__0_ XI2/net029_9_ DECAP_NAND3_G4
XG131 addr_2_ addr__1_ addr_0_ XI2/net029_10_ DECAP_NAND3_G4
XG132 addr_2_ addr__1_ addr__0_ XI2/net029_11_ DECAP_NAND3_G4
XG133 addr__2_ addr_1_ addr_0_ XI2/net029_12_ DECAP_NAND3_G4
XG134 addr__2_ addr_1_ addr__0_ XI2/net029_13_ DECAP_NAND3_G4
XG135 addr__2_ addr__1_ addr_0_ XI2/net029_14_ DECAP_NAND3_G4
XG136 addr__2_ addr__1_ addr__0_ XI2/net029_15_ DECAP_NAND3_G4
XG137 addr_2_ addr_1_ addr_0_ XI2/net029_16_ DECAP_NAND3_G4
XG138 addr_2_ addr_1_ addr__0_ XI2/net029_17_ DECAP_NAND3_G4
XG139 addr_2_ addr__1_ addr_0_ XI2/net029_18_ DECAP_NAND3_G4
XG140 addr_2_ addr__1_ addr__0_ XI2/net029_19_ DECAP_NAND3_G4
XG141 addr__2_ addr_1_ addr_0_ XI2/net029_20_ DECAP_NAND3_G4
XG142 addr__2_ addr_1_ addr__0_ XI2/net029_21_ DECAP_NAND3_G4
XG143 addr__2_ addr__1_ addr_0_ XI2/net029_22_ DECAP_NAND3_G4
XG144 addr__2_ addr__1_ addr__0_ XI2/net029_23_ DECAP_NAND3_G4
XG145 addr_2_ addr_1_ addr_0_ XI2/net029_24_ DECAP_NAND3_G4
XG146 addr_2_ addr_1_ addr__0_ XI2/net029_25_ DECAP_NAND3_G4
XG147 addr_2_ addr__1_ addr_0_ XI2/net029_26_ DECAP_NAND3_G4
XG148 addr_2_ addr__1_ addr__0_ XI2/net029_27_ DECAP_NAND3_G4
XG149 addr__2_ addr_1_ addr_0_ XI2/net029_28_ DECAP_NAND3_G4
XG150 addr__2_ addr_1_ addr__0_ XI2/net029_29_ DECAP_NAND3_G4
XG151 addr__2_ addr__1_ addr_0_ XI2/net029_30_ DECAP_NAND3_G4
XG152 addr__2_ addr__1_ addr__0_ XI2/net029_31_ DECAP_NAND3_G4
XG153 addr_2_ addr_1_ addr_0_ XI2/net029_32_ DECAP_NAND3_G4
XG154 addr_2_ addr_1_ addr__0_ XI2/net029_33_ DECAP_NAND3_G4
XG155 addr_2_ addr__1_ addr_0_ XI2/net029_34_ DECAP_NAND3_G4
XG156 addr_2_ addr__1_ addr__0_ XI2/net029_35_ DECAP_NAND3_G4
XG157 addr__2_ addr_1_ addr_0_ XI2/net029_36_ DECAP_NAND3_G4
XG158 addr__2_ addr_1_ addr__0_ XI2/net029_37_ DECAP_NAND3_G4
XG159 addr__2_ addr__1_ addr_0_ XI2/net029_38_ DECAP_NAND3_G4
XG160 addr__2_ addr__1_ addr__0_ XI2/net029_39_ DECAP_NAND3_G4
XG161 addr_2_ addr_1_ addr_0_ XI2/net029_40_ DECAP_NAND3_G4
XG162 addr_2_ addr_1_ addr__0_ XI2/net029_41_ DECAP_NAND3_G4
XG163 addr_2_ addr__1_ addr_0_ XI2/net029_42_ DECAP_NAND3_G4
XG164 addr_2_ addr__1_ addr__0_ XI2/net029_43_ DECAP_NAND3_G4
XG165 addr__2_ addr_1_ addr_0_ XI2/net029_44_ DECAP_NAND3_G4
XG166 addr__2_ addr_1_ addr__0_ XI2/net029_45_ DECAP_NAND3_G4
XG167 addr__2_ addr__1_ addr_0_ XI2/net029_46_ DECAP_NAND3_G4
XG168 addr__2_ addr__1_ addr__0_ XI2/net029_47_ DECAP_NAND3_G4
XG169 addr_2_ addr_1_ addr_0_ XI2/net029_48_ DECAP_NAND3_G4
XG170 addr_2_ addr_1_ addr__0_ XI2/net029_49_ DECAP_NAND3_G4
XG171 addr_2_ addr__1_ addr_0_ XI2/net029_50_ DECAP_NAND3_G4
XG172 addr_2_ addr__1_ addr__0_ XI2/net029_51_ DECAP_NAND3_G4
XG173 addr__2_ addr_1_ addr_0_ XI2/net029_52_ DECAP_NAND3_G4
XG174 addr__2_ addr_1_ addr__0_ XI2/net029_53_ DECAP_NAND3_G4
XG175 addr__2_ addr__1_ addr_0_ XI2/net029_54_ DECAP_NAND3_G4
XG176 addr__2_ addr__1_ addr__0_ XI2/net029_55_ DECAP_NAND3_G4
XG177 addr_2_ addr_1_ addr_0_ XI2/net029_56_ DECAP_NAND3_G4
XG178 addr_2_ addr_1_ addr__0_ XI2/net029_57_ DECAP_NAND3_G4
XG179 addr_2_ addr__1_ addr_0_ XI2/net029_58_ DECAP_NAND3_G4
XG180 addr_2_ addr__1_ addr__0_ XI2/net029_59_ DECAP_NAND3_G4
XG181 addr__2_ addr_1_ addr_0_ XI2/net029_60_ DECAP_NAND3_G4
XG182 addr__2_ addr_1_ addr__0_ XI2/net029_61_ DECAP_NAND3_G4
XG183 addr__2_ addr__1_ addr_0_ XI2/net029_62_ DECAP_NAND3_G4
XG184 addr__2_ addr__1_ addr__0_ XI2/net029_63_ DECAP_NAND3_G4
XG185 addr_5_ addr_4_ addr_3_ XI2/net026_0_ DECAP_NAND3_G4
XG186 addr_5_ addr_4_ addr_3_ XI2/net026_1_ DECAP_NAND3_G4
XG187 addr_5_ addr_4_ addr_3_ XI2/net026_2_ DECAP_NAND3_G4
XG188 addr_5_ addr_4_ addr_3_ XI2/net026_3_ DECAP_NAND3_G4
XG189 addr_5_ addr_4_ addr_3_ XI2/net026_4_ DECAP_NAND3_G4
XG190 addr_5_ addr_4_ addr_3_ XI2/net026_5_ DECAP_NAND3_G4
XG191 addr_5_ addr_4_ addr_3_ XI2/net026_6_ DECAP_NAND3_G4
XG192 addr_5_ addr_4_ addr_3_ XI2/net026_7_ DECAP_NAND3_G4
XG193 addr_5_ addr_4_ addr__3_ XI2/net026_8_ DECAP_NAND3_G4
XG194 addr_5_ addr_4_ addr__3_ XI2/net026_9_ DECAP_NAND3_G4
XG195 addr_5_ addr_4_ addr__3_ XI2/net026_10_ DECAP_NAND3_G4
XG196 addr_5_ addr_4_ addr__3_ XI2/net026_11_ DECAP_NAND3_G4
XG197 addr_5_ addr_4_ addr__3_ XI2/net026_12_ DECAP_NAND3_G4
XG198 addr_5_ addr_4_ addr__3_ XI2/net026_13_ DECAP_NAND3_G4
XG199 addr_5_ addr_4_ addr__3_ XI2/net026_14_ DECAP_NAND3_G4
XG200 addr_5_ addr_4_ addr__3_ XI2/net026_15_ DECAP_NAND3_G4
XG201 addr_5_ addr__4_ addr_3_ XI2/net026_16_ DECAP_NAND3_G4
XG202 addr_5_ addr__4_ addr_3_ XI2/net026_17_ DECAP_NAND3_G4
XG203 addr_5_ addr__4_ addr_3_ XI2/net026_18_ DECAP_NAND3_G4
XG204 addr_5_ addr__4_ addr_3_ XI2/net026_19_ DECAP_NAND3_G4
XG205 addr_5_ addr__4_ addr_3_ XI2/net026_20_ DECAP_NAND3_G4
XG206 addr_5_ addr__4_ addr_3_ XI2/net026_21_ DECAP_NAND3_G4
XG207 addr_5_ addr__4_ addr_3_ XI2/net026_22_ DECAP_NAND3_G4
XG208 addr_5_ addr__4_ addr_3_ XI2/net026_23_ DECAP_NAND3_G4
XG209 addr_5_ addr__4_ addr__3_ XI2/net026_24_ DECAP_NAND3_G4
XG210 addr_5_ addr__4_ addr__3_ XI2/net026_25_ DECAP_NAND3_G4
XG211 addr_5_ addr__4_ addr__3_ XI2/net026_26_ DECAP_NAND3_G4
XG212 addr_5_ addr__4_ addr__3_ XI2/net026_27_ DECAP_NAND3_G4
XG213 addr_5_ addr__4_ addr__3_ XI2/net026_28_ DECAP_NAND3_G4
XG214 addr_5_ addr__4_ addr__3_ XI2/net026_29_ DECAP_NAND3_G4
XG215 addr_5_ addr__4_ addr__3_ XI2/net026_30_ DECAP_NAND3_G4
XG216 addr_5_ addr__4_ addr__3_ XI2/net026_31_ DECAP_NAND3_G4
XG217 addr__5_ addr_4_ addr_3_ XI2/net026_32_ DECAP_NAND3_G4
XG218 addr__5_ addr_4_ addr_3_ XI2/net026_33_ DECAP_NAND3_G4
XG219 addr__5_ addr_4_ addr_3_ XI2/net026_34_ DECAP_NAND3_G4
XG220 addr__5_ addr_4_ addr_3_ XI2/net026_35_ DECAP_NAND3_G4
XG221 addr__5_ addr_4_ addr_3_ XI2/net026_36_ DECAP_NAND3_G4
XG222 addr__5_ addr_4_ addr_3_ XI2/net026_37_ DECAP_NAND3_G4
XG223 addr__5_ addr_4_ addr_3_ XI2/net026_38_ DECAP_NAND3_G4
XG224 addr__5_ addr_4_ addr_3_ XI2/net026_39_ DECAP_NAND3_G4
XG225 addr__5_ addr_4_ addr__3_ XI2/net026_40_ DECAP_NAND3_G4
XG226 addr__5_ addr_4_ addr__3_ XI2/net026_41_ DECAP_NAND3_G4
XG227 addr__5_ addr_4_ addr__3_ XI2/net026_42_ DECAP_NAND3_G4
XG228 addr__5_ addr_4_ addr__3_ XI2/net026_43_ DECAP_NAND3_G4
XG229 addr__5_ addr_4_ addr__3_ XI2/net026_44_ DECAP_NAND3_G4
XG230 addr__5_ addr_4_ addr__3_ XI2/net026_45_ DECAP_NAND3_G4
XG231 addr__5_ addr_4_ addr__3_ XI2/net026_46_ DECAP_NAND3_G4
XG232 addr__5_ addr_4_ addr__3_ XI2/net026_47_ DECAP_NAND3_G4
XG233 addr__5_ addr__4_ addr_3_ XI2/net026_48_ DECAP_NAND3_G4
XG234 addr__5_ addr__4_ addr_3_ XI2/net026_49_ DECAP_NAND3_G4
XG235 addr__5_ addr__4_ addr_3_ XI2/net026_50_ DECAP_NAND3_G4
XG236 addr__5_ addr__4_ addr_3_ XI2/net026_51_ DECAP_NAND3_G4
XG237 addr__5_ addr__4_ addr_3_ XI2/net026_52_ DECAP_NAND3_G4
XG238 addr__5_ addr__4_ addr_3_ XI2/net026_53_ DECAP_NAND3_G4
XG239 addr__5_ addr__4_ addr_3_ XI2/net026_54_ DECAP_NAND3_G4
XG240 addr__5_ addr__4_ addr_3_ XI2/net026_55_ DECAP_NAND3_G4
XG241 addr__5_ addr__4_ addr__3_ XI2/net026_56_ DECAP_NAND3_G4
XG242 addr__5_ addr__4_ addr__3_ XI2/net026_57_ DECAP_NAND3_G4
XG243 addr__5_ addr__4_ addr__3_ XI2/net026_58_ DECAP_NAND3_G4
XG244 addr__5_ addr__4_ addr__3_ XI2/net026_59_ DECAP_NAND3_G4
XG245 addr__5_ addr__4_ addr__3_ XI2/net026_60_ DECAP_NAND3_G4
XG246 addr__5_ addr__4_ addr__3_ XI2/net026_61_ DECAP_NAND3_G4
XG247 addr__5_ addr__4_ addr__3_ XI2/net026_62_ DECAP_NAND3_G4
XG248 addr__5_ addr__4_ addr__3_ XI2/net026_63_ DECAP_NAND3_G4
XG249 XI6/net018_0_ XI6/net017_0_ XI6/net014_0_ DECAP_NOR2_G3
XG250 XI6/net018_1_ XI6/net017_1_ XI6/net014_1_ DECAP_NOR2_G3
XG251 XI6/net018_2_ XI6/net017_2_ XI6/net014_2_ DECAP_NOR2_G3
XG252 XI6/net018_3_ XI6/net017_3_ XI6/net014_3_ DECAP_NOR2_G3
XG253 XI6/net018_4_ XI6/net017_4_ XI6/net014_4_ DECAP_NOR2_G3
XG254 XI6/net018_5_ XI6/net017_5_ XI6/net014_5_ DECAP_NOR2_G3
XG255 XI6/net018_6_ XI6/net017_6_ XI6/net014_6_ DECAP_NOR2_G3
XG256 XI6/net018_7_ XI6/net017_7_ XI6/net014_7_ DECAP_NOR2_G3
XG257 XI6/net018_8_ XI6/net017_8_ XI6/net014_8_ DECAP_NOR2_G3
XG258 XI6/net018_9_ XI6/net017_9_ XI6/net014_9_ DECAP_NOR2_G3
XG259 XI6/net018_10_ XI6/net017_10_ XI6/net014_10_ DECAP_NOR2_G3
XG260 XI6/net018_11_ XI6/net017_11_ XI6/net014_11_ DECAP_NOR2_G3
XG261 XI6/net018_12_ XI6/net017_12_ XI6/net014_12_ DECAP_NOR2_G3
XG262 XI6/net018_13_ XI6/net017_13_ XI6/net014_13_ DECAP_NOR2_G3
XG263 XI6/net018_14_ XI6/net017_14_ XI6/net014_14_ DECAP_NOR2_G3
XG264 XI6/net018_15_ XI6/net017_15_ XI6/net014_15_ DECAP_NOR2_G5
XG265 addr_7_ addr_6_ XI6/net018_0_ DECAP_NAND2_G6
XG266 addr_7_ XI6/A__6_ XI6/net018_1_ DECAP_NAND2_G6
XG267 addr__7_ addr_6_ XI6/net018_2_ DECAP_NAND2_G6
XG268 addr__7_ XI6/A__6_ XI6/net018_3_ DECAP_NAND2_G6
XG269 addr_7_ addr_6_ XI6/net018_4_ DECAP_NAND2_G6
XG270 addr_7_ XI6/A__6_ XI6/net018_5_ DECAP_NAND2_G6
XG271 addr__7_ addr_6_ XI6/net018_6_ DECAP_NAND2_G6
XG272 addr__7_ XI6/A__6_ XI6/net018_7_ DECAP_NAND2_G6
XG273 addr_7_ addr_6_ XI6/net018_8_ DECAP_NAND2_G6
XG274 addr_7_ XI6/A__6_ XI6/net018_9_ DECAP_NAND2_G6
XG275 addr__7_ addr_6_ XI6/net018_10_ DECAP_NAND2_G6
XG276 addr__7_ XI6/A__6_ XI6/net018_11_ DECAP_NAND2_G6
XG277 addr_7_ addr_6_ XI6/net018_12_ DECAP_NAND2_G6
XG278 addr_7_ XI6/A__6_ XI6/net018_13_ DECAP_NAND2_G6
XG279 addr__7_ addr_6_ XI6/net018_14_ DECAP_NAND2_G6
XG280 addr__7_ XI6/A__6_ XI6/net018_15_ DECAP_NAND2_G6
XG281 addr_9_ addr_8_ XI6/net017_0_ DECAP_NAND2_G6
XG282 addr_9_ addr_8_ XI6/net017_1_ DECAP_NAND2_G6
XG283 addr_9_ addr_8_ XI6/net017_2_ DECAP_NAND2_G6
XG284 addr_9_ addr_8_ XI6/net017_3_ DECAP_NAND2_G6
XG285 addr_9_ addr__8_ XI6/net017_4_ DECAP_NAND2_G6
XG286 addr_9_ addr__8_ XI6/net017_5_ DECAP_NAND2_G6
XG287 addr_9_ addr__8_ XI6/net017_6_ DECAP_NAND2_G6
XG288 addr_9_ addr__8_ XI6/net017_7_ DECAP_NAND2_G6
XG289 addr__9_ addr_8_ XI6/net017_8_ DECAP_NAND2_G6
XG290 addr__9_ addr_8_ XI6/net017_9_ DECAP_NAND2_G6
XG291 addr__9_ addr_8_ XI6/net017_10_ DECAP_NAND2_G6
XG292 addr__9_ addr_8_ XI6/net017_11_ DECAP_NAND2_G6
XG293 addr__9_ addr__8_ XI6/net017_12_ DECAP_NAND2_G6
XG294 addr__9_ addr__8_ XI6/net017_13_ DECAP_NAND2_G6
XG295 addr__9_ addr__8_ XI6/net017_14_ DECAP_NAND2_G6
XG296 addr__9_ addr__8_ XI6/net017_15_ DECAP_NAND2_G6
XG297 XI11_7/XI3/net17 XI11_7/XI3/net5 DECAP_INV_G7
XG298 XI11_7/XI3/net5 XI11_7/preck DECAP_INV_G8
XG299 sck_bar XI11_7/XI3/net018 DECAP_INV_G9
XG300 XI11_7/XI3/net018 XI11_7/XI3/net012 DECAP_INV_G9
XG301 XI11_7/XI3/net014 XI11_7/XI3/net7 DECAP_INV_G9
XG302 XI11_7/XI3/net012 XI11_7/XI3/net014 DECAP_INV_G9
XG303 XI11_7/XI4/net063 XI11_7/XI4/net0112 DECAP_INV_G10
XG304 XI11_7/XI4/net26 XI11_7/XI4/net089 DECAP_INV_G10
XG305 XI11_7/XI4/data_out XI11_7/XI4/data_out_ DECAP_INV_G10
XG306 XI11_7/XI4/net20 XI11_7/XI4/net0103 DECAP_INV_G10
XG307 XI11_7/net12 XI11_7/XI4/net32 DECAP_INV_G7
XG308 XI11_7/net9 XI11_7/XI4/net52 DECAP_INV_G7
XG309 XI11_7/XI4/data_out_ XI11_7/XI4/data_out DECAP_INV_G10
XG310 XI11_7/XI0/XI0_63/d__15_ XI11_7/XI0/XI0_63/d_15_ DECAP_INV_G11
XG311 XI11_7/XI0/XI0_63/d__14_ XI11_7/XI0/XI0_63/d_14_ DECAP_INV_G11
XG312 XI11_7/XI0/XI0_63/d__13_ XI11_7/XI0/XI0_63/d_13_ DECAP_INV_G11
XG313 XI11_7/XI0/XI0_63/d__12_ XI11_7/XI0/XI0_63/d_12_ DECAP_INV_G11
XG314 XI11_7/XI0/XI0_63/d__11_ XI11_7/XI0/XI0_63/d_11_ DECAP_INV_G11
XG315 XI11_7/XI0/XI0_63/d__10_ XI11_7/XI0/XI0_63/d_10_ DECAP_INV_G11
XG316 XI11_7/XI0/XI0_63/d__9_ XI11_7/XI0/XI0_63/d_9_ DECAP_INV_G11
XG317 XI11_7/XI0/XI0_63/d__8_ XI11_7/XI0/XI0_63/d_8_ DECAP_INV_G11
XG318 XI11_7/XI0/XI0_63/d__7_ XI11_7/XI0/XI0_63/d_7_ DECAP_INV_G11
XG319 XI11_7/XI0/XI0_63/d__6_ XI11_7/XI0/XI0_63/d_6_ DECAP_INV_G11
XG320 XI11_7/XI0/XI0_63/d__5_ XI11_7/XI0/XI0_63/d_5_ DECAP_INV_G11
XG321 XI11_7/XI0/XI0_63/d__4_ XI11_7/XI0/XI0_63/d_4_ DECAP_INV_G11
XG322 XI11_7/XI0/XI0_63/d__3_ XI11_7/XI0/XI0_63/d_3_ DECAP_INV_G11
XG323 XI11_7/XI0/XI0_63/d__2_ XI11_7/XI0/XI0_63/d_2_ DECAP_INV_G11
XG324 XI11_7/XI0/XI0_63/d__1_ XI11_7/XI0/XI0_63/d_1_ DECAP_INV_G11
XG325 XI11_7/XI0/XI0_63/d__0_ XI11_7/XI0/XI0_63/d_0_ DECAP_INV_G11
XG326 XI11_7/XI0/XI0_63/d_15_ XI11_7/XI0/XI0_63/d__15_ DECAP_INV_G11
XG327 XI11_7/XI0/XI0_63/d_14_ XI11_7/XI0/XI0_63/d__14_ DECAP_INV_G11
XG328 XI11_7/XI0/XI0_63/d_13_ XI11_7/XI0/XI0_63/d__13_ DECAP_INV_G11
XG329 XI11_7/XI0/XI0_63/d_12_ XI11_7/XI0/XI0_63/d__12_ DECAP_INV_G11
XG330 XI11_7/XI0/XI0_63/d_11_ XI11_7/XI0/XI0_63/d__11_ DECAP_INV_G11
XG331 XI11_7/XI0/XI0_63/d_10_ XI11_7/XI0/XI0_63/d__10_ DECAP_INV_G11
XG332 XI11_7/XI0/XI0_63/d_9_ XI11_7/XI0/XI0_63/d__9_ DECAP_INV_G11
XG333 XI11_7/XI0/XI0_63/d_8_ XI11_7/XI0/XI0_63/d__8_ DECAP_INV_G11
XG334 XI11_7/XI0/XI0_63/d_7_ XI11_7/XI0/XI0_63/d__7_ DECAP_INV_G11
XG335 XI11_7/XI0/XI0_63/d_6_ XI11_7/XI0/XI0_63/d__6_ DECAP_INV_G11
XG336 XI11_7/XI0/XI0_63/d_5_ XI11_7/XI0/XI0_63/d__5_ DECAP_INV_G11
XG337 XI11_7/XI0/XI0_63/d_4_ XI11_7/XI0/XI0_63/d__4_ DECAP_INV_G11
XG338 XI11_7/XI0/XI0_63/d_3_ XI11_7/XI0/XI0_63/d__3_ DECAP_INV_G11
XG339 XI11_7/XI0/XI0_63/d_2_ XI11_7/XI0/XI0_63/d__2_ DECAP_INV_G11
XG340 XI11_7/XI0/XI0_63/d_1_ XI11_7/XI0/XI0_63/d__1_ DECAP_INV_G11
XG341 XI11_7/XI0/XI0_63/d_0_ XI11_7/XI0/XI0_63/d__0_ DECAP_INV_G11
XG342 XI11_7/XI0/XI0_62/d__15_ XI11_7/XI0/XI0_62/d_15_ DECAP_INV_G11
XG343 XI11_7/XI0/XI0_62/d__14_ XI11_7/XI0/XI0_62/d_14_ DECAP_INV_G11
XG344 XI11_7/XI0/XI0_62/d__13_ XI11_7/XI0/XI0_62/d_13_ DECAP_INV_G11
XG345 XI11_7/XI0/XI0_62/d__12_ XI11_7/XI0/XI0_62/d_12_ DECAP_INV_G11
XG346 XI11_7/XI0/XI0_62/d__11_ XI11_7/XI0/XI0_62/d_11_ DECAP_INV_G11
XG347 XI11_7/XI0/XI0_62/d__10_ XI11_7/XI0/XI0_62/d_10_ DECAP_INV_G11
XG348 XI11_7/XI0/XI0_62/d__9_ XI11_7/XI0/XI0_62/d_9_ DECAP_INV_G11
XG349 XI11_7/XI0/XI0_62/d__8_ XI11_7/XI0/XI0_62/d_8_ DECAP_INV_G11
XG350 XI11_7/XI0/XI0_62/d__7_ XI11_7/XI0/XI0_62/d_7_ DECAP_INV_G11
XG351 XI11_7/XI0/XI0_62/d__6_ XI11_7/XI0/XI0_62/d_6_ DECAP_INV_G11
XG352 XI11_7/XI0/XI0_62/d__5_ XI11_7/XI0/XI0_62/d_5_ DECAP_INV_G11
XG353 XI11_7/XI0/XI0_62/d__4_ XI11_7/XI0/XI0_62/d_4_ DECAP_INV_G11
XG354 XI11_7/XI0/XI0_62/d__3_ XI11_7/XI0/XI0_62/d_3_ DECAP_INV_G11
XG355 XI11_7/XI0/XI0_62/d__2_ XI11_7/XI0/XI0_62/d_2_ DECAP_INV_G11
XG356 XI11_7/XI0/XI0_62/d__1_ XI11_7/XI0/XI0_62/d_1_ DECAP_INV_G11
XG357 XI11_7/XI0/XI0_62/d__0_ XI11_7/XI0/XI0_62/d_0_ DECAP_INV_G11
XG358 XI11_7/XI0/XI0_62/d_15_ XI11_7/XI0/XI0_62/d__15_ DECAP_INV_G11
XG359 XI11_7/XI0/XI0_62/d_14_ XI11_7/XI0/XI0_62/d__14_ DECAP_INV_G11
XG360 XI11_7/XI0/XI0_62/d_13_ XI11_7/XI0/XI0_62/d__13_ DECAP_INV_G11
XG361 XI11_7/XI0/XI0_62/d_12_ XI11_7/XI0/XI0_62/d__12_ DECAP_INV_G11
XG362 XI11_7/XI0/XI0_62/d_11_ XI11_7/XI0/XI0_62/d__11_ DECAP_INV_G11
XG363 XI11_7/XI0/XI0_62/d_10_ XI11_7/XI0/XI0_62/d__10_ DECAP_INV_G11
XG364 XI11_7/XI0/XI0_62/d_9_ XI11_7/XI0/XI0_62/d__9_ DECAP_INV_G11
XG365 XI11_7/XI0/XI0_62/d_8_ XI11_7/XI0/XI0_62/d__8_ DECAP_INV_G11
XG366 XI11_7/XI0/XI0_62/d_7_ XI11_7/XI0/XI0_62/d__7_ DECAP_INV_G11
XG367 XI11_7/XI0/XI0_62/d_6_ XI11_7/XI0/XI0_62/d__6_ DECAP_INV_G11
XG368 XI11_7/XI0/XI0_62/d_5_ XI11_7/XI0/XI0_62/d__5_ DECAP_INV_G11
XG369 XI11_7/XI0/XI0_62/d_4_ XI11_7/XI0/XI0_62/d__4_ DECAP_INV_G11
XG370 XI11_7/XI0/XI0_62/d_3_ XI11_7/XI0/XI0_62/d__3_ DECAP_INV_G11
XG371 XI11_7/XI0/XI0_62/d_2_ XI11_7/XI0/XI0_62/d__2_ DECAP_INV_G11
XG372 XI11_7/XI0/XI0_62/d_1_ XI11_7/XI0/XI0_62/d__1_ DECAP_INV_G11
XG373 XI11_7/XI0/XI0_62/d_0_ XI11_7/XI0/XI0_62/d__0_ DECAP_INV_G11
XG374 XI11_7/XI0/XI0_61/d__15_ XI11_7/XI0/XI0_61/d_15_ DECAP_INV_G11
XG375 XI11_7/XI0/XI0_61/d__14_ XI11_7/XI0/XI0_61/d_14_ DECAP_INV_G11
XG376 XI11_7/XI0/XI0_61/d__13_ XI11_7/XI0/XI0_61/d_13_ DECAP_INV_G11
XG377 XI11_7/XI0/XI0_61/d__12_ XI11_7/XI0/XI0_61/d_12_ DECAP_INV_G11
XG378 XI11_7/XI0/XI0_61/d__11_ XI11_7/XI0/XI0_61/d_11_ DECAP_INV_G11
XG379 XI11_7/XI0/XI0_61/d__10_ XI11_7/XI0/XI0_61/d_10_ DECAP_INV_G11
XG380 XI11_7/XI0/XI0_61/d__9_ XI11_7/XI0/XI0_61/d_9_ DECAP_INV_G11
XG381 XI11_7/XI0/XI0_61/d__8_ XI11_7/XI0/XI0_61/d_8_ DECAP_INV_G11
XG382 XI11_7/XI0/XI0_61/d__7_ XI11_7/XI0/XI0_61/d_7_ DECAP_INV_G11
XG383 XI11_7/XI0/XI0_61/d__6_ XI11_7/XI0/XI0_61/d_6_ DECAP_INV_G11
XG384 XI11_7/XI0/XI0_61/d__5_ XI11_7/XI0/XI0_61/d_5_ DECAP_INV_G11
XG385 XI11_7/XI0/XI0_61/d__4_ XI11_7/XI0/XI0_61/d_4_ DECAP_INV_G11
XG386 XI11_7/XI0/XI0_61/d__3_ XI11_7/XI0/XI0_61/d_3_ DECAP_INV_G11
XG387 XI11_7/XI0/XI0_61/d__2_ XI11_7/XI0/XI0_61/d_2_ DECAP_INV_G11
XG388 XI11_7/XI0/XI0_61/d__1_ XI11_7/XI0/XI0_61/d_1_ DECAP_INV_G11
XG389 XI11_7/XI0/XI0_61/d__0_ XI11_7/XI0/XI0_61/d_0_ DECAP_INV_G11
XG390 XI11_7/XI0/XI0_61/d_15_ XI11_7/XI0/XI0_61/d__15_ DECAP_INV_G11
XG391 XI11_7/XI0/XI0_61/d_14_ XI11_7/XI0/XI0_61/d__14_ DECAP_INV_G11
XG392 XI11_7/XI0/XI0_61/d_13_ XI11_7/XI0/XI0_61/d__13_ DECAP_INV_G11
XG393 XI11_7/XI0/XI0_61/d_12_ XI11_7/XI0/XI0_61/d__12_ DECAP_INV_G11
XG394 XI11_7/XI0/XI0_61/d_11_ XI11_7/XI0/XI0_61/d__11_ DECAP_INV_G11
XG395 XI11_7/XI0/XI0_61/d_10_ XI11_7/XI0/XI0_61/d__10_ DECAP_INV_G11
XG396 XI11_7/XI0/XI0_61/d_9_ XI11_7/XI0/XI0_61/d__9_ DECAP_INV_G11
XG397 XI11_7/XI0/XI0_61/d_8_ XI11_7/XI0/XI0_61/d__8_ DECAP_INV_G11
XG398 XI11_7/XI0/XI0_61/d_7_ XI11_7/XI0/XI0_61/d__7_ DECAP_INV_G11
XG399 XI11_7/XI0/XI0_61/d_6_ XI11_7/XI0/XI0_61/d__6_ DECAP_INV_G11
XG400 XI11_7/XI0/XI0_61/d_5_ XI11_7/XI0/XI0_61/d__5_ DECAP_INV_G11
XG401 XI11_7/XI0/XI0_61/d_4_ XI11_7/XI0/XI0_61/d__4_ DECAP_INV_G11
XG402 XI11_7/XI0/XI0_61/d_3_ XI11_7/XI0/XI0_61/d__3_ DECAP_INV_G11
XG403 XI11_7/XI0/XI0_61/d_2_ XI11_7/XI0/XI0_61/d__2_ DECAP_INV_G11
XG404 XI11_7/XI0/XI0_61/d_1_ XI11_7/XI0/XI0_61/d__1_ DECAP_INV_G11
XG405 XI11_7/XI0/XI0_61/d_0_ XI11_7/XI0/XI0_61/d__0_ DECAP_INV_G11
XG406 XI11_7/XI0/XI0_60/d__15_ XI11_7/XI0/XI0_60/d_15_ DECAP_INV_G11
XG407 XI11_7/XI0/XI0_60/d__14_ XI11_7/XI0/XI0_60/d_14_ DECAP_INV_G11
XG408 XI11_7/XI0/XI0_60/d__13_ XI11_7/XI0/XI0_60/d_13_ DECAP_INV_G11
XG409 XI11_7/XI0/XI0_60/d__12_ XI11_7/XI0/XI0_60/d_12_ DECAP_INV_G11
XG410 XI11_7/XI0/XI0_60/d__11_ XI11_7/XI0/XI0_60/d_11_ DECAP_INV_G11
XG411 XI11_7/XI0/XI0_60/d__10_ XI11_7/XI0/XI0_60/d_10_ DECAP_INV_G11
XG412 XI11_7/XI0/XI0_60/d__9_ XI11_7/XI0/XI0_60/d_9_ DECAP_INV_G11
XG413 XI11_7/XI0/XI0_60/d__8_ XI11_7/XI0/XI0_60/d_8_ DECAP_INV_G11
XG414 XI11_7/XI0/XI0_60/d__7_ XI11_7/XI0/XI0_60/d_7_ DECAP_INV_G11
XG415 XI11_7/XI0/XI0_60/d__6_ XI11_7/XI0/XI0_60/d_6_ DECAP_INV_G11
XG416 XI11_7/XI0/XI0_60/d__5_ XI11_7/XI0/XI0_60/d_5_ DECAP_INV_G11
XG417 XI11_7/XI0/XI0_60/d__4_ XI11_7/XI0/XI0_60/d_4_ DECAP_INV_G11
XG418 XI11_7/XI0/XI0_60/d__3_ XI11_7/XI0/XI0_60/d_3_ DECAP_INV_G11
XG419 XI11_7/XI0/XI0_60/d__2_ XI11_7/XI0/XI0_60/d_2_ DECAP_INV_G11
XG420 XI11_7/XI0/XI0_60/d__1_ XI11_7/XI0/XI0_60/d_1_ DECAP_INV_G11
XG421 XI11_7/XI0/XI0_60/d__0_ XI11_7/XI0/XI0_60/d_0_ DECAP_INV_G11
XG422 XI11_7/XI0/XI0_60/d_15_ XI11_7/XI0/XI0_60/d__15_ DECAP_INV_G11
XG423 XI11_7/XI0/XI0_60/d_14_ XI11_7/XI0/XI0_60/d__14_ DECAP_INV_G11
XG424 XI11_7/XI0/XI0_60/d_13_ XI11_7/XI0/XI0_60/d__13_ DECAP_INV_G11
XG425 XI11_7/XI0/XI0_60/d_12_ XI11_7/XI0/XI0_60/d__12_ DECAP_INV_G11
XG426 XI11_7/XI0/XI0_60/d_11_ XI11_7/XI0/XI0_60/d__11_ DECAP_INV_G11
XG427 XI11_7/XI0/XI0_60/d_10_ XI11_7/XI0/XI0_60/d__10_ DECAP_INV_G11
XG428 XI11_7/XI0/XI0_60/d_9_ XI11_7/XI0/XI0_60/d__9_ DECAP_INV_G11
XG429 XI11_7/XI0/XI0_60/d_8_ XI11_7/XI0/XI0_60/d__8_ DECAP_INV_G11
XG430 XI11_7/XI0/XI0_60/d_7_ XI11_7/XI0/XI0_60/d__7_ DECAP_INV_G11
XG431 XI11_7/XI0/XI0_60/d_6_ XI11_7/XI0/XI0_60/d__6_ DECAP_INV_G11
XG432 XI11_7/XI0/XI0_60/d_5_ XI11_7/XI0/XI0_60/d__5_ DECAP_INV_G11
XG433 XI11_7/XI0/XI0_60/d_4_ XI11_7/XI0/XI0_60/d__4_ DECAP_INV_G11
XG434 XI11_7/XI0/XI0_60/d_3_ XI11_7/XI0/XI0_60/d__3_ DECAP_INV_G11
XG435 XI11_7/XI0/XI0_60/d_2_ XI11_7/XI0/XI0_60/d__2_ DECAP_INV_G11
XG436 XI11_7/XI0/XI0_60/d_1_ XI11_7/XI0/XI0_60/d__1_ DECAP_INV_G11
XG437 XI11_7/XI0/XI0_60/d_0_ XI11_7/XI0/XI0_60/d__0_ DECAP_INV_G11
XG438 XI11_7/XI0/XI0_59/d__15_ XI11_7/XI0/XI0_59/d_15_ DECAP_INV_G11
XG439 XI11_7/XI0/XI0_59/d__14_ XI11_7/XI0/XI0_59/d_14_ DECAP_INV_G11
XG440 XI11_7/XI0/XI0_59/d__13_ XI11_7/XI0/XI0_59/d_13_ DECAP_INV_G11
XG441 XI11_7/XI0/XI0_59/d__12_ XI11_7/XI0/XI0_59/d_12_ DECAP_INV_G11
XG442 XI11_7/XI0/XI0_59/d__11_ XI11_7/XI0/XI0_59/d_11_ DECAP_INV_G11
XG443 XI11_7/XI0/XI0_59/d__10_ XI11_7/XI0/XI0_59/d_10_ DECAP_INV_G11
XG444 XI11_7/XI0/XI0_59/d__9_ XI11_7/XI0/XI0_59/d_9_ DECAP_INV_G11
XG445 XI11_7/XI0/XI0_59/d__8_ XI11_7/XI0/XI0_59/d_8_ DECAP_INV_G11
XG446 XI11_7/XI0/XI0_59/d__7_ XI11_7/XI0/XI0_59/d_7_ DECAP_INV_G11
XG447 XI11_7/XI0/XI0_59/d__6_ XI11_7/XI0/XI0_59/d_6_ DECAP_INV_G11
XG448 XI11_7/XI0/XI0_59/d__5_ XI11_7/XI0/XI0_59/d_5_ DECAP_INV_G11
XG449 XI11_7/XI0/XI0_59/d__4_ XI11_7/XI0/XI0_59/d_4_ DECAP_INV_G11
XG450 XI11_7/XI0/XI0_59/d__3_ XI11_7/XI0/XI0_59/d_3_ DECAP_INV_G11
XG451 XI11_7/XI0/XI0_59/d__2_ XI11_7/XI0/XI0_59/d_2_ DECAP_INV_G11
XG452 XI11_7/XI0/XI0_59/d__1_ XI11_7/XI0/XI0_59/d_1_ DECAP_INV_G11
XG453 XI11_7/XI0/XI0_59/d__0_ XI11_7/XI0/XI0_59/d_0_ DECAP_INV_G11
XG454 XI11_7/XI0/XI0_59/d_15_ XI11_7/XI0/XI0_59/d__15_ DECAP_INV_G11
XG455 XI11_7/XI0/XI0_59/d_14_ XI11_7/XI0/XI0_59/d__14_ DECAP_INV_G11
XG456 XI11_7/XI0/XI0_59/d_13_ XI11_7/XI0/XI0_59/d__13_ DECAP_INV_G11
XG457 XI11_7/XI0/XI0_59/d_12_ XI11_7/XI0/XI0_59/d__12_ DECAP_INV_G11
XG458 XI11_7/XI0/XI0_59/d_11_ XI11_7/XI0/XI0_59/d__11_ DECAP_INV_G11
XG459 XI11_7/XI0/XI0_59/d_10_ XI11_7/XI0/XI0_59/d__10_ DECAP_INV_G11
XG460 XI11_7/XI0/XI0_59/d_9_ XI11_7/XI0/XI0_59/d__9_ DECAP_INV_G11
XG461 XI11_7/XI0/XI0_59/d_8_ XI11_7/XI0/XI0_59/d__8_ DECAP_INV_G11
XG462 XI11_7/XI0/XI0_59/d_7_ XI11_7/XI0/XI0_59/d__7_ DECAP_INV_G11
XG463 XI11_7/XI0/XI0_59/d_6_ XI11_7/XI0/XI0_59/d__6_ DECAP_INV_G11
XG464 XI11_7/XI0/XI0_59/d_5_ XI11_7/XI0/XI0_59/d__5_ DECAP_INV_G11
XG465 XI11_7/XI0/XI0_59/d_4_ XI11_7/XI0/XI0_59/d__4_ DECAP_INV_G11
XG466 XI11_7/XI0/XI0_59/d_3_ XI11_7/XI0/XI0_59/d__3_ DECAP_INV_G11
XG467 XI11_7/XI0/XI0_59/d_2_ XI11_7/XI0/XI0_59/d__2_ DECAP_INV_G11
XG468 XI11_7/XI0/XI0_59/d_1_ XI11_7/XI0/XI0_59/d__1_ DECAP_INV_G11
XG469 XI11_7/XI0/XI0_59/d_0_ XI11_7/XI0/XI0_59/d__0_ DECAP_INV_G11
XG470 XI11_7/XI0/XI0_58/d__15_ XI11_7/XI0/XI0_58/d_15_ DECAP_INV_G11
XG471 XI11_7/XI0/XI0_58/d__14_ XI11_7/XI0/XI0_58/d_14_ DECAP_INV_G11
XG472 XI11_7/XI0/XI0_58/d__13_ XI11_7/XI0/XI0_58/d_13_ DECAP_INV_G11
XG473 XI11_7/XI0/XI0_58/d__12_ XI11_7/XI0/XI0_58/d_12_ DECAP_INV_G11
XG474 XI11_7/XI0/XI0_58/d__11_ XI11_7/XI0/XI0_58/d_11_ DECAP_INV_G11
XG475 XI11_7/XI0/XI0_58/d__10_ XI11_7/XI0/XI0_58/d_10_ DECAP_INV_G11
XG476 XI11_7/XI0/XI0_58/d__9_ XI11_7/XI0/XI0_58/d_9_ DECAP_INV_G11
XG477 XI11_7/XI0/XI0_58/d__8_ XI11_7/XI0/XI0_58/d_8_ DECAP_INV_G11
XG478 XI11_7/XI0/XI0_58/d__7_ XI11_7/XI0/XI0_58/d_7_ DECAP_INV_G11
XG479 XI11_7/XI0/XI0_58/d__6_ XI11_7/XI0/XI0_58/d_6_ DECAP_INV_G11
XG480 XI11_7/XI0/XI0_58/d__5_ XI11_7/XI0/XI0_58/d_5_ DECAP_INV_G11
XG481 XI11_7/XI0/XI0_58/d__4_ XI11_7/XI0/XI0_58/d_4_ DECAP_INV_G11
XG482 XI11_7/XI0/XI0_58/d__3_ XI11_7/XI0/XI0_58/d_3_ DECAP_INV_G11
XG483 XI11_7/XI0/XI0_58/d__2_ XI11_7/XI0/XI0_58/d_2_ DECAP_INV_G11
XG484 XI11_7/XI0/XI0_58/d__1_ XI11_7/XI0/XI0_58/d_1_ DECAP_INV_G11
XG485 XI11_7/XI0/XI0_58/d__0_ XI11_7/XI0/XI0_58/d_0_ DECAP_INV_G11
XG486 XI11_7/XI0/XI0_58/d_15_ XI11_7/XI0/XI0_58/d__15_ DECAP_INV_G11
XG487 XI11_7/XI0/XI0_58/d_14_ XI11_7/XI0/XI0_58/d__14_ DECAP_INV_G11
XG488 XI11_7/XI0/XI0_58/d_13_ XI11_7/XI0/XI0_58/d__13_ DECAP_INV_G11
XG489 XI11_7/XI0/XI0_58/d_12_ XI11_7/XI0/XI0_58/d__12_ DECAP_INV_G11
XG490 XI11_7/XI0/XI0_58/d_11_ XI11_7/XI0/XI0_58/d__11_ DECAP_INV_G11
XG491 XI11_7/XI0/XI0_58/d_10_ XI11_7/XI0/XI0_58/d__10_ DECAP_INV_G11
XG492 XI11_7/XI0/XI0_58/d_9_ XI11_7/XI0/XI0_58/d__9_ DECAP_INV_G11
XG493 XI11_7/XI0/XI0_58/d_8_ XI11_7/XI0/XI0_58/d__8_ DECAP_INV_G11
XG494 XI11_7/XI0/XI0_58/d_7_ XI11_7/XI0/XI0_58/d__7_ DECAP_INV_G11
XG495 XI11_7/XI0/XI0_58/d_6_ XI11_7/XI0/XI0_58/d__6_ DECAP_INV_G11
XG496 XI11_7/XI0/XI0_58/d_5_ XI11_7/XI0/XI0_58/d__5_ DECAP_INV_G11
XG497 XI11_7/XI0/XI0_58/d_4_ XI11_7/XI0/XI0_58/d__4_ DECAP_INV_G11
XG498 XI11_7/XI0/XI0_58/d_3_ XI11_7/XI0/XI0_58/d__3_ DECAP_INV_G11
XG499 XI11_7/XI0/XI0_58/d_2_ XI11_7/XI0/XI0_58/d__2_ DECAP_INV_G11
XG500 XI11_7/XI0/XI0_58/d_1_ XI11_7/XI0/XI0_58/d__1_ DECAP_INV_G11
XG501 XI11_7/XI0/XI0_58/d_0_ XI11_7/XI0/XI0_58/d__0_ DECAP_INV_G11
XG502 XI11_7/XI0/XI0_57/d__15_ XI11_7/XI0/XI0_57/d_15_ DECAP_INV_G11
XG503 XI11_7/XI0/XI0_57/d__14_ XI11_7/XI0/XI0_57/d_14_ DECAP_INV_G11
XG504 XI11_7/XI0/XI0_57/d__13_ XI11_7/XI0/XI0_57/d_13_ DECAP_INV_G11
XG505 XI11_7/XI0/XI0_57/d__12_ XI11_7/XI0/XI0_57/d_12_ DECAP_INV_G11
XG506 XI11_7/XI0/XI0_57/d__11_ XI11_7/XI0/XI0_57/d_11_ DECAP_INV_G11
XG507 XI11_7/XI0/XI0_57/d__10_ XI11_7/XI0/XI0_57/d_10_ DECAP_INV_G11
XG508 XI11_7/XI0/XI0_57/d__9_ XI11_7/XI0/XI0_57/d_9_ DECAP_INV_G11
XG509 XI11_7/XI0/XI0_57/d__8_ XI11_7/XI0/XI0_57/d_8_ DECAP_INV_G11
XG510 XI11_7/XI0/XI0_57/d__7_ XI11_7/XI0/XI0_57/d_7_ DECAP_INV_G11
XG511 XI11_7/XI0/XI0_57/d__6_ XI11_7/XI0/XI0_57/d_6_ DECAP_INV_G11
XG512 XI11_7/XI0/XI0_57/d__5_ XI11_7/XI0/XI0_57/d_5_ DECAP_INV_G11
XG513 XI11_7/XI0/XI0_57/d__4_ XI11_7/XI0/XI0_57/d_4_ DECAP_INV_G11
XG514 XI11_7/XI0/XI0_57/d__3_ XI11_7/XI0/XI0_57/d_3_ DECAP_INV_G11
XG515 XI11_7/XI0/XI0_57/d__2_ XI11_7/XI0/XI0_57/d_2_ DECAP_INV_G11
XG516 XI11_7/XI0/XI0_57/d__1_ XI11_7/XI0/XI0_57/d_1_ DECAP_INV_G11
XG517 XI11_7/XI0/XI0_57/d__0_ XI11_7/XI0/XI0_57/d_0_ DECAP_INV_G11
XG518 XI11_7/XI0/XI0_57/d_15_ XI11_7/XI0/XI0_57/d__15_ DECAP_INV_G11
XG519 XI11_7/XI0/XI0_57/d_14_ XI11_7/XI0/XI0_57/d__14_ DECAP_INV_G11
XG520 XI11_7/XI0/XI0_57/d_13_ XI11_7/XI0/XI0_57/d__13_ DECAP_INV_G11
XG521 XI11_7/XI0/XI0_57/d_12_ XI11_7/XI0/XI0_57/d__12_ DECAP_INV_G11
XG522 XI11_7/XI0/XI0_57/d_11_ XI11_7/XI0/XI0_57/d__11_ DECAP_INV_G11
XG523 XI11_7/XI0/XI0_57/d_10_ XI11_7/XI0/XI0_57/d__10_ DECAP_INV_G11
XG524 XI11_7/XI0/XI0_57/d_9_ XI11_7/XI0/XI0_57/d__9_ DECAP_INV_G11
XG525 XI11_7/XI0/XI0_57/d_8_ XI11_7/XI0/XI0_57/d__8_ DECAP_INV_G11
XG526 XI11_7/XI0/XI0_57/d_7_ XI11_7/XI0/XI0_57/d__7_ DECAP_INV_G11
XG527 XI11_7/XI0/XI0_57/d_6_ XI11_7/XI0/XI0_57/d__6_ DECAP_INV_G11
XG528 XI11_7/XI0/XI0_57/d_5_ XI11_7/XI0/XI0_57/d__5_ DECAP_INV_G11
XG529 XI11_7/XI0/XI0_57/d_4_ XI11_7/XI0/XI0_57/d__4_ DECAP_INV_G11
XG530 XI11_7/XI0/XI0_57/d_3_ XI11_7/XI0/XI0_57/d__3_ DECAP_INV_G11
XG531 XI11_7/XI0/XI0_57/d_2_ XI11_7/XI0/XI0_57/d__2_ DECAP_INV_G11
XG532 XI11_7/XI0/XI0_57/d_1_ XI11_7/XI0/XI0_57/d__1_ DECAP_INV_G11
XG533 XI11_7/XI0/XI0_57/d_0_ XI11_7/XI0/XI0_57/d__0_ DECAP_INV_G11
XG534 XI11_7/XI0/XI0_56/d__15_ XI11_7/XI0/XI0_56/d_15_ DECAP_INV_G11
XG535 XI11_7/XI0/XI0_56/d__14_ XI11_7/XI0/XI0_56/d_14_ DECAP_INV_G11
XG536 XI11_7/XI0/XI0_56/d__13_ XI11_7/XI0/XI0_56/d_13_ DECAP_INV_G11
XG537 XI11_7/XI0/XI0_56/d__12_ XI11_7/XI0/XI0_56/d_12_ DECAP_INV_G11
XG538 XI11_7/XI0/XI0_56/d__11_ XI11_7/XI0/XI0_56/d_11_ DECAP_INV_G11
XG539 XI11_7/XI0/XI0_56/d__10_ XI11_7/XI0/XI0_56/d_10_ DECAP_INV_G11
XG540 XI11_7/XI0/XI0_56/d__9_ XI11_7/XI0/XI0_56/d_9_ DECAP_INV_G11
XG541 XI11_7/XI0/XI0_56/d__8_ XI11_7/XI0/XI0_56/d_8_ DECAP_INV_G11
XG542 XI11_7/XI0/XI0_56/d__7_ XI11_7/XI0/XI0_56/d_7_ DECAP_INV_G11
XG543 XI11_7/XI0/XI0_56/d__6_ XI11_7/XI0/XI0_56/d_6_ DECAP_INV_G11
XG544 XI11_7/XI0/XI0_56/d__5_ XI11_7/XI0/XI0_56/d_5_ DECAP_INV_G11
XG545 XI11_7/XI0/XI0_56/d__4_ XI11_7/XI0/XI0_56/d_4_ DECAP_INV_G11
XG546 XI11_7/XI0/XI0_56/d__3_ XI11_7/XI0/XI0_56/d_3_ DECAP_INV_G11
XG547 XI11_7/XI0/XI0_56/d__2_ XI11_7/XI0/XI0_56/d_2_ DECAP_INV_G11
XG548 XI11_7/XI0/XI0_56/d__1_ XI11_7/XI0/XI0_56/d_1_ DECAP_INV_G11
XG549 XI11_7/XI0/XI0_56/d__0_ XI11_7/XI0/XI0_56/d_0_ DECAP_INV_G11
XG550 XI11_7/XI0/XI0_56/d_15_ XI11_7/XI0/XI0_56/d__15_ DECAP_INV_G11
XG551 XI11_7/XI0/XI0_56/d_14_ XI11_7/XI0/XI0_56/d__14_ DECAP_INV_G11
XG552 XI11_7/XI0/XI0_56/d_13_ XI11_7/XI0/XI0_56/d__13_ DECAP_INV_G11
XG553 XI11_7/XI0/XI0_56/d_12_ XI11_7/XI0/XI0_56/d__12_ DECAP_INV_G11
XG554 XI11_7/XI0/XI0_56/d_11_ XI11_7/XI0/XI0_56/d__11_ DECAP_INV_G11
XG555 XI11_7/XI0/XI0_56/d_10_ XI11_7/XI0/XI0_56/d__10_ DECAP_INV_G11
XG556 XI11_7/XI0/XI0_56/d_9_ XI11_7/XI0/XI0_56/d__9_ DECAP_INV_G11
XG557 XI11_7/XI0/XI0_56/d_8_ XI11_7/XI0/XI0_56/d__8_ DECAP_INV_G11
XG558 XI11_7/XI0/XI0_56/d_7_ XI11_7/XI0/XI0_56/d__7_ DECAP_INV_G11
XG559 XI11_7/XI0/XI0_56/d_6_ XI11_7/XI0/XI0_56/d__6_ DECAP_INV_G11
XG560 XI11_7/XI0/XI0_56/d_5_ XI11_7/XI0/XI0_56/d__5_ DECAP_INV_G11
XG561 XI11_7/XI0/XI0_56/d_4_ XI11_7/XI0/XI0_56/d__4_ DECAP_INV_G11
XG562 XI11_7/XI0/XI0_56/d_3_ XI11_7/XI0/XI0_56/d__3_ DECAP_INV_G11
XG563 XI11_7/XI0/XI0_56/d_2_ XI11_7/XI0/XI0_56/d__2_ DECAP_INV_G11
XG564 XI11_7/XI0/XI0_56/d_1_ XI11_7/XI0/XI0_56/d__1_ DECAP_INV_G11
XG565 XI11_7/XI0/XI0_56/d_0_ XI11_7/XI0/XI0_56/d__0_ DECAP_INV_G11
XG566 XI11_7/XI0/XI0_55/d__15_ XI11_7/XI0/XI0_55/d_15_ DECAP_INV_G11
XG567 XI11_7/XI0/XI0_55/d__14_ XI11_7/XI0/XI0_55/d_14_ DECAP_INV_G11
XG568 XI11_7/XI0/XI0_55/d__13_ XI11_7/XI0/XI0_55/d_13_ DECAP_INV_G11
XG569 XI11_7/XI0/XI0_55/d__12_ XI11_7/XI0/XI0_55/d_12_ DECAP_INV_G11
XG570 XI11_7/XI0/XI0_55/d__11_ XI11_7/XI0/XI0_55/d_11_ DECAP_INV_G11
XG571 XI11_7/XI0/XI0_55/d__10_ XI11_7/XI0/XI0_55/d_10_ DECAP_INV_G11
XG572 XI11_7/XI0/XI0_55/d__9_ XI11_7/XI0/XI0_55/d_9_ DECAP_INV_G11
XG573 XI11_7/XI0/XI0_55/d__8_ XI11_7/XI0/XI0_55/d_8_ DECAP_INV_G11
XG574 XI11_7/XI0/XI0_55/d__7_ XI11_7/XI0/XI0_55/d_7_ DECAP_INV_G11
XG575 XI11_7/XI0/XI0_55/d__6_ XI11_7/XI0/XI0_55/d_6_ DECAP_INV_G11
XG576 XI11_7/XI0/XI0_55/d__5_ XI11_7/XI0/XI0_55/d_5_ DECAP_INV_G11
XG577 XI11_7/XI0/XI0_55/d__4_ XI11_7/XI0/XI0_55/d_4_ DECAP_INV_G11
XG578 XI11_7/XI0/XI0_55/d__3_ XI11_7/XI0/XI0_55/d_3_ DECAP_INV_G11
XG579 XI11_7/XI0/XI0_55/d__2_ XI11_7/XI0/XI0_55/d_2_ DECAP_INV_G11
XG580 XI11_7/XI0/XI0_55/d__1_ XI11_7/XI0/XI0_55/d_1_ DECAP_INV_G11
XG581 XI11_7/XI0/XI0_55/d__0_ XI11_7/XI0/XI0_55/d_0_ DECAP_INV_G11
XG582 XI11_7/XI0/XI0_55/d_15_ XI11_7/XI0/XI0_55/d__15_ DECAP_INV_G11
XG583 XI11_7/XI0/XI0_55/d_14_ XI11_7/XI0/XI0_55/d__14_ DECAP_INV_G11
XG584 XI11_7/XI0/XI0_55/d_13_ XI11_7/XI0/XI0_55/d__13_ DECAP_INV_G11
XG585 XI11_7/XI0/XI0_55/d_12_ XI11_7/XI0/XI0_55/d__12_ DECAP_INV_G11
XG586 XI11_7/XI0/XI0_55/d_11_ XI11_7/XI0/XI0_55/d__11_ DECAP_INV_G11
XG587 XI11_7/XI0/XI0_55/d_10_ XI11_7/XI0/XI0_55/d__10_ DECAP_INV_G11
XG588 XI11_7/XI0/XI0_55/d_9_ XI11_7/XI0/XI0_55/d__9_ DECAP_INV_G11
XG589 XI11_7/XI0/XI0_55/d_8_ XI11_7/XI0/XI0_55/d__8_ DECAP_INV_G11
XG590 XI11_7/XI0/XI0_55/d_7_ XI11_7/XI0/XI0_55/d__7_ DECAP_INV_G11
XG591 XI11_7/XI0/XI0_55/d_6_ XI11_7/XI0/XI0_55/d__6_ DECAP_INV_G11
XG592 XI11_7/XI0/XI0_55/d_5_ XI11_7/XI0/XI0_55/d__5_ DECAP_INV_G11
XG593 XI11_7/XI0/XI0_55/d_4_ XI11_7/XI0/XI0_55/d__4_ DECAP_INV_G11
XG594 XI11_7/XI0/XI0_55/d_3_ XI11_7/XI0/XI0_55/d__3_ DECAP_INV_G11
XG595 XI11_7/XI0/XI0_55/d_2_ XI11_7/XI0/XI0_55/d__2_ DECAP_INV_G11
XG596 XI11_7/XI0/XI0_55/d_1_ XI11_7/XI0/XI0_55/d__1_ DECAP_INV_G11
XG597 XI11_7/XI0/XI0_55/d_0_ XI11_7/XI0/XI0_55/d__0_ DECAP_INV_G11
XG598 XI11_7/XI0/XI0_54/d__15_ XI11_7/XI0/XI0_54/d_15_ DECAP_INV_G11
XG599 XI11_7/XI0/XI0_54/d__14_ XI11_7/XI0/XI0_54/d_14_ DECAP_INV_G11
XG600 XI11_7/XI0/XI0_54/d__13_ XI11_7/XI0/XI0_54/d_13_ DECAP_INV_G11
XG601 XI11_7/XI0/XI0_54/d__12_ XI11_7/XI0/XI0_54/d_12_ DECAP_INV_G11
XG602 XI11_7/XI0/XI0_54/d__11_ XI11_7/XI0/XI0_54/d_11_ DECAP_INV_G11
XG603 XI11_7/XI0/XI0_54/d__10_ XI11_7/XI0/XI0_54/d_10_ DECAP_INV_G11
XG604 XI11_7/XI0/XI0_54/d__9_ XI11_7/XI0/XI0_54/d_9_ DECAP_INV_G11
XG605 XI11_7/XI0/XI0_54/d__8_ XI11_7/XI0/XI0_54/d_8_ DECAP_INV_G11
XG606 XI11_7/XI0/XI0_54/d__7_ XI11_7/XI0/XI0_54/d_7_ DECAP_INV_G11
XG607 XI11_7/XI0/XI0_54/d__6_ XI11_7/XI0/XI0_54/d_6_ DECAP_INV_G11
XG608 XI11_7/XI0/XI0_54/d__5_ XI11_7/XI0/XI0_54/d_5_ DECAP_INV_G11
XG609 XI11_7/XI0/XI0_54/d__4_ XI11_7/XI0/XI0_54/d_4_ DECAP_INV_G11
XG610 XI11_7/XI0/XI0_54/d__3_ XI11_7/XI0/XI0_54/d_3_ DECAP_INV_G11
XG611 XI11_7/XI0/XI0_54/d__2_ XI11_7/XI0/XI0_54/d_2_ DECAP_INV_G11
XG612 XI11_7/XI0/XI0_54/d__1_ XI11_7/XI0/XI0_54/d_1_ DECAP_INV_G11
XG613 XI11_7/XI0/XI0_54/d__0_ XI11_7/XI0/XI0_54/d_0_ DECAP_INV_G11
XG614 XI11_7/XI0/XI0_54/d_15_ XI11_7/XI0/XI0_54/d__15_ DECAP_INV_G11
XG615 XI11_7/XI0/XI0_54/d_14_ XI11_7/XI0/XI0_54/d__14_ DECAP_INV_G11
XG616 XI11_7/XI0/XI0_54/d_13_ XI11_7/XI0/XI0_54/d__13_ DECAP_INV_G11
XG617 XI11_7/XI0/XI0_54/d_12_ XI11_7/XI0/XI0_54/d__12_ DECAP_INV_G11
XG618 XI11_7/XI0/XI0_54/d_11_ XI11_7/XI0/XI0_54/d__11_ DECAP_INV_G11
XG619 XI11_7/XI0/XI0_54/d_10_ XI11_7/XI0/XI0_54/d__10_ DECAP_INV_G11
XG620 XI11_7/XI0/XI0_54/d_9_ XI11_7/XI0/XI0_54/d__9_ DECAP_INV_G11
XG621 XI11_7/XI0/XI0_54/d_8_ XI11_7/XI0/XI0_54/d__8_ DECAP_INV_G11
XG622 XI11_7/XI0/XI0_54/d_7_ XI11_7/XI0/XI0_54/d__7_ DECAP_INV_G11
XG623 XI11_7/XI0/XI0_54/d_6_ XI11_7/XI0/XI0_54/d__6_ DECAP_INV_G11
XG624 XI11_7/XI0/XI0_54/d_5_ XI11_7/XI0/XI0_54/d__5_ DECAP_INV_G11
XG625 XI11_7/XI0/XI0_54/d_4_ XI11_7/XI0/XI0_54/d__4_ DECAP_INV_G11
XG626 XI11_7/XI0/XI0_54/d_3_ XI11_7/XI0/XI0_54/d__3_ DECAP_INV_G11
XG627 XI11_7/XI0/XI0_54/d_2_ XI11_7/XI0/XI0_54/d__2_ DECAP_INV_G11
XG628 XI11_7/XI0/XI0_54/d_1_ XI11_7/XI0/XI0_54/d__1_ DECAP_INV_G11
XG629 XI11_7/XI0/XI0_54/d_0_ XI11_7/XI0/XI0_54/d__0_ DECAP_INV_G11
XG630 XI11_7/XI0/XI0_53/d__15_ XI11_7/XI0/XI0_53/d_15_ DECAP_INV_G11
XG631 XI11_7/XI0/XI0_53/d__14_ XI11_7/XI0/XI0_53/d_14_ DECAP_INV_G11
XG632 XI11_7/XI0/XI0_53/d__13_ XI11_7/XI0/XI0_53/d_13_ DECAP_INV_G11
XG633 XI11_7/XI0/XI0_53/d__12_ XI11_7/XI0/XI0_53/d_12_ DECAP_INV_G11
XG634 XI11_7/XI0/XI0_53/d__11_ XI11_7/XI0/XI0_53/d_11_ DECAP_INV_G11
XG635 XI11_7/XI0/XI0_53/d__10_ XI11_7/XI0/XI0_53/d_10_ DECAP_INV_G11
XG636 XI11_7/XI0/XI0_53/d__9_ XI11_7/XI0/XI0_53/d_9_ DECAP_INV_G11
XG637 XI11_7/XI0/XI0_53/d__8_ XI11_7/XI0/XI0_53/d_8_ DECAP_INV_G11
XG638 XI11_7/XI0/XI0_53/d__7_ XI11_7/XI0/XI0_53/d_7_ DECAP_INV_G11
XG639 XI11_7/XI0/XI0_53/d__6_ XI11_7/XI0/XI0_53/d_6_ DECAP_INV_G11
XG640 XI11_7/XI0/XI0_53/d__5_ XI11_7/XI0/XI0_53/d_5_ DECAP_INV_G11
XG641 XI11_7/XI0/XI0_53/d__4_ XI11_7/XI0/XI0_53/d_4_ DECAP_INV_G11
XG642 XI11_7/XI0/XI0_53/d__3_ XI11_7/XI0/XI0_53/d_3_ DECAP_INV_G11
XG643 XI11_7/XI0/XI0_53/d__2_ XI11_7/XI0/XI0_53/d_2_ DECAP_INV_G11
XG644 XI11_7/XI0/XI0_53/d__1_ XI11_7/XI0/XI0_53/d_1_ DECAP_INV_G11
XG645 XI11_7/XI0/XI0_53/d__0_ XI11_7/XI0/XI0_53/d_0_ DECAP_INV_G11
XG646 XI11_7/XI0/XI0_53/d_15_ XI11_7/XI0/XI0_53/d__15_ DECAP_INV_G11
XG647 XI11_7/XI0/XI0_53/d_14_ XI11_7/XI0/XI0_53/d__14_ DECAP_INV_G11
XG648 XI11_7/XI0/XI0_53/d_13_ XI11_7/XI0/XI0_53/d__13_ DECAP_INV_G11
XG649 XI11_7/XI0/XI0_53/d_12_ XI11_7/XI0/XI0_53/d__12_ DECAP_INV_G11
XG650 XI11_7/XI0/XI0_53/d_11_ XI11_7/XI0/XI0_53/d__11_ DECAP_INV_G11
XG651 XI11_7/XI0/XI0_53/d_10_ XI11_7/XI0/XI0_53/d__10_ DECAP_INV_G11
XG652 XI11_7/XI0/XI0_53/d_9_ XI11_7/XI0/XI0_53/d__9_ DECAP_INV_G11
XG653 XI11_7/XI0/XI0_53/d_8_ XI11_7/XI0/XI0_53/d__8_ DECAP_INV_G11
XG654 XI11_7/XI0/XI0_53/d_7_ XI11_7/XI0/XI0_53/d__7_ DECAP_INV_G11
XG655 XI11_7/XI0/XI0_53/d_6_ XI11_7/XI0/XI0_53/d__6_ DECAP_INV_G11
XG656 XI11_7/XI0/XI0_53/d_5_ XI11_7/XI0/XI0_53/d__5_ DECAP_INV_G11
XG657 XI11_7/XI0/XI0_53/d_4_ XI11_7/XI0/XI0_53/d__4_ DECAP_INV_G11
XG658 XI11_7/XI0/XI0_53/d_3_ XI11_7/XI0/XI0_53/d__3_ DECAP_INV_G11
XG659 XI11_7/XI0/XI0_53/d_2_ XI11_7/XI0/XI0_53/d__2_ DECAP_INV_G11
XG660 XI11_7/XI0/XI0_53/d_1_ XI11_7/XI0/XI0_53/d__1_ DECAP_INV_G11
XG661 XI11_7/XI0/XI0_53/d_0_ XI11_7/XI0/XI0_53/d__0_ DECAP_INV_G11
XG662 XI11_7/XI0/XI0_52/d__15_ XI11_7/XI0/XI0_52/d_15_ DECAP_INV_G11
XG663 XI11_7/XI0/XI0_52/d__14_ XI11_7/XI0/XI0_52/d_14_ DECAP_INV_G11
XG664 XI11_7/XI0/XI0_52/d__13_ XI11_7/XI0/XI0_52/d_13_ DECAP_INV_G11
XG665 XI11_7/XI0/XI0_52/d__12_ XI11_7/XI0/XI0_52/d_12_ DECAP_INV_G11
XG666 XI11_7/XI0/XI0_52/d__11_ XI11_7/XI0/XI0_52/d_11_ DECAP_INV_G11
XG667 XI11_7/XI0/XI0_52/d__10_ XI11_7/XI0/XI0_52/d_10_ DECAP_INV_G11
XG668 XI11_7/XI0/XI0_52/d__9_ XI11_7/XI0/XI0_52/d_9_ DECAP_INV_G11
XG669 XI11_7/XI0/XI0_52/d__8_ XI11_7/XI0/XI0_52/d_8_ DECAP_INV_G11
XG670 XI11_7/XI0/XI0_52/d__7_ XI11_7/XI0/XI0_52/d_7_ DECAP_INV_G11
XG671 XI11_7/XI0/XI0_52/d__6_ XI11_7/XI0/XI0_52/d_6_ DECAP_INV_G11
XG672 XI11_7/XI0/XI0_52/d__5_ XI11_7/XI0/XI0_52/d_5_ DECAP_INV_G11
XG673 XI11_7/XI0/XI0_52/d__4_ XI11_7/XI0/XI0_52/d_4_ DECAP_INV_G11
XG674 XI11_7/XI0/XI0_52/d__3_ XI11_7/XI0/XI0_52/d_3_ DECAP_INV_G11
XG675 XI11_7/XI0/XI0_52/d__2_ XI11_7/XI0/XI0_52/d_2_ DECAP_INV_G11
XG676 XI11_7/XI0/XI0_52/d__1_ XI11_7/XI0/XI0_52/d_1_ DECAP_INV_G11
XG677 XI11_7/XI0/XI0_52/d__0_ XI11_7/XI0/XI0_52/d_0_ DECAP_INV_G11
XG678 XI11_7/XI0/XI0_52/d_15_ XI11_7/XI0/XI0_52/d__15_ DECAP_INV_G11
XG679 XI11_7/XI0/XI0_52/d_14_ XI11_7/XI0/XI0_52/d__14_ DECAP_INV_G11
XG680 XI11_7/XI0/XI0_52/d_13_ XI11_7/XI0/XI0_52/d__13_ DECAP_INV_G11
XG681 XI11_7/XI0/XI0_52/d_12_ XI11_7/XI0/XI0_52/d__12_ DECAP_INV_G11
XG682 XI11_7/XI0/XI0_52/d_11_ XI11_7/XI0/XI0_52/d__11_ DECAP_INV_G11
XG683 XI11_7/XI0/XI0_52/d_10_ XI11_7/XI0/XI0_52/d__10_ DECAP_INV_G11
XG684 XI11_7/XI0/XI0_52/d_9_ XI11_7/XI0/XI0_52/d__9_ DECAP_INV_G11
XG685 XI11_7/XI0/XI0_52/d_8_ XI11_7/XI0/XI0_52/d__8_ DECAP_INV_G11
XG686 XI11_7/XI0/XI0_52/d_7_ XI11_7/XI0/XI0_52/d__7_ DECAP_INV_G11
XG687 XI11_7/XI0/XI0_52/d_6_ XI11_7/XI0/XI0_52/d__6_ DECAP_INV_G11
XG688 XI11_7/XI0/XI0_52/d_5_ XI11_7/XI0/XI0_52/d__5_ DECAP_INV_G11
XG689 XI11_7/XI0/XI0_52/d_4_ XI11_7/XI0/XI0_52/d__4_ DECAP_INV_G11
XG690 XI11_7/XI0/XI0_52/d_3_ XI11_7/XI0/XI0_52/d__3_ DECAP_INV_G11
XG691 XI11_7/XI0/XI0_52/d_2_ XI11_7/XI0/XI0_52/d__2_ DECAP_INV_G11
XG692 XI11_7/XI0/XI0_52/d_1_ XI11_7/XI0/XI0_52/d__1_ DECAP_INV_G11
XG693 XI11_7/XI0/XI0_52/d_0_ XI11_7/XI0/XI0_52/d__0_ DECAP_INV_G11
XG694 XI11_7/XI0/XI0_51/d__15_ XI11_7/XI0/XI0_51/d_15_ DECAP_INV_G11
XG695 XI11_7/XI0/XI0_51/d__14_ XI11_7/XI0/XI0_51/d_14_ DECAP_INV_G11
XG696 XI11_7/XI0/XI0_51/d__13_ XI11_7/XI0/XI0_51/d_13_ DECAP_INV_G11
XG697 XI11_7/XI0/XI0_51/d__12_ XI11_7/XI0/XI0_51/d_12_ DECAP_INV_G11
XG698 XI11_7/XI0/XI0_51/d__11_ XI11_7/XI0/XI0_51/d_11_ DECAP_INV_G11
XG699 XI11_7/XI0/XI0_51/d__10_ XI11_7/XI0/XI0_51/d_10_ DECAP_INV_G11
XG700 XI11_7/XI0/XI0_51/d__9_ XI11_7/XI0/XI0_51/d_9_ DECAP_INV_G11
XG701 XI11_7/XI0/XI0_51/d__8_ XI11_7/XI0/XI0_51/d_8_ DECAP_INV_G11
XG702 XI11_7/XI0/XI0_51/d__7_ XI11_7/XI0/XI0_51/d_7_ DECAP_INV_G11
XG703 XI11_7/XI0/XI0_51/d__6_ XI11_7/XI0/XI0_51/d_6_ DECAP_INV_G11
XG704 XI11_7/XI0/XI0_51/d__5_ XI11_7/XI0/XI0_51/d_5_ DECAP_INV_G11
XG705 XI11_7/XI0/XI0_51/d__4_ XI11_7/XI0/XI0_51/d_4_ DECAP_INV_G11
XG706 XI11_7/XI0/XI0_51/d__3_ XI11_7/XI0/XI0_51/d_3_ DECAP_INV_G11
XG707 XI11_7/XI0/XI0_51/d__2_ XI11_7/XI0/XI0_51/d_2_ DECAP_INV_G11
XG708 XI11_7/XI0/XI0_51/d__1_ XI11_7/XI0/XI0_51/d_1_ DECAP_INV_G11
XG709 XI11_7/XI0/XI0_51/d__0_ XI11_7/XI0/XI0_51/d_0_ DECAP_INV_G11
XG710 XI11_7/XI0/XI0_51/d_15_ XI11_7/XI0/XI0_51/d__15_ DECAP_INV_G11
XG711 XI11_7/XI0/XI0_51/d_14_ XI11_7/XI0/XI0_51/d__14_ DECAP_INV_G11
XG712 XI11_7/XI0/XI0_51/d_13_ XI11_7/XI0/XI0_51/d__13_ DECAP_INV_G11
XG713 XI11_7/XI0/XI0_51/d_12_ XI11_7/XI0/XI0_51/d__12_ DECAP_INV_G11
XG714 XI11_7/XI0/XI0_51/d_11_ XI11_7/XI0/XI0_51/d__11_ DECAP_INV_G11
XG715 XI11_7/XI0/XI0_51/d_10_ XI11_7/XI0/XI0_51/d__10_ DECAP_INV_G11
XG716 XI11_7/XI0/XI0_51/d_9_ XI11_7/XI0/XI0_51/d__9_ DECAP_INV_G11
XG717 XI11_7/XI0/XI0_51/d_8_ XI11_7/XI0/XI0_51/d__8_ DECAP_INV_G11
XG718 XI11_7/XI0/XI0_51/d_7_ XI11_7/XI0/XI0_51/d__7_ DECAP_INV_G11
XG719 XI11_7/XI0/XI0_51/d_6_ XI11_7/XI0/XI0_51/d__6_ DECAP_INV_G11
XG720 XI11_7/XI0/XI0_51/d_5_ XI11_7/XI0/XI0_51/d__5_ DECAP_INV_G11
XG721 XI11_7/XI0/XI0_51/d_4_ XI11_7/XI0/XI0_51/d__4_ DECAP_INV_G11
XG722 XI11_7/XI0/XI0_51/d_3_ XI11_7/XI0/XI0_51/d__3_ DECAP_INV_G11
XG723 XI11_7/XI0/XI0_51/d_2_ XI11_7/XI0/XI0_51/d__2_ DECAP_INV_G11
XG724 XI11_7/XI0/XI0_51/d_1_ XI11_7/XI0/XI0_51/d__1_ DECAP_INV_G11
XG725 XI11_7/XI0/XI0_51/d_0_ XI11_7/XI0/XI0_51/d__0_ DECAP_INV_G11
XG726 XI11_7/XI0/XI0_50/d__15_ XI11_7/XI0/XI0_50/d_15_ DECAP_INV_G11
XG727 XI11_7/XI0/XI0_50/d__14_ XI11_7/XI0/XI0_50/d_14_ DECAP_INV_G11
XG728 XI11_7/XI0/XI0_50/d__13_ XI11_7/XI0/XI0_50/d_13_ DECAP_INV_G11
XG729 XI11_7/XI0/XI0_50/d__12_ XI11_7/XI0/XI0_50/d_12_ DECAP_INV_G11
XG730 XI11_7/XI0/XI0_50/d__11_ XI11_7/XI0/XI0_50/d_11_ DECAP_INV_G11
XG731 XI11_7/XI0/XI0_50/d__10_ XI11_7/XI0/XI0_50/d_10_ DECAP_INV_G11
XG732 XI11_7/XI0/XI0_50/d__9_ XI11_7/XI0/XI0_50/d_9_ DECAP_INV_G11
XG733 XI11_7/XI0/XI0_50/d__8_ XI11_7/XI0/XI0_50/d_8_ DECAP_INV_G11
XG734 XI11_7/XI0/XI0_50/d__7_ XI11_7/XI0/XI0_50/d_7_ DECAP_INV_G11
XG735 XI11_7/XI0/XI0_50/d__6_ XI11_7/XI0/XI0_50/d_6_ DECAP_INV_G11
XG736 XI11_7/XI0/XI0_50/d__5_ XI11_7/XI0/XI0_50/d_5_ DECAP_INV_G11
XG737 XI11_7/XI0/XI0_50/d__4_ XI11_7/XI0/XI0_50/d_4_ DECAP_INV_G11
XG738 XI11_7/XI0/XI0_50/d__3_ XI11_7/XI0/XI0_50/d_3_ DECAP_INV_G11
XG739 XI11_7/XI0/XI0_50/d__2_ XI11_7/XI0/XI0_50/d_2_ DECAP_INV_G11
XG740 XI11_7/XI0/XI0_50/d__1_ XI11_7/XI0/XI0_50/d_1_ DECAP_INV_G11
XG741 XI11_7/XI0/XI0_50/d__0_ XI11_7/XI0/XI0_50/d_0_ DECAP_INV_G11
XG742 XI11_7/XI0/XI0_50/d_15_ XI11_7/XI0/XI0_50/d__15_ DECAP_INV_G11
XG743 XI11_7/XI0/XI0_50/d_14_ XI11_7/XI0/XI0_50/d__14_ DECAP_INV_G11
XG744 XI11_7/XI0/XI0_50/d_13_ XI11_7/XI0/XI0_50/d__13_ DECAP_INV_G11
XG745 XI11_7/XI0/XI0_50/d_12_ XI11_7/XI0/XI0_50/d__12_ DECAP_INV_G11
XG746 XI11_7/XI0/XI0_50/d_11_ XI11_7/XI0/XI0_50/d__11_ DECAP_INV_G11
XG747 XI11_7/XI0/XI0_50/d_10_ XI11_7/XI0/XI0_50/d__10_ DECAP_INV_G11
XG748 XI11_7/XI0/XI0_50/d_9_ XI11_7/XI0/XI0_50/d__9_ DECAP_INV_G11
XG749 XI11_7/XI0/XI0_50/d_8_ XI11_7/XI0/XI0_50/d__8_ DECAP_INV_G11
XG750 XI11_7/XI0/XI0_50/d_7_ XI11_7/XI0/XI0_50/d__7_ DECAP_INV_G11
XG751 XI11_7/XI0/XI0_50/d_6_ XI11_7/XI0/XI0_50/d__6_ DECAP_INV_G11
XG752 XI11_7/XI0/XI0_50/d_5_ XI11_7/XI0/XI0_50/d__5_ DECAP_INV_G11
XG753 XI11_7/XI0/XI0_50/d_4_ XI11_7/XI0/XI0_50/d__4_ DECAP_INV_G11
XG754 XI11_7/XI0/XI0_50/d_3_ XI11_7/XI0/XI0_50/d__3_ DECAP_INV_G11
XG755 XI11_7/XI0/XI0_50/d_2_ XI11_7/XI0/XI0_50/d__2_ DECAP_INV_G11
XG756 XI11_7/XI0/XI0_50/d_1_ XI11_7/XI0/XI0_50/d__1_ DECAP_INV_G11
XG757 XI11_7/XI0/XI0_50/d_0_ XI11_7/XI0/XI0_50/d__0_ DECAP_INV_G11
XG758 XI11_7/XI0/XI0_49/d__15_ XI11_7/XI0/XI0_49/d_15_ DECAP_INV_G11
XG759 XI11_7/XI0/XI0_49/d__14_ XI11_7/XI0/XI0_49/d_14_ DECAP_INV_G11
XG760 XI11_7/XI0/XI0_49/d__13_ XI11_7/XI0/XI0_49/d_13_ DECAP_INV_G11
XG761 XI11_7/XI0/XI0_49/d__12_ XI11_7/XI0/XI0_49/d_12_ DECAP_INV_G11
XG762 XI11_7/XI0/XI0_49/d__11_ XI11_7/XI0/XI0_49/d_11_ DECAP_INV_G11
XG763 XI11_7/XI0/XI0_49/d__10_ XI11_7/XI0/XI0_49/d_10_ DECAP_INV_G11
XG764 XI11_7/XI0/XI0_49/d__9_ XI11_7/XI0/XI0_49/d_9_ DECAP_INV_G11
XG765 XI11_7/XI0/XI0_49/d__8_ XI11_7/XI0/XI0_49/d_8_ DECAP_INV_G11
XG766 XI11_7/XI0/XI0_49/d__7_ XI11_7/XI0/XI0_49/d_7_ DECAP_INV_G11
XG767 XI11_7/XI0/XI0_49/d__6_ XI11_7/XI0/XI0_49/d_6_ DECAP_INV_G11
XG768 XI11_7/XI0/XI0_49/d__5_ XI11_7/XI0/XI0_49/d_5_ DECAP_INV_G11
XG769 XI11_7/XI0/XI0_49/d__4_ XI11_7/XI0/XI0_49/d_4_ DECAP_INV_G11
XG770 XI11_7/XI0/XI0_49/d__3_ XI11_7/XI0/XI0_49/d_3_ DECAP_INV_G11
XG771 XI11_7/XI0/XI0_49/d__2_ XI11_7/XI0/XI0_49/d_2_ DECAP_INV_G11
XG772 XI11_7/XI0/XI0_49/d__1_ XI11_7/XI0/XI0_49/d_1_ DECAP_INV_G11
XG773 XI11_7/XI0/XI0_49/d__0_ XI11_7/XI0/XI0_49/d_0_ DECAP_INV_G11
XG774 XI11_7/XI0/XI0_49/d_15_ XI11_7/XI0/XI0_49/d__15_ DECAP_INV_G11
XG775 XI11_7/XI0/XI0_49/d_14_ XI11_7/XI0/XI0_49/d__14_ DECAP_INV_G11
XG776 XI11_7/XI0/XI0_49/d_13_ XI11_7/XI0/XI0_49/d__13_ DECAP_INV_G11
XG777 XI11_7/XI0/XI0_49/d_12_ XI11_7/XI0/XI0_49/d__12_ DECAP_INV_G11
XG778 XI11_7/XI0/XI0_49/d_11_ XI11_7/XI0/XI0_49/d__11_ DECAP_INV_G11
XG779 XI11_7/XI0/XI0_49/d_10_ XI11_7/XI0/XI0_49/d__10_ DECAP_INV_G11
XG780 XI11_7/XI0/XI0_49/d_9_ XI11_7/XI0/XI0_49/d__9_ DECAP_INV_G11
XG781 XI11_7/XI0/XI0_49/d_8_ XI11_7/XI0/XI0_49/d__8_ DECAP_INV_G11
XG782 XI11_7/XI0/XI0_49/d_7_ XI11_7/XI0/XI0_49/d__7_ DECAP_INV_G11
XG783 XI11_7/XI0/XI0_49/d_6_ XI11_7/XI0/XI0_49/d__6_ DECAP_INV_G11
XG784 XI11_7/XI0/XI0_49/d_5_ XI11_7/XI0/XI0_49/d__5_ DECAP_INV_G11
XG785 XI11_7/XI0/XI0_49/d_4_ XI11_7/XI0/XI0_49/d__4_ DECAP_INV_G11
XG786 XI11_7/XI0/XI0_49/d_3_ XI11_7/XI0/XI0_49/d__3_ DECAP_INV_G11
XG787 XI11_7/XI0/XI0_49/d_2_ XI11_7/XI0/XI0_49/d__2_ DECAP_INV_G11
XG788 XI11_7/XI0/XI0_49/d_1_ XI11_7/XI0/XI0_49/d__1_ DECAP_INV_G11
XG789 XI11_7/XI0/XI0_49/d_0_ XI11_7/XI0/XI0_49/d__0_ DECAP_INV_G11
XG790 XI11_7/XI0/XI0_48/d__15_ XI11_7/XI0/XI0_48/d_15_ DECAP_INV_G11
XG791 XI11_7/XI0/XI0_48/d__14_ XI11_7/XI0/XI0_48/d_14_ DECAP_INV_G11
XG792 XI11_7/XI0/XI0_48/d__13_ XI11_7/XI0/XI0_48/d_13_ DECAP_INV_G11
XG793 XI11_7/XI0/XI0_48/d__12_ XI11_7/XI0/XI0_48/d_12_ DECAP_INV_G11
XG794 XI11_7/XI0/XI0_48/d__11_ XI11_7/XI0/XI0_48/d_11_ DECAP_INV_G11
XG795 XI11_7/XI0/XI0_48/d__10_ XI11_7/XI0/XI0_48/d_10_ DECAP_INV_G11
XG796 XI11_7/XI0/XI0_48/d__9_ XI11_7/XI0/XI0_48/d_9_ DECAP_INV_G11
XG797 XI11_7/XI0/XI0_48/d__8_ XI11_7/XI0/XI0_48/d_8_ DECAP_INV_G11
XG798 XI11_7/XI0/XI0_48/d__7_ XI11_7/XI0/XI0_48/d_7_ DECAP_INV_G11
XG799 XI11_7/XI0/XI0_48/d__6_ XI11_7/XI0/XI0_48/d_6_ DECAP_INV_G11
XG800 XI11_7/XI0/XI0_48/d__5_ XI11_7/XI0/XI0_48/d_5_ DECAP_INV_G11
XG801 XI11_7/XI0/XI0_48/d__4_ XI11_7/XI0/XI0_48/d_4_ DECAP_INV_G11
XG802 XI11_7/XI0/XI0_48/d__3_ XI11_7/XI0/XI0_48/d_3_ DECAP_INV_G11
XG803 XI11_7/XI0/XI0_48/d__2_ XI11_7/XI0/XI0_48/d_2_ DECAP_INV_G11
XG804 XI11_7/XI0/XI0_48/d__1_ XI11_7/XI0/XI0_48/d_1_ DECAP_INV_G11
XG805 XI11_7/XI0/XI0_48/d__0_ XI11_7/XI0/XI0_48/d_0_ DECAP_INV_G11
XG806 XI11_7/XI0/XI0_48/d_15_ XI11_7/XI0/XI0_48/d__15_ DECAP_INV_G11
XG807 XI11_7/XI0/XI0_48/d_14_ XI11_7/XI0/XI0_48/d__14_ DECAP_INV_G11
XG808 XI11_7/XI0/XI0_48/d_13_ XI11_7/XI0/XI0_48/d__13_ DECAP_INV_G11
XG809 XI11_7/XI0/XI0_48/d_12_ XI11_7/XI0/XI0_48/d__12_ DECAP_INV_G11
XG810 XI11_7/XI0/XI0_48/d_11_ XI11_7/XI0/XI0_48/d__11_ DECAP_INV_G11
XG811 XI11_7/XI0/XI0_48/d_10_ XI11_7/XI0/XI0_48/d__10_ DECAP_INV_G11
XG812 XI11_7/XI0/XI0_48/d_9_ XI11_7/XI0/XI0_48/d__9_ DECAP_INV_G11
XG813 XI11_7/XI0/XI0_48/d_8_ XI11_7/XI0/XI0_48/d__8_ DECAP_INV_G11
XG814 XI11_7/XI0/XI0_48/d_7_ XI11_7/XI0/XI0_48/d__7_ DECAP_INV_G11
XG815 XI11_7/XI0/XI0_48/d_6_ XI11_7/XI0/XI0_48/d__6_ DECAP_INV_G11
XG816 XI11_7/XI0/XI0_48/d_5_ XI11_7/XI0/XI0_48/d__5_ DECAP_INV_G11
XG817 XI11_7/XI0/XI0_48/d_4_ XI11_7/XI0/XI0_48/d__4_ DECAP_INV_G11
XG818 XI11_7/XI0/XI0_48/d_3_ XI11_7/XI0/XI0_48/d__3_ DECAP_INV_G11
XG819 XI11_7/XI0/XI0_48/d_2_ XI11_7/XI0/XI0_48/d__2_ DECAP_INV_G11
XG820 XI11_7/XI0/XI0_48/d_1_ XI11_7/XI0/XI0_48/d__1_ DECAP_INV_G11
XG821 XI11_7/XI0/XI0_48/d_0_ XI11_7/XI0/XI0_48/d__0_ DECAP_INV_G11
XG822 XI11_7/XI0/XI0_47/d__15_ XI11_7/XI0/XI0_47/d_15_ DECAP_INV_G11
XG823 XI11_7/XI0/XI0_47/d__14_ XI11_7/XI0/XI0_47/d_14_ DECAP_INV_G11
XG824 XI11_7/XI0/XI0_47/d__13_ XI11_7/XI0/XI0_47/d_13_ DECAP_INV_G11
XG825 XI11_7/XI0/XI0_47/d__12_ XI11_7/XI0/XI0_47/d_12_ DECAP_INV_G11
XG826 XI11_7/XI0/XI0_47/d__11_ XI11_7/XI0/XI0_47/d_11_ DECAP_INV_G11
XG827 XI11_7/XI0/XI0_47/d__10_ XI11_7/XI0/XI0_47/d_10_ DECAP_INV_G11
XG828 XI11_7/XI0/XI0_47/d__9_ XI11_7/XI0/XI0_47/d_9_ DECAP_INV_G11
XG829 XI11_7/XI0/XI0_47/d__8_ XI11_7/XI0/XI0_47/d_8_ DECAP_INV_G11
XG830 XI11_7/XI0/XI0_47/d__7_ XI11_7/XI0/XI0_47/d_7_ DECAP_INV_G11
XG831 XI11_7/XI0/XI0_47/d__6_ XI11_7/XI0/XI0_47/d_6_ DECAP_INV_G11
XG832 XI11_7/XI0/XI0_47/d__5_ XI11_7/XI0/XI0_47/d_5_ DECAP_INV_G11
XG833 XI11_7/XI0/XI0_47/d__4_ XI11_7/XI0/XI0_47/d_4_ DECAP_INV_G11
XG834 XI11_7/XI0/XI0_47/d__3_ XI11_7/XI0/XI0_47/d_3_ DECAP_INV_G11
XG835 XI11_7/XI0/XI0_47/d__2_ XI11_7/XI0/XI0_47/d_2_ DECAP_INV_G11
XG836 XI11_7/XI0/XI0_47/d__1_ XI11_7/XI0/XI0_47/d_1_ DECAP_INV_G11
XG837 XI11_7/XI0/XI0_47/d__0_ XI11_7/XI0/XI0_47/d_0_ DECAP_INV_G11
XG838 XI11_7/XI0/XI0_47/d_15_ XI11_7/XI0/XI0_47/d__15_ DECAP_INV_G11
XG839 XI11_7/XI0/XI0_47/d_14_ XI11_7/XI0/XI0_47/d__14_ DECAP_INV_G11
XG840 XI11_7/XI0/XI0_47/d_13_ XI11_7/XI0/XI0_47/d__13_ DECAP_INV_G11
XG841 XI11_7/XI0/XI0_47/d_12_ XI11_7/XI0/XI0_47/d__12_ DECAP_INV_G11
XG842 XI11_7/XI0/XI0_47/d_11_ XI11_7/XI0/XI0_47/d__11_ DECAP_INV_G11
XG843 XI11_7/XI0/XI0_47/d_10_ XI11_7/XI0/XI0_47/d__10_ DECAP_INV_G11
XG844 XI11_7/XI0/XI0_47/d_9_ XI11_7/XI0/XI0_47/d__9_ DECAP_INV_G11
XG845 XI11_7/XI0/XI0_47/d_8_ XI11_7/XI0/XI0_47/d__8_ DECAP_INV_G11
XG846 XI11_7/XI0/XI0_47/d_7_ XI11_7/XI0/XI0_47/d__7_ DECAP_INV_G11
XG847 XI11_7/XI0/XI0_47/d_6_ XI11_7/XI0/XI0_47/d__6_ DECAP_INV_G11
XG848 XI11_7/XI0/XI0_47/d_5_ XI11_7/XI0/XI0_47/d__5_ DECAP_INV_G11
XG849 XI11_7/XI0/XI0_47/d_4_ XI11_7/XI0/XI0_47/d__4_ DECAP_INV_G11
XG850 XI11_7/XI0/XI0_47/d_3_ XI11_7/XI0/XI0_47/d__3_ DECAP_INV_G11
XG851 XI11_7/XI0/XI0_47/d_2_ XI11_7/XI0/XI0_47/d__2_ DECAP_INV_G11
XG852 XI11_7/XI0/XI0_47/d_1_ XI11_7/XI0/XI0_47/d__1_ DECAP_INV_G11
XG853 XI11_7/XI0/XI0_47/d_0_ XI11_7/XI0/XI0_47/d__0_ DECAP_INV_G11
XG854 XI11_7/XI0/XI0_46/d__15_ XI11_7/XI0/XI0_46/d_15_ DECAP_INV_G11
XG855 XI11_7/XI0/XI0_46/d__14_ XI11_7/XI0/XI0_46/d_14_ DECAP_INV_G11
XG856 XI11_7/XI0/XI0_46/d__13_ XI11_7/XI0/XI0_46/d_13_ DECAP_INV_G11
XG857 XI11_7/XI0/XI0_46/d__12_ XI11_7/XI0/XI0_46/d_12_ DECAP_INV_G11
XG858 XI11_7/XI0/XI0_46/d__11_ XI11_7/XI0/XI0_46/d_11_ DECAP_INV_G11
XG859 XI11_7/XI0/XI0_46/d__10_ XI11_7/XI0/XI0_46/d_10_ DECAP_INV_G11
XG860 XI11_7/XI0/XI0_46/d__9_ XI11_7/XI0/XI0_46/d_9_ DECAP_INV_G11
XG861 XI11_7/XI0/XI0_46/d__8_ XI11_7/XI0/XI0_46/d_8_ DECAP_INV_G11
XG862 XI11_7/XI0/XI0_46/d__7_ XI11_7/XI0/XI0_46/d_7_ DECAP_INV_G11
XG863 XI11_7/XI0/XI0_46/d__6_ XI11_7/XI0/XI0_46/d_6_ DECAP_INV_G11
XG864 XI11_7/XI0/XI0_46/d__5_ XI11_7/XI0/XI0_46/d_5_ DECAP_INV_G11
XG865 XI11_7/XI0/XI0_46/d__4_ XI11_7/XI0/XI0_46/d_4_ DECAP_INV_G11
XG866 XI11_7/XI0/XI0_46/d__3_ XI11_7/XI0/XI0_46/d_3_ DECAP_INV_G11
XG867 XI11_7/XI0/XI0_46/d__2_ XI11_7/XI0/XI0_46/d_2_ DECAP_INV_G11
XG868 XI11_7/XI0/XI0_46/d__1_ XI11_7/XI0/XI0_46/d_1_ DECAP_INV_G11
XG869 XI11_7/XI0/XI0_46/d__0_ XI11_7/XI0/XI0_46/d_0_ DECAP_INV_G11
XG870 XI11_7/XI0/XI0_46/d_15_ XI11_7/XI0/XI0_46/d__15_ DECAP_INV_G11
XG871 XI11_7/XI0/XI0_46/d_14_ XI11_7/XI0/XI0_46/d__14_ DECAP_INV_G11
XG872 XI11_7/XI0/XI0_46/d_13_ XI11_7/XI0/XI0_46/d__13_ DECAP_INV_G11
XG873 XI11_7/XI0/XI0_46/d_12_ XI11_7/XI0/XI0_46/d__12_ DECAP_INV_G11
XG874 XI11_7/XI0/XI0_46/d_11_ XI11_7/XI0/XI0_46/d__11_ DECAP_INV_G11
XG875 XI11_7/XI0/XI0_46/d_10_ XI11_7/XI0/XI0_46/d__10_ DECAP_INV_G11
XG876 XI11_7/XI0/XI0_46/d_9_ XI11_7/XI0/XI0_46/d__9_ DECAP_INV_G11
XG877 XI11_7/XI0/XI0_46/d_8_ XI11_7/XI0/XI0_46/d__8_ DECAP_INV_G11
XG878 XI11_7/XI0/XI0_46/d_7_ XI11_7/XI0/XI0_46/d__7_ DECAP_INV_G11
XG879 XI11_7/XI0/XI0_46/d_6_ XI11_7/XI0/XI0_46/d__6_ DECAP_INV_G11
XG880 XI11_7/XI0/XI0_46/d_5_ XI11_7/XI0/XI0_46/d__5_ DECAP_INV_G11
XG881 XI11_7/XI0/XI0_46/d_4_ XI11_7/XI0/XI0_46/d__4_ DECAP_INV_G11
XG882 XI11_7/XI0/XI0_46/d_3_ XI11_7/XI0/XI0_46/d__3_ DECAP_INV_G11
XG883 XI11_7/XI0/XI0_46/d_2_ XI11_7/XI0/XI0_46/d__2_ DECAP_INV_G11
XG884 XI11_7/XI0/XI0_46/d_1_ XI11_7/XI0/XI0_46/d__1_ DECAP_INV_G11
XG885 XI11_7/XI0/XI0_46/d_0_ XI11_7/XI0/XI0_46/d__0_ DECAP_INV_G11
XG886 XI11_7/XI0/XI0_45/d__15_ XI11_7/XI0/XI0_45/d_15_ DECAP_INV_G11
XG887 XI11_7/XI0/XI0_45/d__14_ XI11_7/XI0/XI0_45/d_14_ DECAP_INV_G11
XG888 XI11_7/XI0/XI0_45/d__13_ XI11_7/XI0/XI0_45/d_13_ DECAP_INV_G11
XG889 XI11_7/XI0/XI0_45/d__12_ XI11_7/XI0/XI0_45/d_12_ DECAP_INV_G11
XG890 XI11_7/XI0/XI0_45/d__11_ XI11_7/XI0/XI0_45/d_11_ DECAP_INV_G11
XG891 XI11_7/XI0/XI0_45/d__10_ XI11_7/XI0/XI0_45/d_10_ DECAP_INV_G11
XG892 XI11_7/XI0/XI0_45/d__9_ XI11_7/XI0/XI0_45/d_9_ DECAP_INV_G11
XG893 XI11_7/XI0/XI0_45/d__8_ XI11_7/XI0/XI0_45/d_8_ DECAP_INV_G11
XG894 XI11_7/XI0/XI0_45/d__7_ XI11_7/XI0/XI0_45/d_7_ DECAP_INV_G11
XG895 XI11_7/XI0/XI0_45/d__6_ XI11_7/XI0/XI0_45/d_6_ DECAP_INV_G11
XG896 XI11_7/XI0/XI0_45/d__5_ XI11_7/XI0/XI0_45/d_5_ DECAP_INV_G11
XG897 XI11_7/XI0/XI0_45/d__4_ XI11_7/XI0/XI0_45/d_4_ DECAP_INV_G11
XG898 XI11_7/XI0/XI0_45/d__3_ XI11_7/XI0/XI0_45/d_3_ DECAP_INV_G11
XG899 XI11_7/XI0/XI0_45/d__2_ XI11_7/XI0/XI0_45/d_2_ DECAP_INV_G11
XG900 XI11_7/XI0/XI0_45/d__1_ XI11_7/XI0/XI0_45/d_1_ DECAP_INV_G11
XG901 XI11_7/XI0/XI0_45/d__0_ XI11_7/XI0/XI0_45/d_0_ DECAP_INV_G11
XG902 XI11_7/XI0/XI0_45/d_15_ XI11_7/XI0/XI0_45/d__15_ DECAP_INV_G11
XG903 XI11_7/XI0/XI0_45/d_14_ XI11_7/XI0/XI0_45/d__14_ DECAP_INV_G11
XG904 XI11_7/XI0/XI0_45/d_13_ XI11_7/XI0/XI0_45/d__13_ DECAP_INV_G11
XG905 XI11_7/XI0/XI0_45/d_12_ XI11_7/XI0/XI0_45/d__12_ DECAP_INV_G11
XG906 XI11_7/XI0/XI0_45/d_11_ XI11_7/XI0/XI0_45/d__11_ DECAP_INV_G11
XG907 XI11_7/XI0/XI0_45/d_10_ XI11_7/XI0/XI0_45/d__10_ DECAP_INV_G11
XG908 XI11_7/XI0/XI0_45/d_9_ XI11_7/XI0/XI0_45/d__9_ DECAP_INV_G11
XG909 XI11_7/XI0/XI0_45/d_8_ XI11_7/XI0/XI0_45/d__8_ DECAP_INV_G11
XG910 XI11_7/XI0/XI0_45/d_7_ XI11_7/XI0/XI0_45/d__7_ DECAP_INV_G11
XG911 XI11_7/XI0/XI0_45/d_6_ XI11_7/XI0/XI0_45/d__6_ DECAP_INV_G11
XG912 XI11_7/XI0/XI0_45/d_5_ XI11_7/XI0/XI0_45/d__5_ DECAP_INV_G11
XG913 XI11_7/XI0/XI0_45/d_4_ XI11_7/XI0/XI0_45/d__4_ DECAP_INV_G11
XG914 XI11_7/XI0/XI0_45/d_3_ XI11_7/XI0/XI0_45/d__3_ DECAP_INV_G11
XG915 XI11_7/XI0/XI0_45/d_2_ XI11_7/XI0/XI0_45/d__2_ DECAP_INV_G11
XG916 XI11_7/XI0/XI0_45/d_1_ XI11_7/XI0/XI0_45/d__1_ DECAP_INV_G11
XG917 XI11_7/XI0/XI0_45/d_0_ XI11_7/XI0/XI0_45/d__0_ DECAP_INV_G11
XG918 XI11_7/XI0/XI0_44/d__15_ XI11_7/XI0/XI0_44/d_15_ DECAP_INV_G11
XG919 XI11_7/XI0/XI0_44/d__14_ XI11_7/XI0/XI0_44/d_14_ DECAP_INV_G11
XG920 XI11_7/XI0/XI0_44/d__13_ XI11_7/XI0/XI0_44/d_13_ DECAP_INV_G11
XG921 XI11_7/XI0/XI0_44/d__12_ XI11_7/XI0/XI0_44/d_12_ DECAP_INV_G11
XG922 XI11_7/XI0/XI0_44/d__11_ XI11_7/XI0/XI0_44/d_11_ DECAP_INV_G11
XG923 XI11_7/XI0/XI0_44/d__10_ XI11_7/XI0/XI0_44/d_10_ DECAP_INV_G11
XG924 XI11_7/XI0/XI0_44/d__9_ XI11_7/XI0/XI0_44/d_9_ DECAP_INV_G11
XG925 XI11_7/XI0/XI0_44/d__8_ XI11_7/XI0/XI0_44/d_8_ DECAP_INV_G11
XG926 XI11_7/XI0/XI0_44/d__7_ XI11_7/XI0/XI0_44/d_7_ DECAP_INV_G11
XG927 XI11_7/XI0/XI0_44/d__6_ XI11_7/XI0/XI0_44/d_6_ DECAP_INV_G11
XG928 XI11_7/XI0/XI0_44/d__5_ XI11_7/XI0/XI0_44/d_5_ DECAP_INV_G11
XG929 XI11_7/XI0/XI0_44/d__4_ XI11_7/XI0/XI0_44/d_4_ DECAP_INV_G11
XG930 XI11_7/XI0/XI0_44/d__3_ XI11_7/XI0/XI0_44/d_3_ DECAP_INV_G11
XG931 XI11_7/XI0/XI0_44/d__2_ XI11_7/XI0/XI0_44/d_2_ DECAP_INV_G11
XG932 XI11_7/XI0/XI0_44/d__1_ XI11_7/XI0/XI0_44/d_1_ DECAP_INV_G11
XG933 XI11_7/XI0/XI0_44/d__0_ XI11_7/XI0/XI0_44/d_0_ DECAP_INV_G11
XG934 XI11_7/XI0/XI0_44/d_15_ XI11_7/XI0/XI0_44/d__15_ DECAP_INV_G11
XG935 XI11_7/XI0/XI0_44/d_14_ XI11_7/XI0/XI0_44/d__14_ DECAP_INV_G11
XG936 XI11_7/XI0/XI0_44/d_13_ XI11_7/XI0/XI0_44/d__13_ DECAP_INV_G11
XG937 XI11_7/XI0/XI0_44/d_12_ XI11_7/XI0/XI0_44/d__12_ DECAP_INV_G11
XG938 XI11_7/XI0/XI0_44/d_11_ XI11_7/XI0/XI0_44/d__11_ DECAP_INV_G11
XG939 XI11_7/XI0/XI0_44/d_10_ XI11_7/XI0/XI0_44/d__10_ DECAP_INV_G11
XG940 XI11_7/XI0/XI0_44/d_9_ XI11_7/XI0/XI0_44/d__9_ DECAP_INV_G11
XG941 XI11_7/XI0/XI0_44/d_8_ XI11_7/XI0/XI0_44/d__8_ DECAP_INV_G11
XG942 XI11_7/XI0/XI0_44/d_7_ XI11_7/XI0/XI0_44/d__7_ DECAP_INV_G11
XG943 XI11_7/XI0/XI0_44/d_6_ XI11_7/XI0/XI0_44/d__6_ DECAP_INV_G11
XG944 XI11_7/XI0/XI0_44/d_5_ XI11_7/XI0/XI0_44/d__5_ DECAP_INV_G11
XG945 XI11_7/XI0/XI0_44/d_4_ XI11_7/XI0/XI0_44/d__4_ DECAP_INV_G11
XG946 XI11_7/XI0/XI0_44/d_3_ XI11_7/XI0/XI0_44/d__3_ DECAP_INV_G11
XG947 XI11_7/XI0/XI0_44/d_2_ XI11_7/XI0/XI0_44/d__2_ DECAP_INV_G11
XG948 XI11_7/XI0/XI0_44/d_1_ XI11_7/XI0/XI0_44/d__1_ DECAP_INV_G11
XG949 XI11_7/XI0/XI0_44/d_0_ XI11_7/XI0/XI0_44/d__0_ DECAP_INV_G11
XG950 XI11_7/XI0/XI0_43/d__15_ XI11_7/XI0/XI0_43/d_15_ DECAP_INV_G11
XG951 XI11_7/XI0/XI0_43/d__14_ XI11_7/XI0/XI0_43/d_14_ DECAP_INV_G11
XG952 XI11_7/XI0/XI0_43/d__13_ XI11_7/XI0/XI0_43/d_13_ DECAP_INV_G11
XG953 XI11_7/XI0/XI0_43/d__12_ XI11_7/XI0/XI0_43/d_12_ DECAP_INV_G11
XG954 XI11_7/XI0/XI0_43/d__11_ XI11_7/XI0/XI0_43/d_11_ DECAP_INV_G11
XG955 XI11_7/XI0/XI0_43/d__10_ XI11_7/XI0/XI0_43/d_10_ DECAP_INV_G11
XG956 XI11_7/XI0/XI0_43/d__9_ XI11_7/XI0/XI0_43/d_9_ DECAP_INV_G11
XG957 XI11_7/XI0/XI0_43/d__8_ XI11_7/XI0/XI0_43/d_8_ DECAP_INV_G11
XG958 XI11_7/XI0/XI0_43/d__7_ XI11_7/XI0/XI0_43/d_7_ DECAP_INV_G11
XG959 XI11_7/XI0/XI0_43/d__6_ XI11_7/XI0/XI0_43/d_6_ DECAP_INV_G11
XG960 XI11_7/XI0/XI0_43/d__5_ XI11_7/XI0/XI0_43/d_5_ DECAP_INV_G11
XG961 XI11_7/XI0/XI0_43/d__4_ XI11_7/XI0/XI0_43/d_4_ DECAP_INV_G11
XG962 XI11_7/XI0/XI0_43/d__3_ XI11_7/XI0/XI0_43/d_3_ DECAP_INV_G11
XG963 XI11_7/XI0/XI0_43/d__2_ XI11_7/XI0/XI0_43/d_2_ DECAP_INV_G11
XG964 XI11_7/XI0/XI0_43/d__1_ XI11_7/XI0/XI0_43/d_1_ DECAP_INV_G11
XG965 XI11_7/XI0/XI0_43/d__0_ XI11_7/XI0/XI0_43/d_0_ DECAP_INV_G11
XG966 XI11_7/XI0/XI0_43/d_15_ XI11_7/XI0/XI0_43/d__15_ DECAP_INV_G11
XG967 XI11_7/XI0/XI0_43/d_14_ XI11_7/XI0/XI0_43/d__14_ DECAP_INV_G11
XG968 XI11_7/XI0/XI0_43/d_13_ XI11_7/XI0/XI0_43/d__13_ DECAP_INV_G11
XG969 XI11_7/XI0/XI0_43/d_12_ XI11_7/XI0/XI0_43/d__12_ DECAP_INV_G11
XG970 XI11_7/XI0/XI0_43/d_11_ XI11_7/XI0/XI0_43/d__11_ DECAP_INV_G11
XG971 XI11_7/XI0/XI0_43/d_10_ XI11_7/XI0/XI0_43/d__10_ DECAP_INV_G11
XG972 XI11_7/XI0/XI0_43/d_9_ XI11_7/XI0/XI0_43/d__9_ DECAP_INV_G11
XG973 XI11_7/XI0/XI0_43/d_8_ XI11_7/XI0/XI0_43/d__8_ DECAP_INV_G11
XG974 XI11_7/XI0/XI0_43/d_7_ XI11_7/XI0/XI0_43/d__7_ DECAP_INV_G11
XG975 XI11_7/XI0/XI0_43/d_6_ XI11_7/XI0/XI0_43/d__6_ DECAP_INV_G11
XG976 XI11_7/XI0/XI0_43/d_5_ XI11_7/XI0/XI0_43/d__5_ DECAP_INV_G11
XG977 XI11_7/XI0/XI0_43/d_4_ XI11_7/XI0/XI0_43/d__4_ DECAP_INV_G11
XG978 XI11_7/XI0/XI0_43/d_3_ XI11_7/XI0/XI0_43/d__3_ DECAP_INV_G11
XG979 XI11_7/XI0/XI0_43/d_2_ XI11_7/XI0/XI0_43/d__2_ DECAP_INV_G11
XG980 XI11_7/XI0/XI0_43/d_1_ XI11_7/XI0/XI0_43/d__1_ DECAP_INV_G11
XG981 XI11_7/XI0/XI0_43/d_0_ XI11_7/XI0/XI0_43/d__0_ DECAP_INV_G11
XG982 XI11_7/XI0/XI0_42/d__15_ XI11_7/XI0/XI0_42/d_15_ DECAP_INV_G11
XG983 XI11_7/XI0/XI0_42/d__14_ XI11_7/XI0/XI0_42/d_14_ DECAP_INV_G11
XG984 XI11_7/XI0/XI0_42/d__13_ XI11_7/XI0/XI0_42/d_13_ DECAP_INV_G11
XG985 XI11_7/XI0/XI0_42/d__12_ XI11_7/XI0/XI0_42/d_12_ DECAP_INV_G11
XG986 XI11_7/XI0/XI0_42/d__11_ XI11_7/XI0/XI0_42/d_11_ DECAP_INV_G11
XG987 XI11_7/XI0/XI0_42/d__10_ XI11_7/XI0/XI0_42/d_10_ DECAP_INV_G11
XG988 XI11_7/XI0/XI0_42/d__9_ XI11_7/XI0/XI0_42/d_9_ DECAP_INV_G11
XG989 XI11_7/XI0/XI0_42/d__8_ XI11_7/XI0/XI0_42/d_8_ DECAP_INV_G11
XG990 XI11_7/XI0/XI0_42/d__7_ XI11_7/XI0/XI0_42/d_7_ DECAP_INV_G11
XG991 XI11_7/XI0/XI0_42/d__6_ XI11_7/XI0/XI0_42/d_6_ DECAP_INV_G11
XG992 XI11_7/XI0/XI0_42/d__5_ XI11_7/XI0/XI0_42/d_5_ DECAP_INV_G11
XG993 XI11_7/XI0/XI0_42/d__4_ XI11_7/XI0/XI0_42/d_4_ DECAP_INV_G11
XG994 XI11_7/XI0/XI0_42/d__3_ XI11_7/XI0/XI0_42/d_3_ DECAP_INV_G11
XG995 XI11_7/XI0/XI0_42/d__2_ XI11_7/XI0/XI0_42/d_2_ DECAP_INV_G11
XG996 XI11_7/XI0/XI0_42/d__1_ XI11_7/XI0/XI0_42/d_1_ DECAP_INV_G11
XG997 XI11_7/XI0/XI0_42/d__0_ XI11_7/XI0/XI0_42/d_0_ DECAP_INV_G11
XG998 XI11_7/XI0/XI0_42/d_15_ XI11_7/XI0/XI0_42/d__15_ DECAP_INV_G11
XG999 XI11_7/XI0/XI0_42/d_14_ XI11_7/XI0/XI0_42/d__14_ DECAP_INV_G11
XG1000 XI11_7/XI0/XI0_42/d_13_ XI11_7/XI0/XI0_42/d__13_ DECAP_INV_G11
XG1001 XI11_7/XI0/XI0_42/d_12_ XI11_7/XI0/XI0_42/d__12_ DECAP_INV_G11
XG1002 XI11_7/XI0/XI0_42/d_11_ XI11_7/XI0/XI0_42/d__11_ DECAP_INV_G11
XG1003 XI11_7/XI0/XI0_42/d_10_ XI11_7/XI0/XI0_42/d__10_ DECAP_INV_G11
XG1004 XI11_7/XI0/XI0_42/d_9_ XI11_7/XI0/XI0_42/d__9_ DECAP_INV_G11
XG1005 XI11_7/XI0/XI0_42/d_8_ XI11_7/XI0/XI0_42/d__8_ DECAP_INV_G11
XG1006 XI11_7/XI0/XI0_42/d_7_ XI11_7/XI0/XI0_42/d__7_ DECAP_INV_G11
XG1007 XI11_7/XI0/XI0_42/d_6_ XI11_7/XI0/XI0_42/d__6_ DECAP_INV_G11
XG1008 XI11_7/XI0/XI0_42/d_5_ XI11_7/XI0/XI0_42/d__5_ DECAP_INV_G11
XG1009 XI11_7/XI0/XI0_42/d_4_ XI11_7/XI0/XI0_42/d__4_ DECAP_INV_G11
XG1010 XI11_7/XI0/XI0_42/d_3_ XI11_7/XI0/XI0_42/d__3_ DECAP_INV_G11
XG1011 XI11_7/XI0/XI0_42/d_2_ XI11_7/XI0/XI0_42/d__2_ DECAP_INV_G11
XG1012 XI11_7/XI0/XI0_42/d_1_ XI11_7/XI0/XI0_42/d__1_ DECAP_INV_G11
XG1013 XI11_7/XI0/XI0_42/d_0_ XI11_7/XI0/XI0_42/d__0_ DECAP_INV_G11
XG1014 XI11_7/XI0/XI0_41/d__15_ XI11_7/XI0/XI0_41/d_15_ DECAP_INV_G11
XG1015 XI11_7/XI0/XI0_41/d__14_ XI11_7/XI0/XI0_41/d_14_ DECAP_INV_G11
XG1016 XI11_7/XI0/XI0_41/d__13_ XI11_7/XI0/XI0_41/d_13_ DECAP_INV_G11
XG1017 XI11_7/XI0/XI0_41/d__12_ XI11_7/XI0/XI0_41/d_12_ DECAP_INV_G11
XG1018 XI11_7/XI0/XI0_41/d__11_ XI11_7/XI0/XI0_41/d_11_ DECAP_INV_G11
XG1019 XI11_7/XI0/XI0_41/d__10_ XI11_7/XI0/XI0_41/d_10_ DECAP_INV_G11
XG1020 XI11_7/XI0/XI0_41/d__9_ XI11_7/XI0/XI0_41/d_9_ DECAP_INV_G11
XG1021 XI11_7/XI0/XI0_41/d__8_ XI11_7/XI0/XI0_41/d_8_ DECAP_INV_G11
XG1022 XI11_7/XI0/XI0_41/d__7_ XI11_7/XI0/XI0_41/d_7_ DECAP_INV_G11
XG1023 XI11_7/XI0/XI0_41/d__6_ XI11_7/XI0/XI0_41/d_6_ DECAP_INV_G11
XG1024 XI11_7/XI0/XI0_41/d__5_ XI11_7/XI0/XI0_41/d_5_ DECAP_INV_G11
XG1025 XI11_7/XI0/XI0_41/d__4_ XI11_7/XI0/XI0_41/d_4_ DECAP_INV_G11
XG1026 XI11_7/XI0/XI0_41/d__3_ XI11_7/XI0/XI0_41/d_3_ DECAP_INV_G11
XG1027 XI11_7/XI0/XI0_41/d__2_ XI11_7/XI0/XI0_41/d_2_ DECAP_INV_G11
XG1028 XI11_7/XI0/XI0_41/d__1_ XI11_7/XI0/XI0_41/d_1_ DECAP_INV_G11
XG1029 XI11_7/XI0/XI0_41/d__0_ XI11_7/XI0/XI0_41/d_0_ DECAP_INV_G11
XG1030 XI11_7/XI0/XI0_41/d_15_ XI11_7/XI0/XI0_41/d__15_ DECAP_INV_G11
XG1031 XI11_7/XI0/XI0_41/d_14_ XI11_7/XI0/XI0_41/d__14_ DECAP_INV_G11
XG1032 XI11_7/XI0/XI0_41/d_13_ XI11_7/XI0/XI0_41/d__13_ DECAP_INV_G11
XG1033 XI11_7/XI0/XI0_41/d_12_ XI11_7/XI0/XI0_41/d__12_ DECAP_INV_G11
XG1034 XI11_7/XI0/XI0_41/d_11_ XI11_7/XI0/XI0_41/d__11_ DECAP_INV_G11
XG1035 XI11_7/XI0/XI0_41/d_10_ XI11_7/XI0/XI0_41/d__10_ DECAP_INV_G11
XG1036 XI11_7/XI0/XI0_41/d_9_ XI11_7/XI0/XI0_41/d__9_ DECAP_INV_G11
XG1037 XI11_7/XI0/XI0_41/d_8_ XI11_7/XI0/XI0_41/d__8_ DECAP_INV_G11
XG1038 XI11_7/XI0/XI0_41/d_7_ XI11_7/XI0/XI0_41/d__7_ DECAP_INV_G11
XG1039 XI11_7/XI0/XI0_41/d_6_ XI11_7/XI0/XI0_41/d__6_ DECAP_INV_G11
XG1040 XI11_7/XI0/XI0_41/d_5_ XI11_7/XI0/XI0_41/d__5_ DECAP_INV_G11
XG1041 XI11_7/XI0/XI0_41/d_4_ XI11_7/XI0/XI0_41/d__4_ DECAP_INV_G11
XG1042 XI11_7/XI0/XI0_41/d_3_ XI11_7/XI0/XI0_41/d__3_ DECAP_INV_G11
XG1043 XI11_7/XI0/XI0_41/d_2_ XI11_7/XI0/XI0_41/d__2_ DECAP_INV_G11
XG1044 XI11_7/XI0/XI0_41/d_1_ XI11_7/XI0/XI0_41/d__1_ DECAP_INV_G11
XG1045 XI11_7/XI0/XI0_41/d_0_ XI11_7/XI0/XI0_41/d__0_ DECAP_INV_G11
XG1046 XI11_7/XI0/XI0_40/d__15_ XI11_7/XI0/XI0_40/d_15_ DECAP_INV_G11
XG1047 XI11_7/XI0/XI0_40/d__14_ XI11_7/XI0/XI0_40/d_14_ DECAP_INV_G11
XG1048 XI11_7/XI0/XI0_40/d__13_ XI11_7/XI0/XI0_40/d_13_ DECAP_INV_G11
XG1049 XI11_7/XI0/XI0_40/d__12_ XI11_7/XI0/XI0_40/d_12_ DECAP_INV_G11
XG1050 XI11_7/XI0/XI0_40/d__11_ XI11_7/XI0/XI0_40/d_11_ DECAP_INV_G11
XG1051 XI11_7/XI0/XI0_40/d__10_ XI11_7/XI0/XI0_40/d_10_ DECAP_INV_G11
XG1052 XI11_7/XI0/XI0_40/d__9_ XI11_7/XI0/XI0_40/d_9_ DECAP_INV_G11
XG1053 XI11_7/XI0/XI0_40/d__8_ XI11_7/XI0/XI0_40/d_8_ DECAP_INV_G11
XG1054 XI11_7/XI0/XI0_40/d__7_ XI11_7/XI0/XI0_40/d_7_ DECAP_INV_G11
XG1055 XI11_7/XI0/XI0_40/d__6_ XI11_7/XI0/XI0_40/d_6_ DECAP_INV_G11
XG1056 XI11_7/XI0/XI0_40/d__5_ XI11_7/XI0/XI0_40/d_5_ DECAP_INV_G11
XG1057 XI11_7/XI0/XI0_40/d__4_ XI11_7/XI0/XI0_40/d_4_ DECAP_INV_G11
XG1058 XI11_7/XI0/XI0_40/d__3_ XI11_7/XI0/XI0_40/d_3_ DECAP_INV_G11
XG1059 XI11_7/XI0/XI0_40/d__2_ XI11_7/XI0/XI0_40/d_2_ DECAP_INV_G11
XG1060 XI11_7/XI0/XI0_40/d__1_ XI11_7/XI0/XI0_40/d_1_ DECAP_INV_G11
XG1061 XI11_7/XI0/XI0_40/d__0_ XI11_7/XI0/XI0_40/d_0_ DECAP_INV_G11
XG1062 XI11_7/XI0/XI0_40/d_15_ XI11_7/XI0/XI0_40/d__15_ DECAP_INV_G11
XG1063 XI11_7/XI0/XI0_40/d_14_ XI11_7/XI0/XI0_40/d__14_ DECAP_INV_G11
XG1064 XI11_7/XI0/XI0_40/d_13_ XI11_7/XI0/XI0_40/d__13_ DECAP_INV_G11
XG1065 XI11_7/XI0/XI0_40/d_12_ XI11_7/XI0/XI0_40/d__12_ DECAP_INV_G11
XG1066 XI11_7/XI0/XI0_40/d_11_ XI11_7/XI0/XI0_40/d__11_ DECAP_INV_G11
XG1067 XI11_7/XI0/XI0_40/d_10_ XI11_7/XI0/XI0_40/d__10_ DECAP_INV_G11
XG1068 XI11_7/XI0/XI0_40/d_9_ XI11_7/XI0/XI0_40/d__9_ DECAP_INV_G11
XG1069 XI11_7/XI0/XI0_40/d_8_ XI11_7/XI0/XI0_40/d__8_ DECAP_INV_G11
XG1070 XI11_7/XI0/XI0_40/d_7_ XI11_7/XI0/XI0_40/d__7_ DECAP_INV_G11
XG1071 XI11_7/XI0/XI0_40/d_6_ XI11_7/XI0/XI0_40/d__6_ DECAP_INV_G11
XG1072 XI11_7/XI0/XI0_40/d_5_ XI11_7/XI0/XI0_40/d__5_ DECAP_INV_G11
XG1073 XI11_7/XI0/XI0_40/d_4_ XI11_7/XI0/XI0_40/d__4_ DECAP_INV_G11
XG1074 XI11_7/XI0/XI0_40/d_3_ XI11_7/XI0/XI0_40/d__3_ DECAP_INV_G11
XG1075 XI11_7/XI0/XI0_40/d_2_ XI11_7/XI0/XI0_40/d__2_ DECAP_INV_G11
XG1076 XI11_7/XI0/XI0_40/d_1_ XI11_7/XI0/XI0_40/d__1_ DECAP_INV_G11
XG1077 XI11_7/XI0/XI0_40/d_0_ XI11_7/XI0/XI0_40/d__0_ DECAP_INV_G11
XG1078 XI11_7/XI0/XI0_39/d__15_ XI11_7/XI0/XI0_39/d_15_ DECAP_INV_G11
XG1079 XI11_7/XI0/XI0_39/d__14_ XI11_7/XI0/XI0_39/d_14_ DECAP_INV_G11
XG1080 XI11_7/XI0/XI0_39/d__13_ XI11_7/XI0/XI0_39/d_13_ DECAP_INV_G11
XG1081 XI11_7/XI0/XI0_39/d__12_ XI11_7/XI0/XI0_39/d_12_ DECAP_INV_G11
XG1082 XI11_7/XI0/XI0_39/d__11_ XI11_7/XI0/XI0_39/d_11_ DECAP_INV_G11
XG1083 XI11_7/XI0/XI0_39/d__10_ XI11_7/XI0/XI0_39/d_10_ DECAP_INV_G11
XG1084 XI11_7/XI0/XI0_39/d__9_ XI11_7/XI0/XI0_39/d_9_ DECAP_INV_G11
XG1085 XI11_7/XI0/XI0_39/d__8_ XI11_7/XI0/XI0_39/d_8_ DECAP_INV_G11
XG1086 XI11_7/XI0/XI0_39/d__7_ XI11_7/XI0/XI0_39/d_7_ DECAP_INV_G11
XG1087 XI11_7/XI0/XI0_39/d__6_ XI11_7/XI0/XI0_39/d_6_ DECAP_INV_G11
XG1088 XI11_7/XI0/XI0_39/d__5_ XI11_7/XI0/XI0_39/d_5_ DECAP_INV_G11
XG1089 XI11_7/XI0/XI0_39/d__4_ XI11_7/XI0/XI0_39/d_4_ DECAP_INV_G11
XG1090 XI11_7/XI0/XI0_39/d__3_ XI11_7/XI0/XI0_39/d_3_ DECAP_INV_G11
XG1091 XI11_7/XI0/XI0_39/d__2_ XI11_7/XI0/XI0_39/d_2_ DECAP_INV_G11
XG1092 XI11_7/XI0/XI0_39/d__1_ XI11_7/XI0/XI0_39/d_1_ DECAP_INV_G11
XG1093 XI11_7/XI0/XI0_39/d__0_ XI11_7/XI0/XI0_39/d_0_ DECAP_INV_G11
XG1094 XI11_7/XI0/XI0_39/d_15_ XI11_7/XI0/XI0_39/d__15_ DECAP_INV_G11
XG1095 XI11_7/XI0/XI0_39/d_14_ XI11_7/XI0/XI0_39/d__14_ DECAP_INV_G11
XG1096 XI11_7/XI0/XI0_39/d_13_ XI11_7/XI0/XI0_39/d__13_ DECAP_INV_G11
XG1097 XI11_7/XI0/XI0_39/d_12_ XI11_7/XI0/XI0_39/d__12_ DECAP_INV_G11
XG1098 XI11_7/XI0/XI0_39/d_11_ XI11_7/XI0/XI0_39/d__11_ DECAP_INV_G11
XG1099 XI11_7/XI0/XI0_39/d_10_ XI11_7/XI0/XI0_39/d__10_ DECAP_INV_G11
XG1100 XI11_7/XI0/XI0_39/d_9_ XI11_7/XI0/XI0_39/d__9_ DECAP_INV_G11
XG1101 XI11_7/XI0/XI0_39/d_8_ XI11_7/XI0/XI0_39/d__8_ DECAP_INV_G11
XG1102 XI11_7/XI0/XI0_39/d_7_ XI11_7/XI0/XI0_39/d__7_ DECAP_INV_G11
XG1103 XI11_7/XI0/XI0_39/d_6_ XI11_7/XI0/XI0_39/d__6_ DECAP_INV_G11
XG1104 XI11_7/XI0/XI0_39/d_5_ XI11_7/XI0/XI0_39/d__5_ DECAP_INV_G11
XG1105 XI11_7/XI0/XI0_39/d_4_ XI11_7/XI0/XI0_39/d__4_ DECAP_INV_G11
XG1106 XI11_7/XI0/XI0_39/d_3_ XI11_7/XI0/XI0_39/d__3_ DECAP_INV_G11
XG1107 XI11_7/XI0/XI0_39/d_2_ XI11_7/XI0/XI0_39/d__2_ DECAP_INV_G11
XG1108 XI11_7/XI0/XI0_39/d_1_ XI11_7/XI0/XI0_39/d__1_ DECAP_INV_G11
XG1109 XI11_7/XI0/XI0_39/d_0_ XI11_7/XI0/XI0_39/d__0_ DECAP_INV_G11
XG1110 XI11_7/XI0/XI0_38/d__15_ XI11_7/XI0/XI0_38/d_15_ DECAP_INV_G11
XG1111 XI11_7/XI0/XI0_38/d__14_ XI11_7/XI0/XI0_38/d_14_ DECAP_INV_G11
XG1112 XI11_7/XI0/XI0_38/d__13_ XI11_7/XI0/XI0_38/d_13_ DECAP_INV_G11
XG1113 XI11_7/XI0/XI0_38/d__12_ XI11_7/XI0/XI0_38/d_12_ DECAP_INV_G11
XG1114 XI11_7/XI0/XI0_38/d__11_ XI11_7/XI0/XI0_38/d_11_ DECAP_INV_G11
XG1115 XI11_7/XI0/XI0_38/d__10_ XI11_7/XI0/XI0_38/d_10_ DECAP_INV_G11
XG1116 XI11_7/XI0/XI0_38/d__9_ XI11_7/XI0/XI0_38/d_9_ DECAP_INV_G11
XG1117 XI11_7/XI0/XI0_38/d__8_ XI11_7/XI0/XI0_38/d_8_ DECAP_INV_G11
XG1118 XI11_7/XI0/XI0_38/d__7_ XI11_7/XI0/XI0_38/d_7_ DECAP_INV_G11
XG1119 XI11_7/XI0/XI0_38/d__6_ XI11_7/XI0/XI0_38/d_6_ DECAP_INV_G11
XG1120 XI11_7/XI0/XI0_38/d__5_ XI11_7/XI0/XI0_38/d_5_ DECAP_INV_G11
XG1121 XI11_7/XI0/XI0_38/d__4_ XI11_7/XI0/XI0_38/d_4_ DECAP_INV_G11
XG1122 XI11_7/XI0/XI0_38/d__3_ XI11_7/XI0/XI0_38/d_3_ DECAP_INV_G11
XG1123 XI11_7/XI0/XI0_38/d__2_ XI11_7/XI0/XI0_38/d_2_ DECAP_INV_G11
XG1124 XI11_7/XI0/XI0_38/d__1_ XI11_7/XI0/XI0_38/d_1_ DECAP_INV_G11
XG1125 XI11_7/XI0/XI0_38/d__0_ XI11_7/XI0/XI0_38/d_0_ DECAP_INV_G11
XG1126 XI11_7/XI0/XI0_38/d_15_ XI11_7/XI0/XI0_38/d__15_ DECAP_INV_G11
XG1127 XI11_7/XI0/XI0_38/d_14_ XI11_7/XI0/XI0_38/d__14_ DECAP_INV_G11
XG1128 XI11_7/XI0/XI0_38/d_13_ XI11_7/XI0/XI0_38/d__13_ DECAP_INV_G11
XG1129 XI11_7/XI0/XI0_38/d_12_ XI11_7/XI0/XI0_38/d__12_ DECAP_INV_G11
XG1130 XI11_7/XI0/XI0_38/d_11_ XI11_7/XI0/XI0_38/d__11_ DECAP_INV_G11
XG1131 XI11_7/XI0/XI0_38/d_10_ XI11_7/XI0/XI0_38/d__10_ DECAP_INV_G11
XG1132 XI11_7/XI0/XI0_38/d_9_ XI11_7/XI0/XI0_38/d__9_ DECAP_INV_G11
XG1133 XI11_7/XI0/XI0_38/d_8_ XI11_7/XI0/XI0_38/d__8_ DECAP_INV_G11
XG1134 XI11_7/XI0/XI0_38/d_7_ XI11_7/XI0/XI0_38/d__7_ DECAP_INV_G11
XG1135 XI11_7/XI0/XI0_38/d_6_ XI11_7/XI0/XI0_38/d__6_ DECAP_INV_G11
XG1136 XI11_7/XI0/XI0_38/d_5_ XI11_7/XI0/XI0_38/d__5_ DECAP_INV_G11
XG1137 XI11_7/XI0/XI0_38/d_4_ XI11_7/XI0/XI0_38/d__4_ DECAP_INV_G11
XG1138 XI11_7/XI0/XI0_38/d_3_ XI11_7/XI0/XI0_38/d__3_ DECAP_INV_G11
XG1139 XI11_7/XI0/XI0_38/d_2_ XI11_7/XI0/XI0_38/d__2_ DECAP_INV_G11
XG1140 XI11_7/XI0/XI0_38/d_1_ XI11_7/XI0/XI0_38/d__1_ DECAP_INV_G11
XG1141 XI11_7/XI0/XI0_38/d_0_ XI11_7/XI0/XI0_38/d__0_ DECAP_INV_G11
XG1142 XI11_7/XI0/XI0_37/d__15_ XI11_7/XI0/XI0_37/d_15_ DECAP_INV_G11
XG1143 XI11_7/XI0/XI0_37/d__14_ XI11_7/XI0/XI0_37/d_14_ DECAP_INV_G11
XG1144 XI11_7/XI0/XI0_37/d__13_ XI11_7/XI0/XI0_37/d_13_ DECAP_INV_G11
XG1145 XI11_7/XI0/XI0_37/d__12_ XI11_7/XI0/XI0_37/d_12_ DECAP_INV_G11
XG1146 XI11_7/XI0/XI0_37/d__11_ XI11_7/XI0/XI0_37/d_11_ DECAP_INV_G11
XG1147 XI11_7/XI0/XI0_37/d__10_ XI11_7/XI0/XI0_37/d_10_ DECAP_INV_G11
XG1148 XI11_7/XI0/XI0_37/d__9_ XI11_7/XI0/XI0_37/d_9_ DECAP_INV_G11
XG1149 XI11_7/XI0/XI0_37/d__8_ XI11_7/XI0/XI0_37/d_8_ DECAP_INV_G11
XG1150 XI11_7/XI0/XI0_37/d__7_ XI11_7/XI0/XI0_37/d_7_ DECAP_INV_G11
XG1151 XI11_7/XI0/XI0_37/d__6_ XI11_7/XI0/XI0_37/d_6_ DECAP_INV_G11
XG1152 XI11_7/XI0/XI0_37/d__5_ XI11_7/XI0/XI0_37/d_5_ DECAP_INV_G11
XG1153 XI11_7/XI0/XI0_37/d__4_ XI11_7/XI0/XI0_37/d_4_ DECAP_INV_G11
XG1154 XI11_7/XI0/XI0_37/d__3_ XI11_7/XI0/XI0_37/d_3_ DECAP_INV_G11
XG1155 XI11_7/XI0/XI0_37/d__2_ XI11_7/XI0/XI0_37/d_2_ DECAP_INV_G11
XG1156 XI11_7/XI0/XI0_37/d__1_ XI11_7/XI0/XI0_37/d_1_ DECAP_INV_G11
XG1157 XI11_7/XI0/XI0_37/d__0_ XI11_7/XI0/XI0_37/d_0_ DECAP_INV_G11
XG1158 XI11_7/XI0/XI0_37/d_15_ XI11_7/XI0/XI0_37/d__15_ DECAP_INV_G11
XG1159 XI11_7/XI0/XI0_37/d_14_ XI11_7/XI0/XI0_37/d__14_ DECAP_INV_G11
XG1160 XI11_7/XI0/XI0_37/d_13_ XI11_7/XI0/XI0_37/d__13_ DECAP_INV_G11
XG1161 XI11_7/XI0/XI0_37/d_12_ XI11_7/XI0/XI0_37/d__12_ DECAP_INV_G11
XG1162 XI11_7/XI0/XI0_37/d_11_ XI11_7/XI0/XI0_37/d__11_ DECAP_INV_G11
XG1163 XI11_7/XI0/XI0_37/d_10_ XI11_7/XI0/XI0_37/d__10_ DECAP_INV_G11
XG1164 XI11_7/XI0/XI0_37/d_9_ XI11_7/XI0/XI0_37/d__9_ DECAP_INV_G11
XG1165 XI11_7/XI0/XI0_37/d_8_ XI11_7/XI0/XI0_37/d__8_ DECAP_INV_G11
XG1166 XI11_7/XI0/XI0_37/d_7_ XI11_7/XI0/XI0_37/d__7_ DECAP_INV_G11
XG1167 XI11_7/XI0/XI0_37/d_6_ XI11_7/XI0/XI0_37/d__6_ DECAP_INV_G11
XG1168 XI11_7/XI0/XI0_37/d_5_ XI11_7/XI0/XI0_37/d__5_ DECAP_INV_G11
XG1169 XI11_7/XI0/XI0_37/d_4_ XI11_7/XI0/XI0_37/d__4_ DECAP_INV_G11
XG1170 XI11_7/XI0/XI0_37/d_3_ XI11_7/XI0/XI0_37/d__3_ DECAP_INV_G11
XG1171 XI11_7/XI0/XI0_37/d_2_ XI11_7/XI0/XI0_37/d__2_ DECAP_INV_G11
XG1172 XI11_7/XI0/XI0_37/d_1_ XI11_7/XI0/XI0_37/d__1_ DECAP_INV_G11
XG1173 XI11_7/XI0/XI0_37/d_0_ XI11_7/XI0/XI0_37/d__0_ DECAP_INV_G11
XG1174 XI11_7/XI0/XI0_36/d__15_ XI11_7/XI0/XI0_36/d_15_ DECAP_INV_G11
XG1175 XI11_7/XI0/XI0_36/d__14_ XI11_7/XI0/XI0_36/d_14_ DECAP_INV_G11
XG1176 XI11_7/XI0/XI0_36/d__13_ XI11_7/XI0/XI0_36/d_13_ DECAP_INV_G11
XG1177 XI11_7/XI0/XI0_36/d__12_ XI11_7/XI0/XI0_36/d_12_ DECAP_INV_G11
XG1178 XI11_7/XI0/XI0_36/d__11_ XI11_7/XI0/XI0_36/d_11_ DECAP_INV_G11
XG1179 XI11_7/XI0/XI0_36/d__10_ XI11_7/XI0/XI0_36/d_10_ DECAP_INV_G11
XG1180 XI11_7/XI0/XI0_36/d__9_ XI11_7/XI0/XI0_36/d_9_ DECAP_INV_G11
XG1181 XI11_7/XI0/XI0_36/d__8_ XI11_7/XI0/XI0_36/d_8_ DECAP_INV_G11
XG1182 XI11_7/XI0/XI0_36/d__7_ XI11_7/XI0/XI0_36/d_7_ DECAP_INV_G11
XG1183 XI11_7/XI0/XI0_36/d__6_ XI11_7/XI0/XI0_36/d_6_ DECAP_INV_G11
XG1184 XI11_7/XI0/XI0_36/d__5_ XI11_7/XI0/XI0_36/d_5_ DECAP_INV_G11
XG1185 XI11_7/XI0/XI0_36/d__4_ XI11_7/XI0/XI0_36/d_4_ DECAP_INV_G11
XG1186 XI11_7/XI0/XI0_36/d__3_ XI11_7/XI0/XI0_36/d_3_ DECAP_INV_G11
XG1187 XI11_7/XI0/XI0_36/d__2_ XI11_7/XI0/XI0_36/d_2_ DECAP_INV_G11
XG1188 XI11_7/XI0/XI0_36/d__1_ XI11_7/XI0/XI0_36/d_1_ DECAP_INV_G11
XG1189 XI11_7/XI0/XI0_36/d__0_ XI11_7/XI0/XI0_36/d_0_ DECAP_INV_G11
XG1190 XI11_7/XI0/XI0_36/d_15_ XI11_7/XI0/XI0_36/d__15_ DECAP_INV_G11
XG1191 XI11_7/XI0/XI0_36/d_14_ XI11_7/XI0/XI0_36/d__14_ DECAP_INV_G11
XG1192 XI11_7/XI0/XI0_36/d_13_ XI11_7/XI0/XI0_36/d__13_ DECAP_INV_G11
XG1193 XI11_7/XI0/XI0_36/d_12_ XI11_7/XI0/XI0_36/d__12_ DECAP_INV_G11
XG1194 XI11_7/XI0/XI0_36/d_11_ XI11_7/XI0/XI0_36/d__11_ DECAP_INV_G11
XG1195 XI11_7/XI0/XI0_36/d_10_ XI11_7/XI0/XI0_36/d__10_ DECAP_INV_G11
XG1196 XI11_7/XI0/XI0_36/d_9_ XI11_7/XI0/XI0_36/d__9_ DECAP_INV_G11
XG1197 XI11_7/XI0/XI0_36/d_8_ XI11_7/XI0/XI0_36/d__8_ DECAP_INV_G11
XG1198 XI11_7/XI0/XI0_36/d_7_ XI11_7/XI0/XI0_36/d__7_ DECAP_INV_G11
XG1199 XI11_7/XI0/XI0_36/d_6_ XI11_7/XI0/XI0_36/d__6_ DECAP_INV_G11
XG1200 XI11_7/XI0/XI0_36/d_5_ XI11_7/XI0/XI0_36/d__5_ DECAP_INV_G11
XG1201 XI11_7/XI0/XI0_36/d_4_ XI11_7/XI0/XI0_36/d__4_ DECAP_INV_G11
XG1202 XI11_7/XI0/XI0_36/d_3_ XI11_7/XI0/XI0_36/d__3_ DECAP_INV_G11
XG1203 XI11_7/XI0/XI0_36/d_2_ XI11_7/XI0/XI0_36/d__2_ DECAP_INV_G11
XG1204 XI11_7/XI0/XI0_36/d_1_ XI11_7/XI0/XI0_36/d__1_ DECAP_INV_G11
XG1205 XI11_7/XI0/XI0_36/d_0_ XI11_7/XI0/XI0_36/d__0_ DECAP_INV_G11
XG1206 XI11_7/XI0/XI0_35/d__15_ XI11_7/XI0/XI0_35/d_15_ DECAP_INV_G11
XG1207 XI11_7/XI0/XI0_35/d__14_ XI11_7/XI0/XI0_35/d_14_ DECAP_INV_G11
XG1208 XI11_7/XI0/XI0_35/d__13_ XI11_7/XI0/XI0_35/d_13_ DECAP_INV_G11
XG1209 XI11_7/XI0/XI0_35/d__12_ XI11_7/XI0/XI0_35/d_12_ DECAP_INV_G11
XG1210 XI11_7/XI0/XI0_35/d__11_ XI11_7/XI0/XI0_35/d_11_ DECAP_INV_G11
XG1211 XI11_7/XI0/XI0_35/d__10_ XI11_7/XI0/XI0_35/d_10_ DECAP_INV_G11
XG1212 XI11_7/XI0/XI0_35/d__9_ XI11_7/XI0/XI0_35/d_9_ DECAP_INV_G11
XG1213 XI11_7/XI0/XI0_35/d__8_ XI11_7/XI0/XI0_35/d_8_ DECAP_INV_G11
XG1214 XI11_7/XI0/XI0_35/d__7_ XI11_7/XI0/XI0_35/d_7_ DECAP_INV_G11
XG1215 XI11_7/XI0/XI0_35/d__6_ XI11_7/XI0/XI0_35/d_6_ DECAP_INV_G11
XG1216 XI11_7/XI0/XI0_35/d__5_ XI11_7/XI0/XI0_35/d_5_ DECAP_INV_G11
XG1217 XI11_7/XI0/XI0_35/d__4_ XI11_7/XI0/XI0_35/d_4_ DECAP_INV_G11
XG1218 XI11_7/XI0/XI0_35/d__3_ XI11_7/XI0/XI0_35/d_3_ DECAP_INV_G11
XG1219 XI11_7/XI0/XI0_35/d__2_ XI11_7/XI0/XI0_35/d_2_ DECAP_INV_G11
XG1220 XI11_7/XI0/XI0_35/d__1_ XI11_7/XI0/XI0_35/d_1_ DECAP_INV_G11
XG1221 XI11_7/XI0/XI0_35/d__0_ XI11_7/XI0/XI0_35/d_0_ DECAP_INV_G11
XG1222 XI11_7/XI0/XI0_35/d_15_ XI11_7/XI0/XI0_35/d__15_ DECAP_INV_G11
XG1223 XI11_7/XI0/XI0_35/d_14_ XI11_7/XI0/XI0_35/d__14_ DECAP_INV_G11
XG1224 XI11_7/XI0/XI0_35/d_13_ XI11_7/XI0/XI0_35/d__13_ DECAP_INV_G11
XG1225 XI11_7/XI0/XI0_35/d_12_ XI11_7/XI0/XI0_35/d__12_ DECAP_INV_G11
XG1226 XI11_7/XI0/XI0_35/d_11_ XI11_7/XI0/XI0_35/d__11_ DECAP_INV_G11
XG1227 XI11_7/XI0/XI0_35/d_10_ XI11_7/XI0/XI0_35/d__10_ DECAP_INV_G11
XG1228 XI11_7/XI0/XI0_35/d_9_ XI11_7/XI0/XI0_35/d__9_ DECAP_INV_G11
XG1229 XI11_7/XI0/XI0_35/d_8_ XI11_7/XI0/XI0_35/d__8_ DECAP_INV_G11
XG1230 XI11_7/XI0/XI0_35/d_7_ XI11_7/XI0/XI0_35/d__7_ DECAP_INV_G11
XG1231 XI11_7/XI0/XI0_35/d_6_ XI11_7/XI0/XI0_35/d__6_ DECAP_INV_G11
XG1232 XI11_7/XI0/XI0_35/d_5_ XI11_7/XI0/XI0_35/d__5_ DECAP_INV_G11
XG1233 XI11_7/XI0/XI0_35/d_4_ XI11_7/XI0/XI0_35/d__4_ DECAP_INV_G11
XG1234 XI11_7/XI0/XI0_35/d_3_ XI11_7/XI0/XI0_35/d__3_ DECAP_INV_G11
XG1235 XI11_7/XI0/XI0_35/d_2_ XI11_7/XI0/XI0_35/d__2_ DECAP_INV_G11
XG1236 XI11_7/XI0/XI0_35/d_1_ XI11_7/XI0/XI0_35/d__1_ DECAP_INV_G11
XG1237 XI11_7/XI0/XI0_35/d_0_ XI11_7/XI0/XI0_35/d__0_ DECAP_INV_G11
XG1238 XI11_7/XI0/XI0_34/d__15_ XI11_7/XI0/XI0_34/d_15_ DECAP_INV_G11
XG1239 XI11_7/XI0/XI0_34/d__14_ XI11_7/XI0/XI0_34/d_14_ DECAP_INV_G11
XG1240 XI11_7/XI0/XI0_34/d__13_ XI11_7/XI0/XI0_34/d_13_ DECAP_INV_G11
XG1241 XI11_7/XI0/XI0_34/d__12_ XI11_7/XI0/XI0_34/d_12_ DECAP_INV_G11
XG1242 XI11_7/XI0/XI0_34/d__11_ XI11_7/XI0/XI0_34/d_11_ DECAP_INV_G11
XG1243 XI11_7/XI0/XI0_34/d__10_ XI11_7/XI0/XI0_34/d_10_ DECAP_INV_G11
XG1244 XI11_7/XI0/XI0_34/d__9_ XI11_7/XI0/XI0_34/d_9_ DECAP_INV_G11
XG1245 XI11_7/XI0/XI0_34/d__8_ XI11_7/XI0/XI0_34/d_8_ DECAP_INV_G11
XG1246 XI11_7/XI0/XI0_34/d__7_ XI11_7/XI0/XI0_34/d_7_ DECAP_INV_G11
XG1247 XI11_7/XI0/XI0_34/d__6_ XI11_7/XI0/XI0_34/d_6_ DECAP_INV_G11
XG1248 XI11_7/XI0/XI0_34/d__5_ XI11_7/XI0/XI0_34/d_5_ DECAP_INV_G11
XG1249 XI11_7/XI0/XI0_34/d__4_ XI11_7/XI0/XI0_34/d_4_ DECAP_INV_G11
XG1250 XI11_7/XI0/XI0_34/d__3_ XI11_7/XI0/XI0_34/d_3_ DECAP_INV_G11
XG1251 XI11_7/XI0/XI0_34/d__2_ XI11_7/XI0/XI0_34/d_2_ DECAP_INV_G11
XG1252 XI11_7/XI0/XI0_34/d__1_ XI11_7/XI0/XI0_34/d_1_ DECAP_INV_G11
XG1253 XI11_7/XI0/XI0_34/d__0_ XI11_7/XI0/XI0_34/d_0_ DECAP_INV_G11
XG1254 XI11_7/XI0/XI0_34/d_15_ XI11_7/XI0/XI0_34/d__15_ DECAP_INV_G11
XG1255 XI11_7/XI0/XI0_34/d_14_ XI11_7/XI0/XI0_34/d__14_ DECAP_INV_G11
XG1256 XI11_7/XI0/XI0_34/d_13_ XI11_7/XI0/XI0_34/d__13_ DECAP_INV_G11
XG1257 XI11_7/XI0/XI0_34/d_12_ XI11_7/XI0/XI0_34/d__12_ DECAP_INV_G11
XG1258 XI11_7/XI0/XI0_34/d_11_ XI11_7/XI0/XI0_34/d__11_ DECAP_INV_G11
XG1259 XI11_7/XI0/XI0_34/d_10_ XI11_7/XI0/XI0_34/d__10_ DECAP_INV_G11
XG1260 XI11_7/XI0/XI0_34/d_9_ XI11_7/XI0/XI0_34/d__9_ DECAP_INV_G11
XG1261 XI11_7/XI0/XI0_34/d_8_ XI11_7/XI0/XI0_34/d__8_ DECAP_INV_G11
XG1262 XI11_7/XI0/XI0_34/d_7_ XI11_7/XI0/XI0_34/d__7_ DECAP_INV_G11
XG1263 XI11_7/XI0/XI0_34/d_6_ XI11_7/XI0/XI0_34/d__6_ DECAP_INV_G11
XG1264 XI11_7/XI0/XI0_34/d_5_ XI11_7/XI0/XI0_34/d__5_ DECAP_INV_G11
XG1265 XI11_7/XI0/XI0_34/d_4_ XI11_7/XI0/XI0_34/d__4_ DECAP_INV_G11
XG1266 XI11_7/XI0/XI0_34/d_3_ XI11_7/XI0/XI0_34/d__3_ DECAP_INV_G11
XG1267 XI11_7/XI0/XI0_34/d_2_ XI11_7/XI0/XI0_34/d__2_ DECAP_INV_G11
XG1268 XI11_7/XI0/XI0_34/d_1_ XI11_7/XI0/XI0_34/d__1_ DECAP_INV_G11
XG1269 XI11_7/XI0/XI0_34/d_0_ XI11_7/XI0/XI0_34/d__0_ DECAP_INV_G11
XG1270 XI11_7/XI0/XI0_33/d__15_ XI11_7/XI0/XI0_33/d_15_ DECAP_INV_G11
XG1271 XI11_7/XI0/XI0_33/d__14_ XI11_7/XI0/XI0_33/d_14_ DECAP_INV_G11
XG1272 XI11_7/XI0/XI0_33/d__13_ XI11_7/XI0/XI0_33/d_13_ DECAP_INV_G11
XG1273 XI11_7/XI0/XI0_33/d__12_ XI11_7/XI0/XI0_33/d_12_ DECAP_INV_G11
XG1274 XI11_7/XI0/XI0_33/d__11_ XI11_7/XI0/XI0_33/d_11_ DECAP_INV_G11
XG1275 XI11_7/XI0/XI0_33/d__10_ XI11_7/XI0/XI0_33/d_10_ DECAP_INV_G11
XG1276 XI11_7/XI0/XI0_33/d__9_ XI11_7/XI0/XI0_33/d_9_ DECAP_INV_G11
XG1277 XI11_7/XI0/XI0_33/d__8_ XI11_7/XI0/XI0_33/d_8_ DECAP_INV_G11
XG1278 XI11_7/XI0/XI0_33/d__7_ XI11_7/XI0/XI0_33/d_7_ DECAP_INV_G11
XG1279 XI11_7/XI0/XI0_33/d__6_ XI11_7/XI0/XI0_33/d_6_ DECAP_INV_G11
XG1280 XI11_7/XI0/XI0_33/d__5_ XI11_7/XI0/XI0_33/d_5_ DECAP_INV_G11
XG1281 XI11_7/XI0/XI0_33/d__4_ XI11_7/XI0/XI0_33/d_4_ DECAP_INV_G11
XG1282 XI11_7/XI0/XI0_33/d__3_ XI11_7/XI0/XI0_33/d_3_ DECAP_INV_G11
XG1283 XI11_7/XI0/XI0_33/d__2_ XI11_7/XI0/XI0_33/d_2_ DECAP_INV_G11
XG1284 XI11_7/XI0/XI0_33/d__1_ XI11_7/XI0/XI0_33/d_1_ DECAP_INV_G11
XG1285 XI11_7/XI0/XI0_33/d__0_ XI11_7/XI0/XI0_33/d_0_ DECAP_INV_G11
XG1286 XI11_7/XI0/XI0_33/d_15_ XI11_7/XI0/XI0_33/d__15_ DECAP_INV_G11
XG1287 XI11_7/XI0/XI0_33/d_14_ XI11_7/XI0/XI0_33/d__14_ DECAP_INV_G11
XG1288 XI11_7/XI0/XI0_33/d_13_ XI11_7/XI0/XI0_33/d__13_ DECAP_INV_G11
XG1289 XI11_7/XI0/XI0_33/d_12_ XI11_7/XI0/XI0_33/d__12_ DECAP_INV_G11
XG1290 XI11_7/XI0/XI0_33/d_11_ XI11_7/XI0/XI0_33/d__11_ DECAP_INV_G11
XG1291 XI11_7/XI0/XI0_33/d_10_ XI11_7/XI0/XI0_33/d__10_ DECAP_INV_G11
XG1292 XI11_7/XI0/XI0_33/d_9_ XI11_7/XI0/XI0_33/d__9_ DECAP_INV_G11
XG1293 XI11_7/XI0/XI0_33/d_8_ XI11_7/XI0/XI0_33/d__8_ DECAP_INV_G11
XG1294 XI11_7/XI0/XI0_33/d_7_ XI11_7/XI0/XI0_33/d__7_ DECAP_INV_G11
XG1295 XI11_7/XI0/XI0_33/d_6_ XI11_7/XI0/XI0_33/d__6_ DECAP_INV_G11
XG1296 XI11_7/XI0/XI0_33/d_5_ XI11_7/XI0/XI0_33/d__5_ DECAP_INV_G11
XG1297 XI11_7/XI0/XI0_33/d_4_ XI11_7/XI0/XI0_33/d__4_ DECAP_INV_G11
XG1298 XI11_7/XI0/XI0_33/d_3_ XI11_7/XI0/XI0_33/d__3_ DECAP_INV_G11
XG1299 XI11_7/XI0/XI0_33/d_2_ XI11_7/XI0/XI0_33/d__2_ DECAP_INV_G11
XG1300 XI11_7/XI0/XI0_33/d_1_ XI11_7/XI0/XI0_33/d__1_ DECAP_INV_G11
XG1301 XI11_7/XI0/XI0_33/d_0_ XI11_7/XI0/XI0_33/d__0_ DECAP_INV_G11
XG1302 XI11_7/XI0/XI0_32/d__15_ XI11_7/XI0/XI0_32/d_15_ DECAP_INV_G11
XG1303 XI11_7/XI0/XI0_32/d__14_ XI11_7/XI0/XI0_32/d_14_ DECAP_INV_G11
XG1304 XI11_7/XI0/XI0_32/d__13_ XI11_7/XI0/XI0_32/d_13_ DECAP_INV_G11
XG1305 XI11_7/XI0/XI0_32/d__12_ XI11_7/XI0/XI0_32/d_12_ DECAP_INV_G11
XG1306 XI11_7/XI0/XI0_32/d__11_ XI11_7/XI0/XI0_32/d_11_ DECAP_INV_G11
XG1307 XI11_7/XI0/XI0_32/d__10_ XI11_7/XI0/XI0_32/d_10_ DECAP_INV_G11
XG1308 XI11_7/XI0/XI0_32/d__9_ XI11_7/XI0/XI0_32/d_9_ DECAP_INV_G11
XG1309 XI11_7/XI0/XI0_32/d__8_ XI11_7/XI0/XI0_32/d_8_ DECAP_INV_G11
XG1310 XI11_7/XI0/XI0_32/d__7_ XI11_7/XI0/XI0_32/d_7_ DECAP_INV_G11
XG1311 XI11_7/XI0/XI0_32/d__6_ XI11_7/XI0/XI0_32/d_6_ DECAP_INV_G11
XG1312 XI11_7/XI0/XI0_32/d__5_ XI11_7/XI0/XI0_32/d_5_ DECAP_INV_G11
XG1313 XI11_7/XI0/XI0_32/d__4_ XI11_7/XI0/XI0_32/d_4_ DECAP_INV_G11
XG1314 XI11_7/XI0/XI0_32/d__3_ XI11_7/XI0/XI0_32/d_3_ DECAP_INV_G11
XG1315 XI11_7/XI0/XI0_32/d__2_ XI11_7/XI0/XI0_32/d_2_ DECAP_INV_G11
XG1316 XI11_7/XI0/XI0_32/d__1_ XI11_7/XI0/XI0_32/d_1_ DECAP_INV_G11
XG1317 XI11_7/XI0/XI0_32/d__0_ XI11_7/XI0/XI0_32/d_0_ DECAP_INV_G11
XG1318 XI11_7/XI0/XI0_32/d_15_ XI11_7/XI0/XI0_32/d__15_ DECAP_INV_G11
XG1319 XI11_7/XI0/XI0_32/d_14_ XI11_7/XI0/XI0_32/d__14_ DECAP_INV_G11
XG1320 XI11_7/XI0/XI0_32/d_13_ XI11_7/XI0/XI0_32/d__13_ DECAP_INV_G11
XG1321 XI11_7/XI0/XI0_32/d_12_ XI11_7/XI0/XI0_32/d__12_ DECAP_INV_G11
XG1322 XI11_7/XI0/XI0_32/d_11_ XI11_7/XI0/XI0_32/d__11_ DECAP_INV_G11
XG1323 XI11_7/XI0/XI0_32/d_10_ XI11_7/XI0/XI0_32/d__10_ DECAP_INV_G11
XG1324 XI11_7/XI0/XI0_32/d_9_ XI11_7/XI0/XI0_32/d__9_ DECAP_INV_G11
XG1325 XI11_7/XI0/XI0_32/d_8_ XI11_7/XI0/XI0_32/d__8_ DECAP_INV_G11
XG1326 XI11_7/XI0/XI0_32/d_7_ XI11_7/XI0/XI0_32/d__7_ DECAP_INV_G11
XG1327 XI11_7/XI0/XI0_32/d_6_ XI11_7/XI0/XI0_32/d__6_ DECAP_INV_G11
XG1328 XI11_7/XI0/XI0_32/d_5_ XI11_7/XI0/XI0_32/d__5_ DECAP_INV_G11
XG1329 XI11_7/XI0/XI0_32/d_4_ XI11_7/XI0/XI0_32/d__4_ DECAP_INV_G11
XG1330 XI11_7/XI0/XI0_32/d_3_ XI11_7/XI0/XI0_32/d__3_ DECAP_INV_G11
XG1331 XI11_7/XI0/XI0_32/d_2_ XI11_7/XI0/XI0_32/d__2_ DECAP_INV_G11
XG1332 XI11_7/XI0/XI0_32/d_1_ XI11_7/XI0/XI0_32/d__1_ DECAP_INV_G11
XG1333 XI11_7/XI0/XI0_32/d_0_ XI11_7/XI0/XI0_32/d__0_ DECAP_INV_G11
XG1334 XI11_7/XI0/XI0_31/d__15_ XI11_7/XI0/XI0_31/d_15_ DECAP_INV_G11
XG1335 XI11_7/XI0/XI0_31/d__14_ XI11_7/XI0/XI0_31/d_14_ DECAP_INV_G11
XG1336 XI11_7/XI0/XI0_31/d__13_ XI11_7/XI0/XI0_31/d_13_ DECAP_INV_G11
XG1337 XI11_7/XI0/XI0_31/d__12_ XI11_7/XI0/XI0_31/d_12_ DECAP_INV_G11
XG1338 XI11_7/XI0/XI0_31/d__11_ XI11_7/XI0/XI0_31/d_11_ DECAP_INV_G11
XG1339 XI11_7/XI0/XI0_31/d__10_ XI11_7/XI0/XI0_31/d_10_ DECAP_INV_G11
XG1340 XI11_7/XI0/XI0_31/d__9_ XI11_7/XI0/XI0_31/d_9_ DECAP_INV_G11
XG1341 XI11_7/XI0/XI0_31/d__8_ XI11_7/XI0/XI0_31/d_8_ DECAP_INV_G11
XG1342 XI11_7/XI0/XI0_31/d__7_ XI11_7/XI0/XI0_31/d_7_ DECAP_INV_G11
XG1343 XI11_7/XI0/XI0_31/d__6_ XI11_7/XI0/XI0_31/d_6_ DECAP_INV_G11
XG1344 XI11_7/XI0/XI0_31/d__5_ XI11_7/XI0/XI0_31/d_5_ DECAP_INV_G11
XG1345 XI11_7/XI0/XI0_31/d__4_ XI11_7/XI0/XI0_31/d_4_ DECAP_INV_G11
XG1346 XI11_7/XI0/XI0_31/d__3_ XI11_7/XI0/XI0_31/d_3_ DECAP_INV_G11
XG1347 XI11_7/XI0/XI0_31/d__2_ XI11_7/XI0/XI0_31/d_2_ DECAP_INV_G11
XG1348 XI11_7/XI0/XI0_31/d__1_ XI11_7/XI0/XI0_31/d_1_ DECAP_INV_G11
XG1349 XI11_7/XI0/XI0_31/d__0_ XI11_7/XI0/XI0_31/d_0_ DECAP_INV_G11
XG1350 XI11_7/XI0/XI0_31/d_15_ XI11_7/XI0/XI0_31/d__15_ DECAP_INV_G11
XG1351 XI11_7/XI0/XI0_31/d_14_ XI11_7/XI0/XI0_31/d__14_ DECAP_INV_G11
XG1352 XI11_7/XI0/XI0_31/d_13_ XI11_7/XI0/XI0_31/d__13_ DECAP_INV_G11
XG1353 XI11_7/XI0/XI0_31/d_12_ XI11_7/XI0/XI0_31/d__12_ DECAP_INV_G11
XG1354 XI11_7/XI0/XI0_31/d_11_ XI11_7/XI0/XI0_31/d__11_ DECAP_INV_G11
XG1355 XI11_7/XI0/XI0_31/d_10_ XI11_7/XI0/XI0_31/d__10_ DECAP_INV_G11
XG1356 XI11_7/XI0/XI0_31/d_9_ XI11_7/XI0/XI0_31/d__9_ DECAP_INV_G11
XG1357 XI11_7/XI0/XI0_31/d_8_ XI11_7/XI0/XI0_31/d__8_ DECAP_INV_G11
XG1358 XI11_7/XI0/XI0_31/d_7_ XI11_7/XI0/XI0_31/d__7_ DECAP_INV_G11
XG1359 XI11_7/XI0/XI0_31/d_6_ XI11_7/XI0/XI0_31/d__6_ DECAP_INV_G11
XG1360 XI11_7/XI0/XI0_31/d_5_ XI11_7/XI0/XI0_31/d__5_ DECAP_INV_G11
XG1361 XI11_7/XI0/XI0_31/d_4_ XI11_7/XI0/XI0_31/d__4_ DECAP_INV_G11
XG1362 XI11_7/XI0/XI0_31/d_3_ XI11_7/XI0/XI0_31/d__3_ DECAP_INV_G11
XG1363 XI11_7/XI0/XI0_31/d_2_ XI11_7/XI0/XI0_31/d__2_ DECAP_INV_G11
XG1364 XI11_7/XI0/XI0_31/d_1_ XI11_7/XI0/XI0_31/d__1_ DECAP_INV_G11
XG1365 XI11_7/XI0/XI0_31/d_0_ XI11_7/XI0/XI0_31/d__0_ DECAP_INV_G11
XG1366 XI11_7/XI0/XI0_30/d__15_ XI11_7/XI0/XI0_30/d_15_ DECAP_INV_G11
XG1367 XI11_7/XI0/XI0_30/d__14_ XI11_7/XI0/XI0_30/d_14_ DECAP_INV_G11
XG1368 XI11_7/XI0/XI0_30/d__13_ XI11_7/XI0/XI0_30/d_13_ DECAP_INV_G11
XG1369 XI11_7/XI0/XI0_30/d__12_ XI11_7/XI0/XI0_30/d_12_ DECAP_INV_G11
XG1370 XI11_7/XI0/XI0_30/d__11_ XI11_7/XI0/XI0_30/d_11_ DECAP_INV_G11
XG1371 XI11_7/XI0/XI0_30/d__10_ XI11_7/XI0/XI0_30/d_10_ DECAP_INV_G11
XG1372 XI11_7/XI0/XI0_30/d__9_ XI11_7/XI0/XI0_30/d_9_ DECAP_INV_G11
XG1373 XI11_7/XI0/XI0_30/d__8_ XI11_7/XI0/XI0_30/d_8_ DECAP_INV_G11
XG1374 XI11_7/XI0/XI0_30/d__7_ XI11_7/XI0/XI0_30/d_7_ DECAP_INV_G11
XG1375 XI11_7/XI0/XI0_30/d__6_ XI11_7/XI0/XI0_30/d_6_ DECAP_INV_G11
XG1376 XI11_7/XI0/XI0_30/d__5_ XI11_7/XI0/XI0_30/d_5_ DECAP_INV_G11
XG1377 XI11_7/XI0/XI0_30/d__4_ XI11_7/XI0/XI0_30/d_4_ DECAP_INV_G11
XG1378 XI11_7/XI0/XI0_30/d__3_ XI11_7/XI0/XI0_30/d_3_ DECAP_INV_G11
XG1379 XI11_7/XI0/XI0_30/d__2_ XI11_7/XI0/XI0_30/d_2_ DECAP_INV_G11
XG1380 XI11_7/XI0/XI0_30/d__1_ XI11_7/XI0/XI0_30/d_1_ DECAP_INV_G11
XG1381 XI11_7/XI0/XI0_30/d__0_ XI11_7/XI0/XI0_30/d_0_ DECAP_INV_G11
XG1382 XI11_7/XI0/XI0_30/d_15_ XI11_7/XI0/XI0_30/d__15_ DECAP_INV_G11
XG1383 XI11_7/XI0/XI0_30/d_14_ XI11_7/XI0/XI0_30/d__14_ DECAP_INV_G11
XG1384 XI11_7/XI0/XI0_30/d_13_ XI11_7/XI0/XI0_30/d__13_ DECAP_INV_G11
XG1385 XI11_7/XI0/XI0_30/d_12_ XI11_7/XI0/XI0_30/d__12_ DECAP_INV_G11
XG1386 XI11_7/XI0/XI0_30/d_11_ XI11_7/XI0/XI0_30/d__11_ DECAP_INV_G11
XG1387 XI11_7/XI0/XI0_30/d_10_ XI11_7/XI0/XI0_30/d__10_ DECAP_INV_G11
XG1388 XI11_7/XI0/XI0_30/d_9_ XI11_7/XI0/XI0_30/d__9_ DECAP_INV_G11
XG1389 XI11_7/XI0/XI0_30/d_8_ XI11_7/XI0/XI0_30/d__8_ DECAP_INV_G11
XG1390 XI11_7/XI0/XI0_30/d_7_ XI11_7/XI0/XI0_30/d__7_ DECAP_INV_G11
XG1391 XI11_7/XI0/XI0_30/d_6_ XI11_7/XI0/XI0_30/d__6_ DECAP_INV_G11
XG1392 XI11_7/XI0/XI0_30/d_5_ XI11_7/XI0/XI0_30/d__5_ DECAP_INV_G11
XG1393 XI11_7/XI0/XI0_30/d_4_ XI11_7/XI0/XI0_30/d__4_ DECAP_INV_G11
XG1394 XI11_7/XI0/XI0_30/d_3_ XI11_7/XI0/XI0_30/d__3_ DECAP_INV_G11
XG1395 XI11_7/XI0/XI0_30/d_2_ XI11_7/XI0/XI0_30/d__2_ DECAP_INV_G11
XG1396 XI11_7/XI0/XI0_30/d_1_ XI11_7/XI0/XI0_30/d__1_ DECAP_INV_G11
XG1397 XI11_7/XI0/XI0_30/d_0_ XI11_7/XI0/XI0_30/d__0_ DECAP_INV_G11
XG1398 XI11_7/XI0/XI0_29/d__15_ XI11_7/XI0/XI0_29/d_15_ DECAP_INV_G11
XG1399 XI11_7/XI0/XI0_29/d__14_ XI11_7/XI0/XI0_29/d_14_ DECAP_INV_G11
XG1400 XI11_7/XI0/XI0_29/d__13_ XI11_7/XI0/XI0_29/d_13_ DECAP_INV_G11
XG1401 XI11_7/XI0/XI0_29/d__12_ XI11_7/XI0/XI0_29/d_12_ DECAP_INV_G11
XG1402 XI11_7/XI0/XI0_29/d__11_ XI11_7/XI0/XI0_29/d_11_ DECAP_INV_G11
XG1403 XI11_7/XI0/XI0_29/d__10_ XI11_7/XI0/XI0_29/d_10_ DECAP_INV_G11
XG1404 XI11_7/XI0/XI0_29/d__9_ XI11_7/XI0/XI0_29/d_9_ DECAP_INV_G11
XG1405 XI11_7/XI0/XI0_29/d__8_ XI11_7/XI0/XI0_29/d_8_ DECAP_INV_G11
XG1406 XI11_7/XI0/XI0_29/d__7_ XI11_7/XI0/XI0_29/d_7_ DECAP_INV_G11
XG1407 XI11_7/XI0/XI0_29/d__6_ XI11_7/XI0/XI0_29/d_6_ DECAP_INV_G11
XG1408 XI11_7/XI0/XI0_29/d__5_ XI11_7/XI0/XI0_29/d_5_ DECAP_INV_G11
XG1409 XI11_7/XI0/XI0_29/d__4_ XI11_7/XI0/XI0_29/d_4_ DECAP_INV_G11
XG1410 XI11_7/XI0/XI0_29/d__3_ XI11_7/XI0/XI0_29/d_3_ DECAP_INV_G11
XG1411 XI11_7/XI0/XI0_29/d__2_ XI11_7/XI0/XI0_29/d_2_ DECAP_INV_G11
XG1412 XI11_7/XI0/XI0_29/d__1_ XI11_7/XI0/XI0_29/d_1_ DECAP_INV_G11
XG1413 XI11_7/XI0/XI0_29/d__0_ XI11_7/XI0/XI0_29/d_0_ DECAP_INV_G11
XG1414 XI11_7/XI0/XI0_29/d_15_ XI11_7/XI0/XI0_29/d__15_ DECAP_INV_G11
XG1415 XI11_7/XI0/XI0_29/d_14_ XI11_7/XI0/XI0_29/d__14_ DECAP_INV_G11
XG1416 XI11_7/XI0/XI0_29/d_13_ XI11_7/XI0/XI0_29/d__13_ DECAP_INV_G11
XG1417 XI11_7/XI0/XI0_29/d_12_ XI11_7/XI0/XI0_29/d__12_ DECAP_INV_G11
XG1418 XI11_7/XI0/XI0_29/d_11_ XI11_7/XI0/XI0_29/d__11_ DECAP_INV_G11
XG1419 XI11_7/XI0/XI0_29/d_10_ XI11_7/XI0/XI0_29/d__10_ DECAP_INV_G11
XG1420 XI11_7/XI0/XI0_29/d_9_ XI11_7/XI0/XI0_29/d__9_ DECAP_INV_G11
XG1421 XI11_7/XI0/XI0_29/d_8_ XI11_7/XI0/XI0_29/d__8_ DECAP_INV_G11
XG1422 XI11_7/XI0/XI0_29/d_7_ XI11_7/XI0/XI0_29/d__7_ DECAP_INV_G11
XG1423 XI11_7/XI0/XI0_29/d_6_ XI11_7/XI0/XI0_29/d__6_ DECAP_INV_G11
XG1424 XI11_7/XI0/XI0_29/d_5_ XI11_7/XI0/XI0_29/d__5_ DECAP_INV_G11
XG1425 XI11_7/XI0/XI0_29/d_4_ XI11_7/XI0/XI0_29/d__4_ DECAP_INV_G11
XG1426 XI11_7/XI0/XI0_29/d_3_ XI11_7/XI0/XI0_29/d__3_ DECAP_INV_G11
XG1427 XI11_7/XI0/XI0_29/d_2_ XI11_7/XI0/XI0_29/d__2_ DECAP_INV_G11
XG1428 XI11_7/XI0/XI0_29/d_1_ XI11_7/XI0/XI0_29/d__1_ DECAP_INV_G11
XG1429 XI11_7/XI0/XI0_29/d_0_ XI11_7/XI0/XI0_29/d__0_ DECAP_INV_G11
XG1430 XI11_7/XI0/XI0_28/d__15_ XI11_7/XI0/XI0_28/d_15_ DECAP_INV_G11
XG1431 XI11_7/XI0/XI0_28/d__14_ XI11_7/XI0/XI0_28/d_14_ DECAP_INV_G11
XG1432 XI11_7/XI0/XI0_28/d__13_ XI11_7/XI0/XI0_28/d_13_ DECAP_INV_G11
XG1433 XI11_7/XI0/XI0_28/d__12_ XI11_7/XI0/XI0_28/d_12_ DECAP_INV_G11
XG1434 XI11_7/XI0/XI0_28/d__11_ XI11_7/XI0/XI0_28/d_11_ DECAP_INV_G11
XG1435 XI11_7/XI0/XI0_28/d__10_ XI11_7/XI0/XI0_28/d_10_ DECAP_INV_G11
XG1436 XI11_7/XI0/XI0_28/d__9_ XI11_7/XI0/XI0_28/d_9_ DECAP_INV_G11
XG1437 XI11_7/XI0/XI0_28/d__8_ XI11_7/XI0/XI0_28/d_8_ DECAP_INV_G11
XG1438 XI11_7/XI0/XI0_28/d__7_ XI11_7/XI0/XI0_28/d_7_ DECAP_INV_G11
XG1439 XI11_7/XI0/XI0_28/d__6_ XI11_7/XI0/XI0_28/d_6_ DECAP_INV_G11
XG1440 XI11_7/XI0/XI0_28/d__5_ XI11_7/XI0/XI0_28/d_5_ DECAP_INV_G11
XG1441 XI11_7/XI0/XI0_28/d__4_ XI11_7/XI0/XI0_28/d_4_ DECAP_INV_G11
XG1442 XI11_7/XI0/XI0_28/d__3_ XI11_7/XI0/XI0_28/d_3_ DECAP_INV_G11
XG1443 XI11_7/XI0/XI0_28/d__2_ XI11_7/XI0/XI0_28/d_2_ DECAP_INV_G11
XG1444 XI11_7/XI0/XI0_28/d__1_ XI11_7/XI0/XI0_28/d_1_ DECAP_INV_G11
XG1445 XI11_7/XI0/XI0_28/d__0_ XI11_7/XI0/XI0_28/d_0_ DECAP_INV_G11
XG1446 XI11_7/XI0/XI0_28/d_15_ XI11_7/XI0/XI0_28/d__15_ DECAP_INV_G11
XG1447 XI11_7/XI0/XI0_28/d_14_ XI11_7/XI0/XI0_28/d__14_ DECAP_INV_G11
XG1448 XI11_7/XI0/XI0_28/d_13_ XI11_7/XI0/XI0_28/d__13_ DECAP_INV_G11
XG1449 XI11_7/XI0/XI0_28/d_12_ XI11_7/XI0/XI0_28/d__12_ DECAP_INV_G11
XG1450 XI11_7/XI0/XI0_28/d_11_ XI11_7/XI0/XI0_28/d__11_ DECAP_INV_G11
XG1451 XI11_7/XI0/XI0_28/d_10_ XI11_7/XI0/XI0_28/d__10_ DECAP_INV_G11
XG1452 XI11_7/XI0/XI0_28/d_9_ XI11_7/XI0/XI0_28/d__9_ DECAP_INV_G11
XG1453 XI11_7/XI0/XI0_28/d_8_ XI11_7/XI0/XI0_28/d__8_ DECAP_INV_G11
XG1454 XI11_7/XI0/XI0_28/d_7_ XI11_7/XI0/XI0_28/d__7_ DECAP_INV_G11
XG1455 XI11_7/XI0/XI0_28/d_6_ XI11_7/XI0/XI0_28/d__6_ DECAP_INV_G11
XG1456 XI11_7/XI0/XI0_28/d_5_ XI11_7/XI0/XI0_28/d__5_ DECAP_INV_G11
XG1457 XI11_7/XI0/XI0_28/d_4_ XI11_7/XI0/XI0_28/d__4_ DECAP_INV_G11
XG1458 XI11_7/XI0/XI0_28/d_3_ XI11_7/XI0/XI0_28/d__3_ DECAP_INV_G11
XG1459 XI11_7/XI0/XI0_28/d_2_ XI11_7/XI0/XI0_28/d__2_ DECAP_INV_G11
XG1460 XI11_7/XI0/XI0_28/d_1_ XI11_7/XI0/XI0_28/d__1_ DECAP_INV_G11
XG1461 XI11_7/XI0/XI0_28/d_0_ XI11_7/XI0/XI0_28/d__0_ DECAP_INV_G11
XG1462 XI11_7/XI0/XI0_27/d__15_ XI11_7/XI0/XI0_27/d_15_ DECAP_INV_G11
XG1463 XI11_7/XI0/XI0_27/d__14_ XI11_7/XI0/XI0_27/d_14_ DECAP_INV_G11
XG1464 XI11_7/XI0/XI0_27/d__13_ XI11_7/XI0/XI0_27/d_13_ DECAP_INV_G11
XG1465 XI11_7/XI0/XI0_27/d__12_ XI11_7/XI0/XI0_27/d_12_ DECAP_INV_G11
XG1466 XI11_7/XI0/XI0_27/d__11_ XI11_7/XI0/XI0_27/d_11_ DECAP_INV_G11
XG1467 XI11_7/XI0/XI0_27/d__10_ XI11_7/XI0/XI0_27/d_10_ DECAP_INV_G11
XG1468 XI11_7/XI0/XI0_27/d__9_ XI11_7/XI0/XI0_27/d_9_ DECAP_INV_G11
XG1469 XI11_7/XI0/XI0_27/d__8_ XI11_7/XI0/XI0_27/d_8_ DECAP_INV_G11
XG1470 XI11_7/XI0/XI0_27/d__7_ XI11_7/XI0/XI0_27/d_7_ DECAP_INV_G11
XG1471 XI11_7/XI0/XI0_27/d__6_ XI11_7/XI0/XI0_27/d_6_ DECAP_INV_G11
XG1472 XI11_7/XI0/XI0_27/d__5_ XI11_7/XI0/XI0_27/d_5_ DECAP_INV_G11
XG1473 XI11_7/XI0/XI0_27/d__4_ XI11_7/XI0/XI0_27/d_4_ DECAP_INV_G11
XG1474 XI11_7/XI0/XI0_27/d__3_ XI11_7/XI0/XI0_27/d_3_ DECAP_INV_G11
XG1475 XI11_7/XI0/XI0_27/d__2_ XI11_7/XI0/XI0_27/d_2_ DECAP_INV_G11
XG1476 XI11_7/XI0/XI0_27/d__1_ XI11_7/XI0/XI0_27/d_1_ DECAP_INV_G11
XG1477 XI11_7/XI0/XI0_27/d__0_ XI11_7/XI0/XI0_27/d_0_ DECAP_INV_G11
XG1478 XI11_7/XI0/XI0_27/d_15_ XI11_7/XI0/XI0_27/d__15_ DECAP_INV_G11
XG1479 XI11_7/XI0/XI0_27/d_14_ XI11_7/XI0/XI0_27/d__14_ DECAP_INV_G11
XG1480 XI11_7/XI0/XI0_27/d_13_ XI11_7/XI0/XI0_27/d__13_ DECAP_INV_G11
XG1481 XI11_7/XI0/XI0_27/d_12_ XI11_7/XI0/XI0_27/d__12_ DECAP_INV_G11
XG1482 XI11_7/XI0/XI0_27/d_11_ XI11_7/XI0/XI0_27/d__11_ DECAP_INV_G11
XG1483 XI11_7/XI0/XI0_27/d_10_ XI11_7/XI0/XI0_27/d__10_ DECAP_INV_G11
XG1484 XI11_7/XI0/XI0_27/d_9_ XI11_7/XI0/XI0_27/d__9_ DECAP_INV_G11
XG1485 XI11_7/XI0/XI0_27/d_8_ XI11_7/XI0/XI0_27/d__8_ DECAP_INV_G11
XG1486 XI11_7/XI0/XI0_27/d_7_ XI11_7/XI0/XI0_27/d__7_ DECAP_INV_G11
XG1487 XI11_7/XI0/XI0_27/d_6_ XI11_7/XI0/XI0_27/d__6_ DECAP_INV_G11
XG1488 XI11_7/XI0/XI0_27/d_5_ XI11_7/XI0/XI0_27/d__5_ DECAP_INV_G11
XG1489 XI11_7/XI0/XI0_27/d_4_ XI11_7/XI0/XI0_27/d__4_ DECAP_INV_G11
XG1490 XI11_7/XI0/XI0_27/d_3_ XI11_7/XI0/XI0_27/d__3_ DECAP_INV_G11
XG1491 XI11_7/XI0/XI0_27/d_2_ XI11_7/XI0/XI0_27/d__2_ DECAP_INV_G11
XG1492 XI11_7/XI0/XI0_27/d_1_ XI11_7/XI0/XI0_27/d__1_ DECAP_INV_G11
XG1493 XI11_7/XI0/XI0_27/d_0_ XI11_7/XI0/XI0_27/d__0_ DECAP_INV_G11
XG1494 XI11_7/XI0/XI0_26/d__15_ XI11_7/XI0/XI0_26/d_15_ DECAP_INV_G11
XG1495 XI11_7/XI0/XI0_26/d__14_ XI11_7/XI0/XI0_26/d_14_ DECAP_INV_G11
XG1496 XI11_7/XI0/XI0_26/d__13_ XI11_7/XI0/XI0_26/d_13_ DECAP_INV_G11
XG1497 XI11_7/XI0/XI0_26/d__12_ XI11_7/XI0/XI0_26/d_12_ DECAP_INV_G11
XG1498 XI11_7/XI0/XI0_26/d__11_ XI11_7/XI0/XI0_26/d_11_ DECAP_INV_G11
XG1499 XI11_7/XI0/XI0_26/d__10_ XI11_7/XI0/XI0_26/d_10_ DECAP_INV_G11
XG1500 XI11_7/XI0/XI0_26/d__9_ XI11_7/XI0/XI0_26/d_9_ DECAP_INV_G11
XG1501 XI11_7/XI0/XI0_26/d__8_ XI11_7/XI0/XI0_26/d_8_ DECAP_INV_G11
XG1502 XI11_7/XI0/XI0_26/d__7_ XI11_7/XI0/XI0_26/d_7_ DECAP_INV_G11
XG1503 XI11_7/XI0/XI0_26/d__6_ XI11_7/XI0/XI0_26/d_6_ DECAP_INV_G11
XG1504 XI11_7/XI0/XI0_26/d__5_ XI11_7/XI0/XI0_26/d_5_ DECAP_INV_G11
XG1505 XI11_7/XI0/XI0_26/d__4_ XI11_7/XI0/XI0_26/d_4_ DECAP_INV_G11
XG1506 XI11_7/XI0/XI0_26/d__3_ XI11_7/XI0/XI0_26/d_3_ DECAP_INV_G11
XG1507 XI11_7/XI0/XI0_26/d__2_ XI11_7/XI0/XI0_26/d_2_ DECAP_INV_G11
XG1508 XI11_7/XI0/XI0_26/d__1_ XI11_7/XI0/XI0_26/d_1_ DECAP_INV_G11
XG1509 XI11_7/XI0/XI0_26/d__0_ XI11_7/XI0/XI0_26/d_0_ DECAP_INV_G11
XG1510 XI11_7/XI0/XI0_26/d_15_ XI11_7/XI0/XI0_26/d__15_ DECAP_INV_G11
XG1511 XI11_7/XI0/XI0_26/d_14_ XI11_7/XI0/XI0_26/d__14_ DECAP_INV_G11
XG1512 XI11_7/XI0/XI0_26/d_13_ XI11_7/XI0/XI0_26/d__13_ DECAP_INV_G11
XG1513 XI11_7/XI0/XI0_26/d_12_ XI11_7/XI0/XI0_26/d__12_ DECAP_INV_G11
XG1514 XI11_7/XI0/XI0_26/d_11_ XI11_7/XI0/XI0_26/d__11_ DECAP_INV_G11
XG1515 XI11_7/XI0/XI0_26/d_10_ XI11_7/XI0/XI0_26/d__10_ DECAP_INV_G11
XG1516 XI11_7/XI0/XI0_26/d_9_ XI11_7/XI0/XI0_26/d__9_ DECAP_INV_G11
XG1517 XI11_7/XI0/XI0_26/d_8_ XI11_7/XI0/XI0_26/d__8_ DECAP_INV_G11
XG1518 XI11_7/XI0/XI0_26/d_7_ XI11_7/XI0/XI0_26/d__7_ DECAP_INV_G11
XG1519 XI11_7/XI0/XI0_26/d_6_ XI11_7/XI0/XI0_26/d__6_ DECAP_INV_G11
XG1520 XI11_7/XI0/XI0_26/d_5_ XI11_7/XI0/XI0_26/d__5_ DECAP_INV_G11
XG1521 XI11_7/XI0/XI0_26/d_4_ XI11_7/XI0/XI0_26/d__4_ DECAP_INV_G11
XG1522 XI11_7/XI0/XI0_26/d_3_ XI11_7/XI0/XI0_26/d__3_ DECAP_INV_G11
XG1523 XI11_7/XI0/XI0_26/d_2_ XI11_7/XI0/XI0_26/d__2_ DECAP_INV_G11
XG1524 XI11_7/XI0/XI0_26/d_1_ XI11_7/XI0/XI0_26/d__1_ DECAP_INV_G11
XG1525 XI11_7/XI0/XI0_26/d_0_ XI11_7/XI0/XI0_26/d__0_ DECAP_INV_G11
XG1526 XI11_7/XI0/XI0_25/d__15_ XI11_7/XI0/XI0_25/d_15_ DECAP_INV_G11
XG1527 XI11_7/XI0/XI0_25/d__14_ XI11_7/XI0/XI0_25/d_14_ DECAP_INV_G11
XG1528 XI11_7/XI0/XI0_25/d__13_ XI11_7/XI0/XI0_25/d_13_ DECAP_INV_G11
XG1529 XI11_7/XI0/XI0_25/d__12_ XI11_7/XI0/XI0_25/d_12_ DECAP_INV_G11
XG1530 XI11_7/XI0/XI0_25/d__11_ XI11_7/XI0/XI0_25/d_11_ DECAP_INV_G11
XG1531 XI11_7/XI0/XI0_25/d__10_ XI11_7/XI0/XI0_25/d_10_ DECAP_INV_G11
XG1532 XI11_7/XI0/XI0_25/d__9_ XI11_7/XI0/XI0_25/d_9_ DECAP_INV_G11
XG1533 XI11_7/XI0/XI0_25/d__8_ XI11_7/XI0/XI0_25/d_8_ DECAP_INV_G11
XG1534 XI11_7/XI0/XI0_25/d__7_ XI11_7/XI0/XI0_25/d_7_ DECAP_INV_G11
XG1535 XI11_7/XI0/XI0_25/d__6_ XI11_7/XI0/XI0_25/d_6_ DECAP_INV_G11
XG1536 XI11_7/XI0/XI0_25/d__5_ XI11_7/XI0/XI0_25/d_5_ DECAP_INV_G11
XG1537 XI11_7/XI0/XI0_25/d__4_ XI11_7/XI0/XI0_25/d_4_ DECAP_INV_G11
XG1538 XI11_7/XI0/XI0_25/d__3_ XI11_7/XI0/XI0_25/d_3_ DECAP_INV_G11
XG1539 XI11_7/XI0/XI0_25/d__2_ XI11_7/XI0/XI0_25/d_2_ DECAP_INV_G11
XG1540 XI11_7/XI0/XI0_25/d__1_ XI11_7/XI0/XI0_25/d_1_ DECAP_INV_G11
XG1541 XI11_7/XI0/XI0_25/d__0_ XI11_7/XI0/XI0_25/d_0_ DECAP_INV_G11
XG1542 XI11_7/XI0/XI0_25/d_15_ XI11_7/XI0/XI0_25/d__15_ DECAP_INV_G11
XG1543 XI11_7/XI0/XI0_25/d_14_ XI11_7/XI0/XI0_25/d__14_ DECAP_INV_G11
XG1544 XI11_7/XI0/XI0_25/d_13_ XI11_7/XI0/XI0_25/d__13_ DECAP_INV_G11
XG1545 XI11_7/XI0/XI0_25/d_12_ XI11_7/XI0/XI0_25/d__12_ DECAP_INV_G11
XG1546 XI11_7/XI0/XI0_25/d_11_ XI11_7/XI0/XI0_25/d__11_ DECAP_INV_G11
XG1547 XI11_7/XI0/XI0_25/d_10_ XI11_7/XI0/XI0_25/d__10_ DECAP_INV_G11
XG1548 XI11_7/XI0/XI0_25/d_9_ XI11_7/XI0/XI0_25/d__9_ DECAP_INV_G11
XG1549 XI11_7/XI0/XI0_25/d_8_ XI11_7/XI0/XI0_25/d__8_ DECAP_INV_G11
XG1550 XI11_7/XI0/XI0_25/d_7_ XI11_7/XI0/XI0_25/d__7_ DECAP_INV_G11
XG1551 XI11_7/XI0/XI0_25/d_6_ XI11_7/XI0/XI0_25/d__6_ DECAP_INV_G11
XG1552 XI11_7/XI0/XI0_25/d_5_ XI11_7/XI0/XI0_25/d__5_ DECAP_INV_G11
XG1553 XI11_7/XI0/XI0_25/d_4_ XI11_7/XI0/XI0_25/d__4_ DECAP_INV_G11
XG1554 XI11_7/XI0/XI0_25/d_3_ XI11_7/XI0/XI0_25/d__3_ DECAP_INV_G11
XG1555 XI11_7/XI0/XI0_25/d_2_ XI11_7/XI0/XI0_25/d__2_ DECAP_INV_G11
XG1556 XI11_7/XI0/XI0_25/d_1_ XI11_7/XI0/XI0_25/d__1_ DECAP_INV_G11
XG1557 XI11_7/XI0/XI0_25/d_0_ XI11_7/XI0/XI0_25/d__0_ DECAP_INV_G11
XG1558 XI11_7/XI0/XI0_24/d__15_ XI11_7/XI0/XI0_24/d_15_ DECAP_INV_G11
XG1559 XI11_7/XI0/XI0_24/d__14_ XI11_7/XI0/XI0_24/d_14_ DECAP_INV_G11
XG1560 XI11_7/XI0/XI0_24/d__13_ XI11_7/XI0/XI0_24/d_13_ DECAP_INV_G11
XG1561 XI11_7/XI0/XI0_24/d__12_ XI11_7/XI0/XI0_24/d_12_ DECAP_INV_G11
XG1562 XI11_7/XI0/XI0_24/d__11_ XI11_7/XI0/XI0_24/d_11_ DECAP_INV_G11
XG1563 XI11_7/XI0/XI0_24/d__10_ XI11_7/XI0/XI0_24/d_10_ DECAP_INV_G11
XG1564 XI11_7/XI0/XI0_24/d__9_ XI11_7/XI0/XI0_24/d_9_ DECAP_INV_G11
XG1565 XI11_7/XI0/XI0_24/d__8_ XI11_7/XI0/XI0_24/d_8_ DECAP_INV_G11
XG1566 XI11_7/XI0/XI0_24/d__7_ XI11_7/XI0/XI0_24/d_7_ DECAP_INV_G11
XG1567 XI11_7/XI0/XI0_24/d__6_ XI11_7/XI0/XI0_24/d_6_ DECAP_INV_G11
XG1568 XI11_7/XI0/XI0_24/d__5_ XI11_7/XI0/XI0_24/d_5_ DECAP_INV_G11
XG1569 XI11_7/XI0/XI0_24/d__4_ XI11_7/XI0/XI0_24/d_4_ DECAP_INV_G11
XG1570 XI11_7/XI0/XI0_24/d__3_ XI11_7/XI0/XI0_24/d_3_ DECAP_INV_G11
XG1571 XI11_7/XI0/XI0_24/d__2_ XI11_7/XI0/XI0_24/d_2_ DECAP_INV_G11
XG1572 XI11_7/XI0/XI0_24/d__1_ XI11_7/XI0/XI0_24/d_1_ DECAP_INV_G11
XG1573 XI11_7/XI0/XI0_24/d__0_ XI11_7/XI0/XI0_24/d_0_ DECAP_INV_G11
XG1574 XI11_7/XI0/XI0_24/d_15_ XI11_7/XI0/XI0_24/d__15_ DECAP_INV_G11
XG1575 XI11_7/XI0/XI0_24/d_14_ XI11_7/XI0/XI0_24/d__14_ DECAP_INV_G11
XG1576 XI11_7/XI0/XI0_24/d_13_ XI11_7/XI0/XI0_24/d__13_ DECAP_INV_G11
XG1577 XI11_7/XI0/XI0_24/d_12_ XI11_7/XI0/XI0_24/d__12_ DECAP_INV_G11
XG1578 XI11_7/XI0/XI0_24/d_11_ XI11_7/XI0/XI0_24/d__11_ DECAP_INV_G11
XG1579 XI11_7/XI0/XI0_24/d_10_ XI11_7/XI0/XI0_24/d__10_ DECAP_INV_G11
XG1580 XI11_7/XI0/XI0_24/d_9_ XI11_7/XI0/XI0_24/d__9_ DECAP_INV_G11
XG1581 XI11_7/XI0/XI0_24/d_8_ XI11_7/XI0/XI0_24/d__8_ DECAP_INV_G11
XG1582 XI11_7/XI0/XI0_24/d_7_ XI11_7/XI0/XI0_24/d__7_ DECAP_INV_G11
XG1583 XI11_7/XI0/XI0_24/d_6_ XI11_7/XI0/XI0_24/d__6_ DECAP_INV_G11
XG1584 XI11_7/XI0/XI0_24/d_5_ XI11_7/XI0/XI0_24/d__5_ DECAP_INV_G11
XG1585 XI11_7/XI0/XI0_24/d_4_ XI11_7/XI0/XI0_24/d__4_ DECAP_INV_G11
XG1586 XI11_7/XI0/XI0_24/d_3_ XI11_7/XI0/XI0_24/d__3_ DECAP_INV_G11
XG1587 XI11_7/XI0/XI0_24/d_2_ XI11_7/XI0/XI0_24/d__2_ DECAP_INV_G11
XG1588 XI11_7/XI0/XI0_24/d_1_ XI11_7/XI0/XI0_24/d__1_ DECAP_INV_G11
XG1589 XI11_7/XI0/XI0_24/d_0_ XI11_7/XI0/XI0_24/d__0_ DECAP_INV_G11
XG1590 XI11_7/XI0/XI0_23/d__15_ XI11_7/XI0/XI0_23/d_15_ DECAP_INV_G11
XG1591 XI11_7/XI0/XI0_23/d__14_ XI11_7/XI0/XI0_23/d_14_ DECAP_INV_G11
XG1592 XI11_7/XI0/XI0_23/d__13_ XI11_7/XI0/XI0_23/d_13_ DECAP_INV_G11
XG1593 XI11_7/XI0/XI0_23/d__12_ XI11_7/XI0/XI0_23/d_12_ DECAP_INV_G11
XG1594 XI11_7/XI0/XI0_23/d__11_ XI11_7/XI0/XI0_23/d_11_ DECAP_INV_G11
XG1595 XI11_7/XI0/XI0_23/d__10_ XI11_7/XI0/XI0_23/d_10_ DECAP_INV_G11
XG1596 XI11_7/XI0/XI0_23/d__9_ XI11_7/XI0/XI0_23/d_9_ DECAP_INV_G11
XG1597 XI11_7/XI0/XI0_23/d__8_ XI11_7/XI0/XI0_23/d_8_ DECAP_INV_G11
XG1598 XI11_7/XI0/XI0_23/d__7_ XI11_7/XI0/XI0_23/d_7_ DECAP_INV_G11
XG1599 XI11_7/XI0/XI0_23/d__6_ XI11_7/XI0/XI0_23/d_6_ DECAP_INV_G11
XG1600 XI11_7/XI0/XI0_23/d__5_ XI11_7/XI0/XI0_23/d_5_ DECAP_INV_G11
XG1601 XI11_7/XI0/XI0_23/d__4_ XI11_7/XI0/XI0_23/d_4_ DECAP_INV_G11
XG1602 XI11_7/XI0/XI0_23/d__3_ XI11_7/XI0/XI0_23/d_3_ DECAP_INV_G11
XG1603 XI11_7/XI0/XI0_23/d__2_ XI11_7/XI0/XI0_23/d_2_ DECAP_INV_G11
XG1604 XI11_7/XI0/XI0_23/d__1_ XI11_7/XI0/XI0_23/d_1_ DECAP_INV_G11
XG1605 XI11_7/XI0/XI0_23/d__0_ XI11_7/XI0/XI0_23/d_0_ DECAP_INV_G11
XG1606 XI11_7/XI0/XI0_23/d_15_ XI11_7/XI0/XI0_23/d__15_ DECAP_INV_G11
XG1607 XI11_7/XI0/XI0_23/d_14_ XI11_7/XI0/XI0_23/d__14_ DECAP_INV_G11
XG1608 XI11_7/XI0/XI0_23/d_13_ XI11_7/XI0/XI0_23/d__13_ DECAP_INV_G11
XG1609 XI11_7/XI0/XI0_23/d_12_ XI11_7/XI0/XI0_23/d__12_ DECAP_INV_G11
XG1610 XI11_7/XI0/XI0_23/d_11_ XI11_7/XI0/XI0_23/d__11_ DECAP_INV_G11
XG1611 XI11_7/XI0/XI0_23/d_10_ XI11_7/XI0/XI0_23/d__10_ DECAP_INV_G11
XG1612 XI11_7/XI0/XI0_23/d_9_ XI11_7/XI0/XI0_23/d__9_ DECAP_INV_G11
XG1613 XI11_7/XI0/XI0_23/d_8_ XI11_7/XI0/XI0_23/d__8_ DECAP_INV_G11
XG1614 XI11_7/XI0/XI0_23/d_7_ XI11_7/XI0/XI0_23/d__7_ DECAP_INV_G11
XG1615 XI11_7/XI0/XI0_23/d_6_ XI11_7/XI0/XI0_23/d__6_ DECAP_INV_G11
XG1616 XI11_7/XI0/XI0_23/d_5_ XI11_7/XI0/XI0_23/d__5_ DECAP_INV_G11
XG1617 XI11_7/XI0/XI0_23/d_4_ XI11_7/XI0/XI0_23/d__4_ DECAP_INV_G11
XG1618 XI11_7/XI0/XI0_23/d_3_ XI11_7/XI0/XI0_23/d__3_ DECAP_INV_G11
XG1619 XI11_7/XI0/XI0_23/d_2_ XI11_7/XI0/XI0_23/d__2_ DECAP_INV_G11
XG1620 XI11_7/XI0/XI0_23/d_1_ XI11_7/XI0/XI0_23/d__1_ DECAP_INV_G11
XG1621 XI11_7/XI0/XI0_23/d_0_ XI11_7/XI0/XI0_23/d__0_ DECAP_INV_G11
XG1622 XI11_7/XI0/XI0_22/d__15_ XI11_7/XI0/XI0_22/d_15_ DECAP_INV_G11
XG1623 XI11_7/XI0/XI0_22/d__14_ XI11_7/XI0/XI0_22/d_14_ DECAP_INV_G11
XG1624 XI11_7/XI0/XI0_22/d__13_ XI11_7/XI0/XI0_22/d_13_ DECAP_INV_G11
XG1625 XI11_7/XI0/XI0_22/d__12_ XI11_7/XI0/XI0_22/d_12_ DECAP_INV_G11
XG1626 XI11_7/XI0/XI0_22/d__11_ XI11_7/XI0/XI0_22/d_11_ DECAP_INV_G11
XG1627 XI11_7/XI0/XI0_22/d__10_ XI11_7/XI0/XI0_22/d_10_ DECAP_INV_G11
XG1628 XI11_7/XI0/XI0_22/d__9_ XI11_7/XI0/XI0_22/d_9_ DECAP_INV_G11
XG1629 XI11_7/XI0/XI0_22/d__8_ XI11_7/XI0/XI0_22/d_8_ DECAP_INV_G11
XG1630 XI11_7/XI0/XI0_22/d__7_ XI11_7/XI0/XI0_22/d_7_ DECAP_INV_G11
XG1631 XI11_7/XI0/XI0_22/d__6_ XI11_7/XI0/XI0_22/d_6_ DECAP_INV_G11
XG1632 XI11_7/XI0/XI0_22/d__5_ XI11_7/XI0/XI0_22/d_5_ DECAP_INV_G11
XG1633 XI11_7/XI0/XI0_22/d__4_ XI11_7/XI0/XI0_22/d_4_ DECAP_INV_G11
XG1634 XI11_7/XI0/XI0_22/d__3_ XI11_7/XI0/XI0_22/d_3_ DECAP_INV_G11
XG1635 XI11_7/XI0/XI0_22/d__2_ XI11_7/XI0/XI0_22/d_2_ DECAP_INV_G11
XG1636 XI11_7/XI0/XI0_22/d__1_ XI11_7/XI0/XI0_22/d_1_ DECAP_INV_G11
XG1637 XI11_7/XI0/XI0_22/d__0_ XI11_7/XI0/XI0_22/d_0_ DECAP_INV_G11
XG1638 XI11_7/XI0/XI0_22/d_15_ XI11_7/XI0/XI0_22/d__15_ DECAP_INV_G11
XG1639 XI11_7/XI0/XI0_22/d_14_ XI11_7/XI0/XI0_22/d__14_ DECAP_INV_G11
XG1640 XI11_7/XI0/XI0_22/d_13_ XI11_7/XI0/XI0_22/d__13_ DECAP_INV_G11
XG1641 XI11_7/XI0/XI0_22/d_12_ XI11_7/XI0/XI0_22/d__12_ DECAP_INV_G11
XG1642 XI11_7/XI0/XI0_22/d_11_ XI11_7/XI0/XI0_22/d__11_ DECAP_INV_G11
XG1643 XI11_7/XI0/XI0_22/d_10_ XI11_7/XI0/XI0_22/d__10_ DECAP_INV_G11
XG1644 XI11_7/XI0/XI0_22/d_9_ XI11_7/XI0/XI0_22/d__9_ DECAP_INV_G11
XG1645 XI11_7/XI0/XI0_22/d_8_ XI11_7/XI0/XI0_22/d__8_ DECAP_INV_G11
XG1646 XI11_7/XI0/XI0_22/d_7_ XI11_7/XI0/XI0_22/d__7_ DECAP_INV_G11
XG1647 XI11_7/XI0/XI0_22/d_6_ XI11_7/XI0/XI0_22/d__6_ DECAP_INV_G11
XG1648 XI11_7/XI0/XI0_22/d_5_ XI11_7/XI0/XI0_22/d__5_ DECAP_INV_G11
XG1649 XI11_7/XI0/XI0_22/d_4_ XI11_7/XI0/XI0_22/d__4_ DECAP_INV_G11
XG1650 XI11_7/XI0/XI0_22/d_3_ XI11_7/XI0/XI0_22/d__3_ DECAP_INV_G11
XG1651 XI11_7/XI0/XI0_22/d_2_ XI11_7/XI0/XI0_22/d__2_ DECAP_INV_G11
XG1652 XI11_7/XI0/XI0_22/d_1_ XI11_7/XI0/XI0_22/d__1_ DECAP_INV_G11
XG1653 XI11_7/XI0/XI0_22/d_0_ XI11_7/XI0/XI0_22/d__0_ DECAP_INV_G11
XG1654 XI11_7/XI0/XI0_21/d__15_ XI11_7/XI0/XI0_21/d_15_ DECAP_INV_G11
XG1655 XI11_7/XI0/XI0_21/d__14_ XI11_7/XI0/XI0_21/d_14_ DECAP_INV_G11
XG1656 XI11_7/XI0/XI0_21/d__13_ XI11_7/XI0/XI0_21/d_13_ DECAP_INV_G11
XG1657 XI11_7/XI0/XI0_21/d__12_ XI11_7/XI0/XI0_21/d_12_ DECAP_INV_G11
XG1658 XI11_7/XI0/XI0_21/d__11_ XI11_7/XI0/XI0_21/d_11_ DECAP_INV_G11
XG1659 XI11_7/XI0/XI0_21/d__10_ XI11_7/XI0/XI0_21/d_10_ DECAP_INV_G11
XG1660 XI11_7/XI0/XI0_21/d__9_ XI11_7/XI0/XI0_21/d_9_ DECAP_INV_G11
XG1661 XI11_7/XI0/XI0_21/d__8_ XI11_7/XI0/XI0_21/d_8_ DECAP_INV_G11
XG1662 XI11_7/XI0/XI0_21/d__7_ XI11_7/XI0/XI0_21/d_7_ DECAP_INV_G11
XG1663 XI11_7/XI0/XI0_21/d__6_ XI11_7/XI0/XI0_21/d_6_ DECAP_INV_G11
XG1664 XI11_7/XI0/XI0_21/d__5_ XI11_7/XI0/XI0_21/d_5_ DECAP_INV_G11
XG1665 XI11_7/XI0/XI0_21/d__4_ XI11_7/XI0/XI0_21/d_4_ DECAP_INV_G11
XG1666 XI11_7/XI0/XI0_21/d__3_ XI11_7/XI0/XI0_21/d_3_ DECAP_INV_G11
XG1667 XI11_7/XI0/XI0_21/d__2_ XI11_7/XI0/XI0_21/d_2_ DECAP_INV_G11
XG1668 XI11_7/XI0/XI0_21/d__1_ XI11_7/XI0/XI0_21/d_1_ DECAP_INV_G11
XG1669 XI11_7/XI0/XI0_21/d__0_ XI11_7/XI0/XI0_21/d_0_ DECAP_INV_G11
XG1670 XI11_7/XI0/XI0_21/d_15_ XI11_7/XI0/XI0_21/d__15_ DECAP_INV_G11
XG1671 XI11_7/XI0/XI0_21/d_14_ XI11_7/XI0/XI0_21/d__14_ DECAP_INV_G11
XG1672 XI11_7/XI0/XI0_21/d_13_ XI11_7/XI0/XI0_21/d__13_ DECAP_INV_G11
XG1673 XI11_7/XI0/XI0_21/d_12_ XI11_7/XI0/XI0_21/d__12_ DECAP_INV_G11
XG1674 XI11_7/XI0/XI0_21/d_11_ XI11_7/XI0/XI0_21/d__11_ DECAP_INV_G11
XG1675 XI11_7/XI0/XI0_21/d_10_ XI11_7/XI0/XI0_21/d__10_ DECAP_INV_G11
XG1676 XI11_7/XI0/XI0_21/d_9_ XI11_7/XI0/XI0_21/d__9_ DECAP_INV_G11
XG1677 XI11_7/XI0/XI0_21/d_8_ XI11_7/XI0/XI0_21/d__8_ DECAP_INV_G11
XG1678 XI11_7/XI0/XI0_21/d_7_ XI11_7/XI0/XI0_21/d__7_ DECAP_INV_G11
XG1679 XI11_7/XI0/XI0_21/d_6_ XI11_7/XI0/XI0_21/d__6_ DECAP_INV_G11
XG1680 XI11_7/XI0/XI0_21/d_5_ XI11_7/XI0/XI0_21/d__5_ DECAP_INV_G11
XG1681 XI11_7/XI0/XI0_21/d_4_ XI11_7/XI0/XI0_21/d__4_ DECAP_INV_G11
XG1682 XI11_7/XI0/XI0_21/d_3_ XI11_7/XI0/XI0_21/d__3_ DECAP_INV_G11
XG1683 XI11_7/XI0/XI0_21/d_2_ XI11_7/XI0/XI0_21/d__2_ DECAP_INV_G11
XG1684 XI11_7/XI0/XI0_21/d_1_ XI11_7/XI0/XI0_21/d__1_ DECAP_INV_G11
XG1685 XI11_7/XI0/XI0_21/d_0_ XI11_7/XI0/XI0_21/d__0_ DECAP_INV_G11
XG1686 XI11_7/XI0/XI0_20/d__15_ XI11_7/XI0/XI0_20/d_15_ DECAP_INV_G11
XG1687 XI11_7/XI0/XI0_20/d__14_ XI11_7/XI0/XI0_20/d_14_ DECAP_INV_G11
XG1688 XI11_7/XI0/XI0_20/d__13_ XI11_7/XI0/XI0_20/d_13_ DECAP_INV_G11
XG1689 XI11_7/XI0/XI0_20/d__12_ XI11_7/XI0/XI0_20/d_12_ DECAP_INV_G11
XG1690 XI11_7/XI0/XI0_20/d__11_ XI11_7/XI0/XI0_20/d_11_ DECAP_INV_G11
XG1691 XI11_7/XI0/XI0_20/d__10_ XI11_7/XI0/XI0_20/d_10_ DECAP_INV_G11
XG1692 XI11_7/XI0/XI0_20/d__9_ XI11_7/XI0/XI0_20/d_9_ DECAP_INV_G11
XG1693 XI11_7/XI0/XI0_20/d__8_ XI11_7/XI0/XI0_20/d_8_ DECAP_INV_G11
XG1694 XI11_7/XI0/XI0_20/d__7_ XI11_7/XI0/XI0_20/d_7_ DECAP_INV_G11
XG1695 XI11_7/XI0/XI0_20/d__6_ XI11_7/XI0/XI0_20/d_6_ DECAP_INV_G11
XG1696 XI11_7/XI0/XI0_20/d__5_ XI11_7/XI0/XI0_20/d_5_ DECAP_INV_G11
XG1697 XI11_7/XI0/XI0_20/d__4_ XI11_7/XI0/XI0_20/d_4_ DECAP_INV_G11
XG1698 XI11_7/XI0/XI0_20/d__3_ XI11_7/XI0/XI0_20/d_3_ DECAP_INV_G11
XG1699 XI11_7/XI0/XI0_20/d__2_ XI11_7/XI0/XI0_20/d_2_ DECAP_INV_G11
XG1700 XI11_7/XI0/XI0_20/d__1_ XI11_7/XI0/XI0_20/d_1_ DECAP_INV_G11
XG1701 XI11_7/XI0/XI0_20/d__0_ XI11_7/XI0/XI0_20/d_0_ DECAP_INV_G11
XG1702 XI11_7/XI0/XI0_20/d_15_ XI11_7/XI0/XI0_20/d__15_ DECAP_INV_G11
XG1703 XI11_7/XI0/XI0_20/d_14_ XI11_7/XI0/XI0_20/d__14_ DECAP_INV_G11
XG1704 XI11_7/XI0/XI0_20/d_13_ XI11_7/XI0/XI0_20/d__13_ DECAP_INV_G11
XG1705 XI11_7/XI0/XI0_20/d_12_ XI11_7/XI0/XI0_20/d__12_ DECAP_INV_G11
XG1706 XI11_7/XI0/XI0_20/d_11_ XI11_7/XI0/XI0_20/d__11_ DECAP_INV_G11
XG1707 XI11_7/XI0/XI0_20/d_10_ XI11_7/XI0/XI0_20/d__10_ DECAP_INV_G11
XG1708 XI11_7/XI0/XI0_20/d_9_ XI11_7/XI0/XI0_20/d__9_ DECAP_INV_G11
XG1709 XI11_7/XI0/XI0_20/d_8_ XI11_7/XI0/XI0_20/d__8_ DECAP_INV_G11
XG1710 XI11_7/XI0/XI0_20/d_7_ XI11_7/XI0/XI0_20/d__7_ DECAP_INV_G11
XG1711 XI11_7/XI0/XI0_20/d_6_ XI11_7/XI0/XI0_20/d__6_ DECAP_INV_G11
XG1712 XI11_7/XI0/XI0_20/d_5_ XI11_7/XI0/XI0_20/d__5_ DECAP_INV_G11
XG1713 XI11_7/XI0/XI0_20/d_4_ XI11_7/XI0/XI0_20/d__4_ DECAP_INV_G11
XG1714 XI11_7/XI0/XI0_20/d_3_ XI11_7/XI0/XI0_20/d__3_ DECAP_INV_G11
XG1715 XI11_7/XI0/XI0_20/d_2_ XI11_7/XI0/XI0_20/d__2_ DECAP_INV_G11
XG1716 XI11_7/XI0/XI0_20/d_1_ XI11_7/XI0/XI0_20/d__1_ DECAP_INV_G11
XG1717 XI11_7/XI0/XI0_20/d_0_ XI11_7/XI0/XI0_20/d__0_ DECAP_INV_G11
XG1718 XI11_7/XI0/XI0_19/d__15_ XI11_7/XI0/XI0_19/d_15_ DECAP_INV_G11
XG1719 XI11_7/XI0/XI0_19/d__14_ XI11_7/XI0/XI0_19/d_14_ DECAP_INV_G11
XG1720 XI11_7/XI0/XI0_19/d__13_ XI11_7/XI0/XI0_19/d_13_ DECAP_INV_G11
XG1721 XI11_7/XI0/XI0_19/d__12_ XI11_7/XI0/XI0_19/d_12_ DECAP_INV_G11
XG1722 XI11_7/XI0/XI0_19/d__11_ XI11_7/XI0/XI0_19/d_11_ DECAP_INV_G11
XG1723 XI11_7/XI0/XI0_19/d__10_ XI11_7/XI0/XI0_19/d_10_ DECAP_INV_G11
XG1724 XI11_7/XI0/XI0_19/d__9_ XI11_7/XI0/XI0_19/d_9_ DECAP_INV_G11
XG1725 XI11_7/XI0/XI0_19/d__8_ XI11_7/XI0/XI0_19/d_8_ DECAP_INV_G11
XG1726 XI11_7/XI0/XI0_19/d__7_ XI11_7/XI0/XI0_19/d_7_ DECAP_INV_G11
XG1727 XI11_7/XI0/XI0_19/d__6_ XI11_7/XI0/XI0_19/d_6_ DECAP_INV_G11
XG1728 XI11_7/XI0/XI0_19/d__5_ XI11_7/XI0/XI0_19/d_5_ DECAP_INV_G11
XG1729 XI11_7/XI0/XI0_19/d__4_ XI11_7/XI0/XI0_19/d_4_ DECAP_INV_G11
XG1730 XI11_7/XI0/XI0_19/d__3_ XI11_7/XI0/XI0_19/d_3_ DECAP_INV_G11
XG1731 XI11_7/XI0/XI0_19/d__2_ XI11_7/XI0/XI0_19/d_2_ DECAP_INV_G11
XG1732 XI11_7/XI0/XI0_19/d__1_ XI11_7/XI0/XI0_19/d_1_ DECAP_INV_G11
XG1733 XI11_7/XI0/XI0_19/d__0_ XI11_7/XI0/XI0_19/d_0_ DECAP_INV_G11
XG1734 XI11_7/XI0/XI0_19/d_15_ XI11_7/XI0/XI0_19/d__15_ DECAP_INV_G11
XG1735 XI11_7/XI0/XI0_19/d_14_ XI11_7/XI0/XI0_19/d__14_ DECAP_INV_G11
XG1736 XI11_7/XI0/XI0_19/d_13_ XI11_7/XI0/XI0_19/d__13_ DECAP_INV_G11
XG1737 XI11_7/XI0/XI0_19/d_12_ XI11_7/XI0/XI0_19/d__12_ DECAP_INV_G11
XG1738 XI11_7/XI0/XI0_19/d_11_ XI11_7/XI0/XI0_19/d__11_ DECAP_INV_G11
XG1739 XI11_7/XI0/XI0_19/d_10_ XI11_7/XI0/XI0_19/d__10_ DECAP_INV_G11
XG1740 XI11_7/XI0/XI0_19/d_9_ XI11_7/XI0/XI0_19/d__9_ DECAP_INV_G11
XG1741 XI11_7/XI0/XI0_19/d_8_ XI11_7/XI0/XI0_19/d__8_ DECAP_INV_G11
XG1742 XI11_7/XI0/XI0_19/d_7_ XI11_7/XI0/XI0_19/d__7_ DECAP_INV_G11
XG1743 XI11_7/XI0/XI0_19/d_6_ XI11_7/XI0/XI0_19/d__6_ DECAP_INV_G11
XG1744 XI11_7/XI0/XI0_19/d_5_ XI11_7/XI0/XI0_19/d__5_ DECAP_INV_G11
XG1745 XI11_7/XI0/XI0_19/d_4_ XI11_7/XI0/XI0_19/d__4_ DECAP_INV_G11
XG1746 XI11_7/XI0/XI0_19/d_3_ XI11_7/XI0/XI0_19/d__3_ DECAP_INV_G11
XG1747 XI11_7/XI0/XI0_19/d_2_ XI11_7/XI0/XI0_19/d__2_ DECAP_INV_G11
XG1748 XI11_7/XI0/XI0_19/d_1_ XI11_7/XI0/XI0_19/d__1_ DECAP_INV_G11
XG1749 XI11_7/XI0/XI0_19/d_0_ XI11_7/XI0/XI0_19/d__0_ DECAP_INV_G11
XG1750 XI11_7/XI0/XI0_18/d__15_ XI11_7/XI0/XI0_18/d_15_ DECAP_INV_G11
XG1751 XI11_7/XI0/XI0_18/d__14_ XI11_7/XI0/XI0_18/d_14_ DECAP_INV_G11
XG1752 XI11_7/XI0/XI0_18/d__13_ XI11_7/XI0/XI0_18/d_13_ DECAP_INV_G11
XG1753 XI11_7/XI0/XI0_18/d__12_ XI11_7/XI0/XI0_18/d_12_ DECAP_INV_G11
XG1754 XI11_7/XI0/XI0_18/d__11_ XI11_7/XI0/XI0_18/d_11_ DECAP_INV_G11
XG1755 XI11_7/XI0/XI0_18/d__10_ XI11_7/XI0/XI0_18/d_10_ DECAP_INV_G11
XG1756 XI11_7/XI0/XI0_18/d__9_ XI11_7/XI0/XI0_18/d_9_ DECAP_INV_G11
XG1757 XI11_7/XI0/XI0_18/d__8_ XI11_7/XI0/XI0_18/d_8_ DECAP_INV_G11
XG1758 XI11_7/XI0/XI0_18/d__7_ XI11_7/XI0/XI0_18/d_7_ DECAP_INV_G11
XG1759 XI11_7/XI0/XI0_18/d__6_ XI11_7/XI0/XI0_18/d_6_ DECAP_INV_G11
XG1760 XI11_7/XI0/XI0_18/d__5_ XI11_7/XI0/XI0_18/d_5_ DECAP_INV_G11
XG1761 XI11_7/XI0/XI0_18/d__4_ XI11_7/XI0/XI0_18/d_4_ DECAP_INV_G11
XG1762 XI11_7/XI0/XI0_18/d__3_ XI11_7/XI0/XI0_18/d_3_ DECAP_INV_G11
XG1763 XI11_7/XI0/XI0_18/d__2_ XI11_7/XI0/XI0_18/d_2_ DECAP_INV_G11
XG1764 XI11_7/XI0/XI0_18/d__1_ XI11_7/XI0/XI0_18/d_1_ DECAP_INV_G11
XG1765 XI11_7/XI0/XI0_18/d__0_ XI11_7/XI0/XI0_18/d_0_ DECAP_INV_G11
XG1766 XI11_7/XI0/XI0_18/d_15_ XI11_7/XI0/XI0_18/d__15_ DECAP_INV_G11
XG1767 XI11_7/XI0/XI0_18/d_14_ XI11_7/XI0/XI0_18/d__14_ DECAP_INV_G11
XG1768 XI11_7/XI0/XI0_18/d_13_ XI11_7/XI0/XI0_18/d__13_ DECAP_INV_G11
XG1769 XI11_7/XI0/XI0_18/d_12_ XI11_7/XI0/XI0_18/d__12_ DECAP_INV_G11
XG1770 XI11_7/XI0/XI0_18/d_11_ XI11_7/XI0/XI0_18/d__11_ DECAP_INV_G11
XG1771 XI11_7/XI0/XI0_18/d_10_ XI11_7/XI0/XI0_18/d__10_ DECAP_INV_G11
XG1772 XI11_7/XI0/XI0_18/d_9_ XI11_7/XI0/XI0_18/d__9_ DECAP_INV_G11
XG1773 XI11_7/XI0/XI0_18/d_8_ XI11_7/XI0/XI0_18/d__8_ DECAP_INV_G11
XG1774 XI11_7/XI0/XI0_18/d_7_ XI11_7/XI0/XI0_18/d__7_ DECAP_INV_G11
XG1775 XI11_7/XI0/XI0_18/d_6_ XI11_7/XI0/XI0_18/d__6_ DECAP_INV_G11
XG1776 XI11_7/XI0/XI0_18/d_5_ XI11_7/XI0/XI0_18/d__5_ DECAP_INV_G11
XG1777 XI11_7/XI0/XI0_18/d_4_ XI11_7/XI0/XI0_18/d__4_ DECAP_INV_G11
XG1778 XI11_7/XI0/XI0_18/d_3_ XI11_7/XI0/XI0_18/d__3_ DECAP_INV_G11
XG1779 XI11_7/XI0/XI0_18/d_2_ XI11_7/XI0/XI0_18/d__2_ DECAP_INV_G11
XG1780 XI11_7/XI0/XI0_18/d_1_ XI11_7/XI0/XI0_18/d__1_ DECAP_INV_G11
XG1781 XI11_7/XI0/XI0_18/d_0_ XI11_7/XI0/XI0_18/d__0_ DECAP_INV_G11
XG1782 XI11_7/XI0/XI0_17/d__15_ XI11_7/XI0/XI0_17/d_15_ DECAP_INV_G11
XG1783 XI11_7/XI0/XI0_17/d__14_ XI11_7/XI0/XI0_17/d_14_ DECAP_INV_G11
XG1784 XI11_7/XI0/XI0_17/d__13_ XI11_7/XI0/XI0_17/d_13_ DECAP_INV_G11
XG1785 XI11_7/XI0/XI0_17/d__12_ XI11_7/XI0/XI0_17/d_12_ DECAP_INV_G11
XG1786 XI11_7/XI0/XI0_17/d__11_ XI11_7/XI0/XI0_17/d_11_ DECAP_INV_G11
XG1787 XI11_7/XI0/XI0_17/d__10_ XI11_7/XI0/XI0_17/d_10_ DECAP_INV_G11
XG1788 XI11_7/XI0/XI0_17/d__9_ XI11_7/XI0/XI0_17/d_9_ DECAP_INV_G11
XG1789 XI11_7/XI0/XI0_17/d__8_ XI11_7/XI0/XI0_17/d_8_ DECAP_INV_G11
XG1790 XI11_7/XI0/XI0_17/d__7_ XI11_7/XI0/XI0_17/d_7_ DECAP_INV_G11
XG1791 XI11_7/XI0/XI0_17/d__6_ XI11_7/XI0/XI0_17/d_6_ DECAP_INV_G11
XG1792 XI11_7/XI0/XI0_17/d__5_ XI11_7/XI0/XI0_17/d_5_ DECAP_INV_G11
XG1793 XI11_7/XI0/XI0_17/d__4_ XI11_7/XI0/XI0_17/d_4_ DECAP_INV_G11
XG1794 XI11_7/XI0/XI0_17/d__3_ XI11_7/XI0/XI0_17/d_3_ DECAP_INV_G11
XG1795 XI11_7/XI0/XI0_17/d__2_ XI11_7/XI0/XI0_17/d_2_ DECAP_INV_G11
XG1796 XI11_7/XI0/XI0_17/d__1_ XI11_7/XI0/XI0_17/d_1_ DECAP_INV_G11
XG1797 XI11_7/XI0/XI0_17/d__0_ XI11_7/XI0/XI0_17/d_0_ DECAP_INV_G11
XG1798 XI11_7/XI0/XI0_17/d_15_ XI11_7/XI0/XI0_17/d__15_ DECAP_INV_G11
XG1799 XI11_7/XI0/XI0_17/d_14_ XI11_7/XI0/XI0_17/d__14_ DECAP_INV_G11
XG1800 XI11_7/XI0/XI0_17/d_13_ XI11_7/XI0/XI0_17/d__13_ DECAP_INV_G11
XG1801 XI11_7/XI0/XI0_17/d_12_ XI11_7/XI0/XI0_17/d__12_ DECAP_INV_G11
XG1802 XI11_7/XI0/XI0_17/d_11_ XI11_7/XI0/XI0_17/d__11_ DECAP_INV_G11
XG1803 XI11_7/XI0/XI0_17/d_10_ XI11_7/XI0/XI0_17/d__10_ DECAP_INV_G11
XG1804 XI11_7/XI0/XI0_17/d_9_ XI11_7/XI0/XI0_17/d__9_ DECAP_INV_G11
XG1805 XI11_7/XI0/XI0_17/d_8_ XI11_7/XI0/XI0_17/d__8_ DECAP_INV_G11
XG1806 XI11_7/XI0/XI0_17/d_7_ XI11_7/XI0/XI0_17/d__7_ DECAP_INV_G11
XG1807 XI11_7/XI0/XI0_17/d_6_ XI11_7/XI0/XI0_17/d__6_ DECAP_INV_G11
XG1808 XI11_7/XI0/XI0_17/d_5_ XI11_7/XI0/XI0_17/d__5_ DECAP_INV_G11
XG1809 XI11_7/XI0/XI0_17/d_4_ XI11_7/XI0/XI0_17/d__4_ DECAP_INV_G11
XG1810 XI11_7/XI0/XI0_17/d_3_ XI11_7/XI0/XI0_17/d__3_ DECAP_INV_G11
XG1811 XI11_7/XI0/XI0_17/d_2_ XI11_7/XI0/XI0_17/d__2_ DECAP_INV_G11
XG1812 XI11_7/XI0/XI0_17/d_1_ XI11_7/XI0/XI0_17/d__1_ DECAP_INV_G11
XG1813 XI11_7/XI0/XI0_17/d_0_ XI11_7/XI0/XI0_17/d__0_ DECAP_INV_G11
XG1814 XI11_7/XI0/XI0_16/d__15_ XI11_7/XI0/XI0_16/d_15_ DECAP_INV_G11
XG1815 XI11_7/XI0/XI0_16/d__14_ XI11_7/XI0/XI0_16/d_14_ DECAP_INV_G11
XG1816 XI11_7/XI0/XI0_16/d__13_ XI11_7/XI0/XI0_16/d_13_ DECAP_INV_G11
XG1817 XI11_7/XI0/XI0_16/d__12_ XI11_7/XI0/XI0_16/d_12_ DECAP_INV_G11
XG1818 XI11_7/XI0/XI0_16/d__11_ XI11_7/XI0/XI0_16/d_11_ DECAP_INV_G11
XG1819 XI11_7/XI0/XI0_16/d__10_ XI11_7/XI0/XI0_16/d_10_ DECAP_INV_G11
XG1820 XI11_7/XI0/XI0_16/d__9_ XI11_7/XI0/XI0_16/d_9_ DECAP_INV_G11
XG1821 XI11_7/XI0/XI0_16/d__8_ XI11_7/XI0/XI0_16/d_8_ DECAP_INV_G11
XG1822 XI11_7/XI0/XI0_16/d__7_ XI11_7/XI0/XI0_16/d_7_ DECAP_INV_G11
XG1823 XI11_7/XI0/XI0_16/d__6_ XI11_7/XI0/XI0_16/d_6_ DECAP_INV_G11
XG1824 XI11_7/XI0/XI0_16/d__5_ XI11_7/XI0/XI0_16/d_5_ DECAP_INV_G11
XG1825 XI11_7/XI0/XI0_16/d__4_ XI11_7/XI0/XI0_16/d_4_ DECAP_INV_G11
XG1826 XI11_7/XI0/XI0_16/d__3_ XI11_7/XI0/XI0_16/d_3_ DECAP_INV_G11
XG1827 XI11_7/XI0/XI0_16/d__2_ XI11_7/XI0/XI0_16/d_2_ DECAP_INV_G11
XG1828 XI11_7/XI0/XI0_16/d__1_ XI11_7/XI0/XI0_16/d_1_ DECAP_INV_G11
XG1829 XI11_7/XI0/XI0_16/d__0_ XI11_7/XI0/XI0_16/d_0_ DECAP_INV_G11
XG1830 XI11_7/XI0/XI0_16/d_15_ XI11_7/XI0/XI0_16/d__15_ DECAP_INV_G11
XG1831 XI11_7/XI0/XI0_16/d_14_ XI11_7/XI0/XI0_16/d__14_ DECAP_INV_G11
XG1832 XI11_7/XI0/XI0_16/d_13_ XI11_7/XI0/XI0_16/d__13_ DECAP_INV_G11
XG1833 XI11_7/XI0/XI0_16/d_12_ XI11_7/XI0/XI0_16/d__12_ DECAP_INV_G11
XG1834 XI11_7/XI0/XI0_16/d_11_ XI11_7/XI0/XI0_16/d__11_ DECAP_INV_G11
XG1835 XI11_7/XI0/XI0_16/d_10_ XI11_7/XI0/XI0_16/d__10_ DECAP_INV_G11
XG1836 XI11_7/XI0/XI0_16/d_9_ XI11_7/XI0/XI0_16/d__9_ DECAP_INV_G11
XG1837 XI11_7/XI0/XI0_16/d_8_ XI11_7/XI0/XI0_16/d__8_ DECAP_INV_G11
XG1838 XI11_7/XI0/XI0_16/d_7_ XI11_7/XI0/XI0_16/d__7_ DECAP_INV_G11
XG1839 XI11_7/XI0/XI0_16/d_6_ XI11_7/XI0/XI0_16/d__6_ DECAP_INV_G11
XG1840 XI11_7/XI0/XI0_16/d_5_ XI11_7/XI0/XI0_16/d__5_ DECAP_INV_G11
XG1841 XI11_7/XI0/XI0_16/d_4_ XI11_7/XI0/XI0_16/d__4_ DECAP_INV_G11
XG1842 XI11_7/XI0/XI0_16/d_3_ XI11_7/XI0/XI0_16/d__3_ DECAP_INV_G11
XG1843 XI11_7/XI0/XI0_16/d_2_ XI11_7/XI0/XI0_16/d__2_ DECAP_INV_G11
XG1844 XI11_7/XI0/XI0_16/d_1_ XI11_7/XI0/XI0_16/d__1_ DECAP_INV_G11
XG1845 XI11_7/XI0/XI0_16/d_0_ XI11_7/XI0/XI0_16/d__0_ DECAP_INV_G11
XG1846 XI11_7/XI0/XI0_15/d__15_ XI11_7/XI0/XI0_15/d_15_ DECAP_INV_G11
XG1847 XI11_7/XI0/XI0_15/d__14_ XI11_7/XI0/XI0_15/d_14_ DECAP_INV_G11
XG1848 XI11_7/XI0/XI0_15/d__13_ XI11_7/XI0/XI0_15/d_13_ DECAP_INV_G11
XG1849 XI11_7/XI0/XI0_15/d__12_ XI11_7/XI0/XI0_15/d_12_ DECAP_INV_G11
XG1850 XI11_7/XI0/XI0_15/d__11_ XI11_7/XI0/XI0_15/d_11_ DECAP_INV_G11
XG1851 XI11_7/XI0/XI0_15/d__10_ XI11_7/XI0/XI0_15/d_10_ DECAP_INV_G11
XG1852 XI11_7/XI0/XI0_15/d__9_ XI11_7/XI0/XI0_15/d_9_ DECAP_INV_G11
XG1853 XI11_7/XI0/XI0_15/d__8_ XI11_7/XI0/XI0_15/d_8_ DECAP_INV_G11
XG1854 XI11_7/XI0/XI0_15/d__7_ XI11_7/XI0/XI0_15/d_7_ DECAP_INV_G11
XG1855 XI11_7/XI0/XI0_15/d__6_ XI11_7/XI0/XI0_15/d_6_ DECAP_INV_G11
XG1856 XI11_7/XI0/XI0_15/d__5_ XI11_7/XI0/XI0_15/d_5_ DECAP_INV_G11
XG1857 XI11_7/XI0/XI0_15/d__4_ XI11_7/XI0/XI0_15/d_4_ DECAP_INV_G11
XG1858 XI11_7/XI0/XI0_15/d__3_ XI11_7/XI0/XI0_15/d_3_ DECAP_INV_G11
XG1859 XI11_7/XI0/XI0_15/d__2_ XI11_7/XI0/XI0_15/d_2_ DECAP_INV_G11
XG1860 XI11_7/XI0/XI0_15/d__1_ XI11_7/XI0/XI0_15/d_1_ DECAP_INV_G11
XG1861 XI11_7/XI0/XI0_15/d__0_ XI11_7/XI0/XI0_15/d_0_ DECAP_INV_G11
XG1862 XI11_7/XI0/XI0_15/d_15_ XI11_7/XI0/XI0_15/d__15_ DECAP_INV_G11
XG1863 XI11_7/XI0/XI0_15/d_14_ XI11_7/XI0/XI0_15/d__14_ DECAP_INV_G11
XG1864 XI11_7/XI0/XI0_15/d_13_ XI11_7/XI0/XI0_15/d__13_ DECAP_INV_G11
XG1865 XI11_7/XI0/XI0_15/d_12_ XI11_7/XI0/XI0_15/d__12_ DECAP_INV_G11
XG1866 XI11_7/XI0/XI0_15/d_11_ XI11_7/XI0/XI0_15/d__11_ DECAP_INV_G11
XG1867 XI11_7/XI0/XI0_15/d_10_ XI11_7/XI0/XI0_15/d__10_ DECAP_INV_G11
XG1868 XI11_7/XI0/XI0_15/d_9_ XI11_7/XI0/XI0_15/d__9_ DECAP_INV_G11
XG1869 XI11_7/XI0/XI0_15/d_8_ XI11_7/XI0/XI0_15/d__8_ DECAP_INV_G11
XG1870 XI11_7/XI0/XI0_15/d_7_ XI11_7/XI0/XI0_15/d__7_ DECAP_INV_G11
XG1871 XI11_7/XI0/XI0_15/d_6_ XI11_7/XI0/XI0_15/d__6_ DECAP_INV_G11
XG1872 XI11_7/XI0/XI0_15/d_5_ XI11_7/XI0/XI0_15/d__5_ DECAP_INV_G11
XG1873 XI11_7/XI0/XI0_15/d_4_ XI11_7/XI0/XI0_15/d__4_ DECAP_INV_G11
XG1874 XI11_7/XI0/XI0_15/d_3_ XI11_7/XI0/XI0_15/d__3_ DECAP_INV_G11
XG1875 XI11_7/XI0/XI0_15/d_2_ XI11_7/XI0/XI0_15/d__2_ DECAP_INV_G11
XG1876 XI11_7/XI0/XI0_15/d_1_ XI11_7/XI0/XI0_15/d__1_ DECAP_INV_G11
XG1877 XI11_7/XI0/XI0_15/d_0_ XI11_7/XI0/XI0_15/d__0_ DECAP_INV_G11
XG1878 XI11_7/XI0/XI0_14/d__15_ XI11_7/XI0/XI0_14/d_15_ DECAP_INV_G11
XG1879 XI11_7/XI0/XI0_14/d__14_ XI11_7/XI0/XI0_14/d_14_ DECAP_INV_G11
XG1880 XI11_7/XI0/XI0_14/d__13_ XI11_7/XI0/XI0_14/d_13_ DECAP_INV_G11
XG1881 XI11_7/XI0/XI0_14/d__12_ XI11_7/XI0/XI0_14/d_12_ DECAP_INV_G11
XG1882 XI11_7/XI0/XI0_14/d__11_ XI11_7/XI0/XI0_14/d_11_ DECAP_INV_G11
XG1883 XI11_7/XI0/XI0_14/d__10_ XI11_7/XI0/XI0_14/d_10_ DECAP_INV_G11
XG1884 XI11_7/XI0/XI0_14/d__9_ XI11_7/XI0/XI0_14/d_9_ DECAP_INV_G11
XG1885 XI11_7/XI0/XI0_14/d__8_ XI11_7/XI0/XI0_14/d_8_ DECAP_INV_G11
XG1886 XI11_7/XI0/XI0_14/d__7_ XI11_7/XI0/XI0_14/d_7_ DECAP_INV_G11
XG1887 XI11_7/XI0/XI0_14/d__6_ XI11_7/XI0/XI0_14/d_6_ DECAP_INV_G11
XG1888 XI11_7/XI0/XI0_14/d__5_ XI11_7/XI0/XI0_14/d_5_ DECAP_INV_G11
XG1889 XI11_7/XI0/XI0_14/d__4_ XI11_7/XI0/XI0_14/d_4_ DECAP_INV_G11
XG1890 XI11_7/XI0/XI0_14/d__3_ XI11_7/XI0/XI0_14/d_3_ DECAP_INV_G11
XG1891 XI11_7/XI0/XI0_14/d__2_ XI11_7/XI0/XI0_14/d_2_ DECAP_INV_G11
XG1892 XI11_7/XI0/XI0_14/d__1_ XI11_7/XI0/XI0_14/d_1_ DECAP_INV_G11
XG1893 XI11_7/XI0/XI0_14/d__0_ XI11_7/XI0/XI0_14/d_0_ DECAP_INV_G11
XG1894 XI11_7/XI0/XI0_14/d_15_ XI11_7/XI0/XI0_14/d__15_ DECAP_INV_G11
XG1895 XI11_7/XI0/XI0_14/d_14_ XI11_7/XI0/XI0_14/d__14_ DECAP_INV_G11
XG1896 XI11_7/XI0/XI0_14/d_13_ XI11_7/XI0/XI0_14/d__13_ DECAP_INV_G11
XG1897 XI11_7/XI0/XI0_14/d_12_ XI11_7/XI0/XI0_14/d__12_ DECAP_INV_G11
XG1898 XI11_7/XI0/XI0_14/d_11_ XI11_7/XI0/XI0_14/d__11_ DECAP_INV_G11
XG1899 XI11_7/XI0/XI0_14/d_10_ XI11_7/XI0/XI0_14/d__10_ DECAP_INV_G11
XG1900 XI11_7/XI0/XI0_14/d_9_ XI11_7/XI0/XI0_14/d__9_ DECAP_INV_G11
XG1901 XI11_7/XI0/XI0_14/d_8_ XI11_7/XI0/XI0_14/d__8_ DECAP_INV_G11
XG1902 XI11_7/XI0/XI0_14/d_7_ XI11_7/XI0/XI0_14/d__7_ DECAP_INV_G11
XG1903 XI11_7/XI0/XI0_14/d_6_ XI11_7/XI0/XI0_14/d__6_ DECAP_INV_G11
XG1904 XI11_7/XI0/XI0_14/d_5_ XI11_7/XI0/XI0_14/d__5_ DECAP_INV_G11
XG1905 XI11_7/XI0/XI0_14/d_4_ XI11_7/XI0/XI0_14/d__4_ DECAP_INV_G11
XG1906 XI11_7/XI0/XI0_14/d_3_ XI11_7/XI0/XI0_14/d__3_ DECAP_INV_G11
XG1907 XI11_7/XI0/XI0_14/d_2_ XI11_7/XI0/XI0_14/d__2_ DECAP_INV_G11
XG1908 XI11_7/XI0/XI0_14/d_1_ XI11_7/XI0/XI0_14/d__1_ DECAP_INV_G11
XG1909 XI11_7/XI0/XI0_14/d_0_ XI11_7/XI0/XI0_14/d__0_ DECAP_INV_G11
XG1910 XI11_7/XI0/XI0_13/d__15_ XI11_7/XI0/XI0_13/d_15_ DECAP_INV_G11
XG1911 XI11_7/XI0/XI0_13/d__14_ XI11_7/XI0/XI0_13/d_14_ DECAP_INV_G11
XG1912 XI11_7/XI0/XI0_13/d__13_ XI11_7/XI0/XI0_13/d_13_ DECAP_INV_G11
XG1913 XI11_7/XI0/XI0_13/d__12_ XI11_7/XI0/XI0_13/d_12_ DECAP_INV_G11
XG1914 XI11_7/XI0/XI0_13/d__11_ XI11_7/XI0/XI0_13/d_11_ DECAP_INV_G11
XG1915 XI11_7/XI0/XI0_13/d__10_ XI11_7/XI0/XI0_13/d_10_ DECAP_INV_G11
XG1916 XI11_7/XI0/XI0_13/d__9_ XI11_7/XI0/XI0_13/d_9_ DECAP_INV_G11
XG1917 XI11_7/XI0/XI0_13/d__8_ XI11_7/XI0/XI0_13/d_8_ DECAP_INV_G11
XG1918 XI11_7/XI0/XI0_13/d__7_ XI11_7/XI0/XI0_13/d_7_ DECAP_INV_G11
XG1919 XI11_7/XI0/XI0_13/d__6_ XI11_7/XI0/XI0_13/d_6_ DECAP_INV_G11
XG1920 XI11_7/XI0/XI0_13/d__5_ XI11_7/XI0/XI0_13/d_5_ DECAP_INV_G11
XG1921 XI11_7/XI0/XI0_13/d__4_ XI11_7/XI0/XI0_13/d_4_ DECAP_INV_G11
XG1922 XI11_7/XI0/XI0_13/d__3_ XI11_7/XI0/XI0_13/d_3_ DECAP_INV_G11
XG1923 XI11_7/XI0/XI0_13/d__2_ XI11_7/XI0/XI0_13/d_2_ DECAP_INV_G11
XG1924 XI11_7/XI0/XI0_13/d__1_ XI11_7/XI0/XI0_13/d_1_ DECAP_INV_G11
XG1925 XI11_7/XI0/XI0_13/d__0_ XI11_7/XI0/XI0_13/d_0_ DECAP_INV_G11
XG1926 XI11_7/XI0/XI0_13/d_15_ XI11_7/XI0/XI0_13/d__15_ DECAP_INV_G11
XG1927 XI11_7/XI0/XI0_13/d_14_ XI11_7/XI0/XI0_13/d__14_ DECAP_INV_G11
XG1928 XI11_7/XI0/XI0_13/d_13_ XI11_7/XI0/XI0_13/d__13_ DECAP_INV_G11
XG1929 XI11_7/XI0/XI0_13/d_12_ XI11_7/XI0/XI0_13/d__12_ DECAP_INV_G11
XG1930 XI11_7/XI0/XI0_13/d_11_ XI11_7/XI0/XI0_13/d__11_ DECAP_INV_G11
XG1931 XI11_7/XI0/XI0_13/d_10_ XI11_7/XI0/XI0_13/d__10_ DECAP_INV_G11
XG1932 XI11_7/XI0/XI0_13/d_9_ XI11_7/XI0/XI0_13/d__9_ DECAP_INV_G11
XG1933 XI11_7/XI0/XI0_13/d_8_ XI11_7/XI0/XI0_13/d__8_ DECAP_INV_G11
XG1934 XI11_7/XI0/XI0_13/d_7_ XI11_7/XI0/XI0_13/d__7_ DECAP_INV_G11
XG1935 XI11_7/XI0/XI0_13/d_6_ XI11_7/XI0/XI0_13/d__6_ DECAP_INV_G11
XG1936 XI11_7/XI0/XI0_13/d_5_ XI11_7/XI0/XI0_13/d__5_ DECAP_INV_G11
XG1937 XI11_7/XI0/XI0_13/d_4_ XI11_7/XI0/XI0_13/d__4_ DECAP_INV_G11
XG1938 XI11_7/XI0/XI0_13/d_3_ XI11_7/XI0/XI0_13/d__3_ DECAP_INV_G11
XG1939 XI11_7/XI0/XI0_13/d_2_ XI11_7/XI0/XI0_13/d__2_ DECAP_INV_G11
XG1940 XI11_7/XI0/XI0_13/d_1_ XI11_7/XI0/XI0_13/d__1_ DECAP_INV_G11
XG1941 XI11_7/XI0/XI0_13/d_0_ XI11_7/XI0/XI0_13/d__0_ DECAP_INV_G11
XG1942 XI11_7/XI0/XI0_12/d__15_ XI11_7/XI0/XI0_12/d_15_ DECAP_INV_G11
XG1943 XI11_7/XI0/XI0_12/d__14_ XI11_7/XI0/XI0_12/d_14_ DECAP_INV_G11
XG1944 XI11_7/XI0/XI0_12/d__13_ XI11_7/XI0/XI0_12/d_13_ DECAP_INV_G11
XG1945 XI11_7/XI0/XI0_12/d__12_ XI11_7/XI0/XI0_12/d_12_ DECAP_INV_G11
XG1946 XI11_7/XI0/XI0_12/d__11_ XI11_7/XI0/XI0_12/d_11_ DECAP_INV_G11
XG1947 XI11_7/XI0/XI0_12/d__10_ XI11_7/XI0/XI0_12/d_10_ DECAP_INV_G11
XG1948 XI11_7/XI0/XI0_12/d__9_ XI11_7/XI0/XI0_12/d_9_ DECAP_INV_G11
XG1949 XI11_7/XI0/XI0_12/d__8_ XI11_7/XI0/XI0_12/d_8_ DECAP_INV_G11
XG1950 XI11_7/XI0/XI0_12/d__7_ XI11_7/XI0/XI0_12/d_7_ DECAP_INV_G11
XG1951 XI11_7/XI0/XI0_12/d__6_ XI11_7/XI0/XI0_12/d_6_ DECAP_INV_G11
XG1952 XI11_7/XI0/XI0_12/d__5_ XI11_7/XI0/XI0_12/d_5_ DECAP_INV_G11
XG1953 XI11_7/XI0/XI0_12/d__4_ XI11_7/XI0/XI0_12/d_4_ DECAP_INV_G11
XG1954 XI11_7/XI0/XI0_12/d__3_ XI11_7/XI0/XI0_12/d_3_ DECAP_INV_G11
XG1955 XI11_7/XI0/XI0_12/d__2_ XI11_7/XI0/XI0_12/d_2_ DECAP_INV_G11
XG1956 XI11_7/XI0/XI0_12/d__1_ XI11_7/XI0/XI0_12/d_1_ DECAP_INV_G11
XG1957 XI11_7/XI0/XI0_12/d__0_ XI11_7/XI0/XI0_12/d_0_ DECAP_INV_G11
XG1958 XI11_7/XI0/XI0_12/d_15_ XI11_7/XI0/XI0_12/d__15_ DECAP_INV_G11
XG1959 XI11_7/XI0/XI0_12/d_14_ XI11_7/XI0/XI0_12/d__14_ DECAP_INV_G11
XG1960 XI11_7/XI0/XI0_12/d_13_ XI11_7/XI0/XI0_12/d__13_ DECAP_INV_G11
XG1961 XI11_7/XI0/XI0_12/d_12_ XI11_7/XI0/XI0_12/d__12_ DECAP_INV_G11
XG1962 XI11_7/XI0/XI0_12/d_11_ XI11_7/XI0/XI0_12/d__11_ DECAP_INV_G11
XG1963 XI11_7/XI0/XI0_12/d_10_ XI11_7/XI0/XI0_12/d__10_ DECAP_INV_G11
XG1964 XI11_7/XI0/XI0_12/d_9_ XI11_7/XI0/XI0_12/d__9_ DECAP_INV_G11
XG1965 XI11_7/XI0/XI0_12/d_8_ XI11_7/XI0/XI0_12/d__8_ DECAP_INV_G11
XG1966 XI11_7/XI0/XI0_12/d_7_ XI11_7/XI0/XI0_12/d__7_ DECAP_INV_G11
XG1967 XI11_7/XI0/XI0_12/d_6_ XI11_7/XI0/XI0_12/d__6_ DECAP_INV_G11
XG1968 XI11_7/XI0/XI0_12/d_5_ XI11_7/XI0/XI0_12/d__5_ DECAP_INV_G11
XG1969 XI11_7/XI0/XI0_12/d_4_ XI11_7/XI0/XI0_12/d__4_ DECAP_INV_G11
XG1970 XI11_7/XI0/XI0_12/d_3_ XI11_7/XI0/XI0_12/d__3_ DECAP_INV_G11
XG1971 XI11_7/XI0/XI0_12/d_2_ XI11_7/XI0/XI0_12/d__2_ DECAP_INV_G11
XG1972 XI11_7/XI0/XI0_12/d_1_ XI11_7/XI0/XI0_12/d__1_ DECAP_INV_G11
XG1973 XI11_7/XI0/XI0_12/d_0_ XI11_7/XI0/XI0_12/d__0_ DECAP_INV_G11
XG1974 XI11_7/XI0/XI0_11/d__15_ XI11_7/XI0/XI0_11/d_15_ DECAP_INV_G11
XG1975 XI11_7/XI0/XI0_11/d__14_ XI11_7/XI0/XI0_11/d_14_ DECAP_INV_G11
XG1976 XI11_7/XI0/XI0_11/d__13_ XI11_7/XI0/XI0_11/d_13_ DECAP_INV_G11
XG1977 XI11_7/XI0/XI0_11/d__12_ XI11_7/XI0/XI0_11/d_12_ DECAP_INV_G11
XG1978 XI11_7/XI0/XI0_11/d__11_ XI11_7/XI0/XI0_11/d_11_ DECAP_INV_G11
XG1979 XI11_7/XI0/XI0_11/d__10_ XI11_7/XI0/XI0_11/d_10_ DECAP_INV_G11
XG1980 XI11_7/XI0/XI0_11/d__9_ XI11_7/XI0/XI0_11/d_9_ DECAP_INV_G11
XG1981 XI11_7/XI0/XI0_11/d__8_ XI11_7/XI0/XI0_11/d_8_ DECAP_INV_G11
XG1982 XI11_7/XI0/XI0_11/d__7_ XI11_7/XI0/XI0_11/d_7_ DECAP_INV_G11
XG1983 XI11_7/XI0/XI0_11/d__6_ XI11_7/XI0/XI0_11/d_6_ DECAP_INV_G11
XG1984 XI11_7/XI0/XI0_11/d__5_ XI11_7/XI0/XI0_11/d_5_ DECAP_INV_G11
XG1985 XI11_7/XI0/XI0_11/d__4_ XI11_7/XI0/XI0_11/d_4_ DECAP_INV_G11
XG1986 XI11_7/XI0/XI0_11/d__3_ XI11_7/XI0/XI0_11/d_3_ DECAP_INV_G11
XG1987 XI11_7/XI0/XI0_11/d__2_ XI11_7/XI0/XI0_11/d_2_ DECAP_INV_G11
XG1988 XI11_7/XI0/XI0_11/d__1_ XI11_7/XI0/XI0_11/d_1_ DECAP_INV_G11
XG1989 XI11_7/XI0/XI0_11/d__0_ XI11_7/XI0/XI0_11/d_0_ DECAP_INV_G11
XG1990 XI11_7/XI0/XI0_11/d_15_ XI11_7/XI0/XI0_11/d__15_ DECAP_INV_G11
XG1991 XI11_7/XI0/XI0_11/d_14_ XI11_7/XI0/XI0_11/d__14_ DECAP_INV_G11
XG1992 XI11_7/XI0/XI0_11/d_13_ XI11_7/XI0/XI0_11/d__13_ DECAP_INV_G11
XG1993 XI11_7/XI0/XI0_11/d_12_ XI11_7/XI0/XI0_11/d__12_ DECAP_INV_G11
XG1994 XI11_7/XI0/XI0_11/d_11_ XI11_7/XI0/XI0_11/d__11_ DECAP_INV_G11
XG1995 XI11_7/XI0/XI0_11/d_10_ XI11_7/XI0/XI0_11/d__10_ DECAP_INV_G11
XG1996 XI11_7/XI0/XI0_11/d_9_ XI11_7/XI0/XI0_11/d__9_ DECAP_INV_G11
XG1997 XI11_7/XI0/XI0_11/d_8_ XI11_7/XI0/XI0_11/d__8_ DECAP_INV_G11
XG1998 XI11_7/XI0/XI0_11/d_7_ XI11_7/XI0/XI0_11/d__7_ DECAP_INV_G11
XG1999 XI11_7/XI0/XI0_11/d_6_ XI11_7/XI0/XI0_11/d__6_ DECAP_INV_G11
XG2000 XI11_7/XI0/XI0_11/d_5_ XI11_7/XI0/XI0_11/d__5_ DECAP_INV_G11
XG2001 XI11_7/XI0/XI0_11/d_4_ XI11_7/XI0/XI0_11/d__4_ DECAP_INV_G11
XG2002 XI11_7/XI0/XI0_11/d_3_ XI11_7/XI0/XI0_11/d__3_ DECAP_INV_G11
XG2003 XI11_7/XI0/XI0_11/d_2_ XI11_7/XI0/XI0_11/d__2_ DECAP_INV_G11
XG2004 XI11_7/XI0/XI0_11/d_1_ XI11_7/XI0/XI0_11/d__1_ DECAP_INV_G11
XG2005 XI11_7/XI0/XI0_11/d_0_ XI11_7/XI0/XI0_11/d__0_ DECAP_INV_G11
XG2006 XI11_7/XI0/XI0_10/d__15_ XI11_7/XI0/XI0_10/d_15_ DECAP_INV_G11
XG2007 XI11_7/XI0/XI0_10/d__14_ XI11_7/XI0/XI0_10/d_14_ DECAP_INV_G11
XG2008 XI11_7/XI0/XI0_10/d__13_ XI11_7/XI0/XI0_10/d_13_ DECAP_INV_G11
XG2009 XI11_7/XI0/XI0_10/d__12_ XI11_7/XI0/XI0_10/d_12_ DECAP_INV_G11
XG2010 XI11_7/XI0/XI0_10/d__11_ XI11_7/XI0/XI0_10/d_11_ DECAP_INV_G11
XG2011 XI11_7/XI0/XI0_10/d__10_ XI11_7/XI0/XI0_10/d_10_ DECAP_INV_G11
XG2012 XI11_7/XI0/XI0_10/d__9_ XI11_7/XI0/XI0_10/d_9_ DECAP_INV_G11
XG2013 XI11_7/XI0/XI0_10/d__8_ XI11_7/XI0/XI0_10/d_8_ DECAP_INV_G11
XG2014 XI11_7/XI0/XI0_10/d__7_ XI11_7/XI0/XI0_10/d_7_ DECAP_INV_G11
XG2015 XI11_7/XI0/XI0_10/d__6_ XI11_7/XI0/XI0_10/d_6_ DECAP_INV_G11
XG2016 XI11_7/XI0/XI0_10/d__5_ XI11_7/XI0/XI0_10/d_5_ DECAP_INV_G11
XG2017 XI11_7/XI0/XI0_10/d__4_ XI11_7/XI0/XI0_10/d_4_ DECAP_INV_G11
XG2018 XI11_7/XI0/XI0_10/d__3_ XI11_7/XI0/XI0_10/d_3_ DECAP_INV_G11
XG2019 XI11_7/XI0/XI0_10/d__2_ XI11_7/XI0/XI0_10/d_2_ DECAP_INV_G11
XG2020 XI11_7/XI0/XI0_10/d__1_ XI11_7/XI0/XI0_10/d_1_ DECAP_INV_G11
XG2021 XI11_7/XI0/XI0_10/d__0_ XI11_7/XI0/XI0_10/d_0_ DECAP_INV_G11
XG2022 XI11_7/XI0/XI0_10/d_15_ XI11_7/XI0/XI0_10/d__15_ DECAP_INV_G11
XG2023 XI11_7/XI0/XI0_10/d_14_ XI11_7/XI0/XI0_10/d__14_ DECAP_INV_G11
XG2024 XI11_7/XI0/XI0_10/d_13_ XI11_7/XI0/XI0_10/d__13_ DECAP_INV_G11
XG2025 XI11_7/XI0/XI0_10/d_12_ XI11_7/XI0/XI0_10/d__12_ DECAP_INV_G11
XG2026 XI11_7/XI0/XI0_10/d_11_ XI11_7/XI0/XI0_10/d__11_ DECAP_INV_G11
XG2027 XI11_7/XI0/XI0_10/d_10_ XI11_7/XI0/XI0_10/d__10_ DECAP_INV_G11
XG2028 XI11_7/XI0/XI0_10/d_9_ XI11_7/XI0/XI0_10/d__9_ DECAP_INV_G11
XG2029 XI11_7/XI0/XI0_10/d_8_ XI11_7/XI0/XI0_10/d__8_ DECAP_INV_G11
XG2030 XI11_7/XI0/XI0_10/d_7_ XI11_7/XI0/XI0_10/d__7_ DECAP_INV_G11
XG2031 XI11_7/XI0/XI0_10/d_6_ XI11_7/XI0/XI0_10/d__6_ DECAP_INV_G11
XG2032 XI11_7/XI0/XI0_10/d_5_ XI11_7/XI0/XI0_10/d__5_ DECAP_INV_G11
XG2033 XI11_7/XI0/XI0_10/d_4_ XI11_7/XI0/XI0_10/d__4_ DECAP_INV_G11
XG2034 XI11_7/XI0/XI0_10/d_3_ XI11_7/XI0/XI0_10/d__3_ DECAP_INV_G11
XG2035 XI11_7/XI0/XI0_10/d_2_ XI11_7/XI0/XI0_10/d__2_ DECAP_INV_G11
XG2036 XI11_7/XI0/XI0_10/d_1_ XI11_7/XI0/XI0_10/d__1_ DECAP_INV_G11
XG2037 XI11_7/XI0/XI0_10/d_0_ XI11_7/XI0/XI0_10/d__0_ DECAP_INV_G11
XG2038 XI11_7/XI0/XI0_9/d__15_ XI11_7/XI0/XI0_9/d_15_ DECAP_INV_G11
XG2039 XI11_7/XI0/XI0_9/d__14_ XI11_7/XI0/XI0_9/d_14_ DECAP_INV_G11
XG2040 XI11_7/XI0/XI0_9/d__13_ XI11_7/XI0/XI0_9/d_13_ DECAP_INV_G11
XG2041 XI11_7/XI0/XI0_9/d__12_ XI11_7/XI0/XI0_9/d_12_ DECAP_INV_G11
XG2042 XI11_7/XI0/XI0_9/d__11_ XI11_7/XI0/XI0_9/d_11_ DECAP_INV_G11
XG2043 XI11_7/XI0/XI0_9/d__10_ XI11_7/XI0/XI0_9/d_10_ DECAP_INV_G11
XG2044 XI11_7/XI0/XI0_9/d__9_ XI11_7/XI0/XI0_9/d_9_ DECAP_INV_G11
XG2045 XI11_7/XI0/XI0_9/d__8_ XI11_7/XI0/XI0_9/d_8_ DECAP_INV_G11
XG2046 XI11_7/XI0/XI0_9/d__7_ XI11_7/XI0/XI0_9/d_7_ DECAP_INV_G11
XG2047 XI11_7/XI0/XI0_9/d__6_ XI11_7/XI0/XI0_9/d_6_ DECAP_INV_G11
XG2048 XI11_7/XI0/XI0_9/d__5_ XI11_7/XI0/XI0_9/d_5_ DECAP_INV_G11
XG2049 XI11_7/XI0/XI0_9/d__4_ XI11_7/XI0/XI0_9/d_4_ DECAP_INV_G11
XG2050 XI11_7/XI0/XI0_9/d__3_ XI11_7/XI0/XI0_9/d_3_ DECAP_INV_G11
XG2051 XI11_7/XI0/XI0_9/d__2_ XI11_7/XI0/XI0_9/d_2_ DECAP_INV_G11
XG2052 XI11_7/XI0/XI0_9/d__1_ XI11_7/XI0/XI0_9/d_1_ DECAP_INV_G11
XG2053 XI11_7/XI0/XI0_9/d__0_ XI11_7/XI0/XI0_9/d_0_ DECAP_INV_G11
XG2054 XI11_7/XI0/XI0_9/d_15_ XI11_7/XI0/XI0_9/d__15_ DECAP_INV_G11
XG2055 XI11_7/XI0/XI0_9/d_14_ XI11_7/XI0/XI0_9/d__14_ DECAP_INV_G11
XG2056 XI11_7/XI0/XI0_9/d_13_ XI11_7/XI0/XI0_9/d__13_ DECAP_INV_G11
XG2057 XI11_7/XI0/XI0_9/d_12_ XI11_7/XI0/XI0_9/d__12_ DECAP_INV_G11
XG2058 XI11_7/XI0/XI0_9/d_11_ XI11_7/XI0/XI0_9/d__11_ DECAP_INV_G11
XG2059 XI11_7/XI0/XI0_9/d_10_ XI11_7/XI0/XI0_9/d__10_ DECAP_INV_G11
XG2060 XI11_7/XI0/XI0_9/d_9_ XI11_7/XI0/XI0_9/d__9_ DECAP_INV_G11
XG2061 XI11_7/XI0/XI0_9/d_8_ XI11_7/XI0/XI0_9/d__8_ DECAP_INV_G11
XG2062 XI11_7/XI0/XI0_9/d_7_ XI11_7/XI0/XI0_9/d__7_ DECAP_INV_G11
XG2063 XI11_7/XI0/XI0_9/d_6_ XI11_7/XI0/XI0_9/d__6_ DECAP_INV_G11
XG2064 XI11_7/XI0/XI0_9/d_5_ XI11_7/XI0/XI0_9/d__5_ DECAP_INV_G11
XG2065 XI11_7/XI0/XI0_9/d_4_ XI11_7/XI0/XI0_9/d__4_ DECAP_INV_G11
XG2066 XI11_7/XI0/XI0_9/d_3_ XI11_7/XI0/XI0_9/d__3_ DECAP_INV_G11
XG2067 XI11_7/XI0/XI0_9/d_2_ XI11_7/XI0/XI0_9/d__2_ DECAP_INV_G11
XG2068 XI11_7/XI0/XI0_9/d_1_ XI11_7/XI0/XI0_9/d__1_ DECAP_INV_G11
XG2069 XI11_7/XI0/XI0_9/d_0_ XI11_7/XI0/XI0_9/d__0_ DECAP_INV_G11
XG2070 XI11_7/XI0/XI0_8/d__15_ XI11_7/XI0/XI0_8/d_15_ DECAP_INV_G11
XG2071 XI11_7/XI0/XI0_8/d__14_ XI11_7/XI0/XI0_8/d_14_ DECAP_INV_G11
XG2072 XI11_7/XI0/XI0_8/d__13_ XI11_7/XI0/XI0_8/d_13_ DECAP_INV_G11
XG2073 XI11_7/XI0/XI0_8/d__12_ XI11_7/XI0/XI0_8/d_12_ DECAP_INV_G11
XG2074 XI11_7/XI0/XI0_8/d__11_ XI11_7/XI0/XI0_8/d_11_ DECAP_INV_G11
XG2075 XI11_7/XI0/XI0_8/d__10_ XI11_7/XI0/XI0_8/d_10_ DECAP_INV_G11
XG2076 XI11_7/XI0/XI0_8/d__9_ XI11_7/XI0/XI0_8/d_9_ DECAP_INV_G11
XG2077 XI11_7/XI0/XI0_8/d__8_ XI11_7/XI0/XI0_8/d_8_ DECAP_INV_G11
XG2078 XI11_7/XI0/XI0_8/d__7_ XI11_7/XI0/XI0_8/d_7_ DECAP_INV_G11
XG2079 XI11_7/XI0/XI0_8/d__6_ XI11_7/XI0/XI0_8/d_6_ DECAP_INV_G11
XG2080 XI11_7/XI0/XI0_8/d__5_ XI11_7/XI0/XI0_8/d_5_ DECAP_INV_G11
XG2081 XI11_7/XI0/XI0_8/d__4_ XI11_7/XI0/XI0_8/d_4_ DECAP_INV_G11
XG2082 XI11_7/XI0/XI0_8/d__3_ XI11_7/XI0/XI0_8/d_3_ DECAP_INV_G11
XG2083 XI11_7/XI0/XI0_8/d__2_ XI11_7/XI0/XI0_8/d_2_ DECAP_INV_G11
XG2084 XI11_7/XI0/XI0_8/d__1_ XI11_7/XI0/XI0_8/d_1_ DECAP_INV_G11
XG2085 XI11_7/XI0/XI0_8/d__0_ XI11_7/XI0/XI0_8/d_0_ DECAP_INV_G11
XG2086 XI11_7/XI0/XI0_8/d_15_ XI11_7/XI0/XI0_8/d__15_ DECAP_INV_G11
XG2087 XI11_7/XI0/XI0_8/d_14_ XI11_7/XI0/XI0_8/d__14_ DECAP_INV_G11
XG2088 XI11_7/XI0/XI0_8/d_13_ XI11_7/XI0/XI0_8/d__13_ DECAP_INV_G11
XG2089 XI11_7/XI0/XI0_8/d_12_ XI11_7/XI0/XI0_8/d__12_ DECAP_INV_G11
XG2090 XI11_7/XI0/XI0_8/d_11_ XI11_7/XI0/XI0_8/d__11_ DECAP_INV_G11
XG2091 XI11_7/XI0/XI0_8/d_10_ XI11_7/XI0/XI0_8/d__10_ DECAP_INV_G11
XG2092 XI11_7/XI0/XI0_8/d_9_ XI11_7/XI0/XI0_8/d__9_ DECAP_INV_G11
XG2093 XI11_7/XI0/XI0_8/d_8_ XI11_7/XI0/XI0_8/d__8_ DECAP_INV_G11
XG2094 XI11_7/XI0/XI0_8/d_7_ XI11_7/XI0/XI0_8/d__7_ DECAP_INV_G11
XG2095 XI11_7/XI0/XI0_8/d_6_ XI11_7/XI0/XI0_8/d__6_ DECAP_INV_G11
XG2096 XI11_7/XI0/XI0_8/d_5_ XI11_7/XI0/XI0_8/d__5_ DECAP_INV_G11
XG2097 XI11_7/XI0/XI0_8/d_4_ XI11_7/XI0/XI0_8/d__4_ DECAP_INV_G11
XG2098 XI11_7/XI0/XI0_8/d_3_ XI11_7/XI0/XI0_8/d__3_ DECAP_INV_G11
XG2099 XI11_7/XI0/XI0_8/d_2_ XI11_7/XI0/XI0_8/d__2_ DECAP_INV_G11
XG2100 XI11_7/XI0/XI0_8/d_1_ XI11_7/XI0/XI0_8/d__1_ DECAP_INV_G11
XG2101 XI11_7/XI0/XI0_8/d_0_ XI11_7/XI0/XI0_8/d__0_ DECAP_INV_G11
XG2102 XI11_7/XI0/XI0_7/d__15_ XI11_7/XI0/XI0_7/d_15_ DECAP_INV_G11
XG2103 XI11_7/XI0/XI0_7/d__14_ XI11_7/XI0/XI0_7/d_14_ DECAP_INV_G11
XG2104 XI11_7/XI0/XI0_7/d__13_ XI11_7/XI0/XI0_7/d_13_ DECAP_INV_G11
XG2105 XI11_7/XI0/XI0_7/d__12_ XI11_7/XI0/XI0_7/d_12_ DECAP_INV_G11
XG2106 XI11_7/XI0/XI0_7/d__11_ XI11_7/XI0/XI0_7/d_11_ DECAP_INV_G11
XG2107 XI11_7/XI0/XI0_7/d__10_ XI11_7/XI0/XI0_7/d_10_ DECAP_INV_G11
XG2108 XI11_7/XI0/XI0_7/d__9_ XI11_7/XI0/XI0_7/d_9_ DECAP_INV_G11
XG2109 XI11_7/XI0/XI0_7/d__8_ XI11_7/XI0/XI0_7/d_8_ DECAP_INV_G11
XG2110 XI11_7/XI0/XI0_7/d__7_ XI11_7/XI0/XI0_7/d_7_ DECAP_INV_G11
XG2111 XI11_7/XI0/XI0_7/d__6_ XI11_7/XI0/XI0_7/d_6_ DECAP_INV_G11
XG2112 XI11_7/XI0/XI0_7/d__5_ XI11_7/XI0/XI0_7/d_5_ DECAP_INV_G11
XG2113 XI11_7/XI0/XI0_7/d__4_ XI11_7/XI0/XI0_7/d_4_ DECAP_INV_G11
XG2114 XI11_7/XI0/XI0_7/d__3_ XI11_7/XI0/XI0_7/d_3_ DECAP_INV_G11
XG2115 XI11_7/XI0/XI0_7/d__2_ XI11_7/XI0/XI0_7/d_2_ DECAP_INV_G11
XG2116 XI11_7/XI0/XI0_7/d__1_ XI11_7/XI0/XI0_7/d_1_ DECAP_INV_G11
XG2117 XI11_7/XI0/XI0_7/d__0_ XI11_7/XI0/XI0_7/d_0_ DECAP_INV_G11
XG2118 XI11_7/XI0/XI0_7/d_15_ XI11_7/XI0/XI0_7/d__15_ DECAP_INV_G11
XG2119 XI11_7/XI0/XI0_7/d_14_ XI11_7/XI0/XI0_7/d__14_ DECAP_INV_G11
XG2120 XI11_7/XI0/XI0_7/d_13_ XI11_7/XI0/XI0_7/d__13_ DECAP_INV_G11
XG2121 XI11_7/XI0/XI0_7/d_12_ XI11_7/XI0/XI0_7/d__12_ DECAP_INV_G11
XG2122 XI11_7/XI0/XI0_7/d_11_ XI11_7/XI0/XI0_7/d__11_ DECAP_INV_G11
XG2123 XI11_7/XI0/XI0_7/d_10_ XI11_7/XI0/XI0_7/d__10_ DECAP_INV_G11
XG2124 XI11_7/XI0/XI0_7/d_9_ XI11_7/XI0/XI0_7/d__9_ DECAP_INV_G11
XG2125 XI11_7/XI0/XI0_7/d_8_ XI11_7/XI0/XI0_7/d__8_ DECAP_INV_G11
XG2126 XI11_7/XI0/XI0_7/d_7_ XI11_7/XI0/XI0_7/d__7_ DECAP_INV_G11
XG2127 XI11_7/XI0/XI0_7/d_6_ XI11_7/XI0/XI0_7/d__6_ DECAP_INV_G11
XG2128 XI11_7/XI0/XI0_7/d_5_ XI11_7/XI0/XI0_7/d__5_ DECAP_INV_G11
XG2129 XI11_7/XI0/XI0_7/d_4_ XI11_7/XI0/XI0_7/d__4_ DECAP_INV_G11
XG2130 XI11_7/XI0/XI0_7/d_3_ XI11_7/XI0/XI0_7/d__3_ DECAP_INV_G11
XG2131 XI11_7/XI0/XI0_7/d_2_ XI11_7/XI0/XI0_7/d__2_ DECAP_INV_G11
XG2132 XI11_7/XI0/XI0_7/d_1_ XI11_7/XI0/XI0_7/d__1_ DECAP_INV_G11
XG2133 XI11_7/XI0/XI0_7/d_0_ XI11_7/XI0/XI0_7/d__0_ DECAP_INV_G11
XG2134 XI11_7/XI0/XI0_6/d__15_ XI11_7/XI0/XI0_6/d_15_ DECAP_INV_G11
XG2135 XI11_7/XI0/XI0_6/d__14_ XI11_7/XI0/XI0_6/d_14_ DECAP_INV_G11
XG2136 XI11_7/XI0/XI0_6/d__13_ XI11_7/XI0/XI0_6/d_13_ DECAP_INV_G11
XG2137 XI11_7/XI0/XI0_6/d__12_ XI11_7/XI0/XI0_6/d_12_ DECAP_INV_G11
XG2138 XI11_7/XI0/XI0_6/d__11_ XI11_7/XI0/XI0_6/d_11_ DECAP_INV_G11
XG2139 XI11_7/XI0/XI0_6/d__10_ XI11_7/XI0/XI0_6/d_10_ DECAP_INV_G11
XG2140 XI11_7/XI0/XI0_6/d__9_ XI11_7/XI0/XI0_6/d_9_ DECAP_INV_G11
XG2141 XI11_7/XI0/XI0_6/d__8_ XI11_7/XI0/XI0_6/d_8_ DECAP_INV_G11
XG2142 XI11_7/XI0/XI0_6/d__7_ XI11_7/XI0/XI0_6/d_7_ DECAP_INV_G11
XG2143 XI11_7/XI0/XI0_6/d__6_ XI11_7/XI0/XI0_6/d_6_ DECAP_INV_G11
XG2144 XI11_7/XI0/XI0_6/d__5_ XI11_7/XI0/XI0_6/d_5_ DECAP_INV_G11
XG2145 XI11_7/XI0/XI0_6/d__4_ XI11_7/XI0/XI0_6/d_4_ DECAP_INV_G11
XG2146 XI11_7/XI0/XI0_6/d__3_ XI11_7/XI0/XI0_6/d_3_ DECAP_INV_G11
XG2147 XI11_7/XI0/XI0_6/d__2_ XI11_7/XI0/XI0_6/d_2_ DECAP_INV_G11
XG2148 XI11_7/XI0/XI0_6/d__1_ XI11_7/XI0/XI0_6/d_1_ DECAP_INV_G11
XG2149 XI11_7/XI0/XI0_6/d__0_ XI11_7/XI0/XI0_6/d_0_ DECAP_INV_G11
XG2150 XI11_7/XI0/XI0_6/d_15_ XI11_7/XI0/XI0_6/d__15_ DECAP_INV_G11
XG2151 XI11_7/XI0/XI0_6/d_14_ XI11_7/XI0/XI0_6/d__14_ DECAP_INV_G11
XG2152 XI11_7/XI0/XI0_6/d_13_ XI11_7/XI0/XI0_6/d__13_ DECAP_INV_G11
XG2153 XI11_7/XI0/XI0_6/d_12_ XI11_7/XI0/XI0_6/d__12_ DECAP_INV_G11
XG2154 XI11_7/XI0/XI0_6/d_11_ XI11_7/XI0/XI0_6/d__11_ DECAP_INV_G11
XG2155 XI11_7/XI0/XI0_6/d_10_ XI11_7/XI0/XI0_6/d__10_ DECAP_INV_G11
XG2156 XI11_7/XI0/XI0_6/d_9_ XI11_7/XI0/XI0_6/d__9_ DECAP_INV_G11
XG2157 XI11_7/XI0/XI0_6/d_8_ XI11_7/XI0/XI0_6/d__8_ DECAP_INV_G11
XG2158 XI11_7/XI0/XI0_6/d_7_ XI11_7/XI0/XI0_6/d__7_ DECAP_INV_G11
XG2159 XI11_7/XI0/XI0_6/d_6_ XI11_7/XI0/XI0_6/d__6_ DECAP_INV_G11
XG2160 XI11_7/XI0/XI0_6/d_5_ XI11_7/XI0/XI0_6/d__5_ DECAP_INV_G11
XG2161 XI11_7/XI0/XI0_6/d_4_ XI11_7/XI0/XI0_6/d__4_ DECAP_INV_G11
XG2162 XI11_7/XI0/XI0_6/d_3_ XI11_7/XI0/XI0_6/d__3_ DECAP_INV_G11
XG2163 XI11_7/XI0/XI0_6/d_2_ XI11_7/XI0/XI0_6/d__2_ DECAP_INV_G11
XG2164 XI11_7/XI0/XI0_6/d_1_ XI11_7/XI0/XI0_6/d__1_ DECAP_INV_G11
XG2165 XI11_7/XI0/XI0_6/d_0_ XI11_7/XI0/XI0_6/d__0_ DECAP_INV_G11
XG2166 XI11_7/XI0/XI0_5/d__15_ XI11_7/XI0/XI0_5/d_15_ DECAP_INV_G11
XG2167 XI11_7/XI0/XI0_5/d__14_ XI11_7/XI0/XI0_5/d_14_ DECAP_INV_G11
XG2168 XI11_7/XI0/XI0_5/d__13_ XI11_7/XI0/XI0_5/d_13_ DECAP_INV_G11
XG2169 XI11_7/XI0/XI0_5/d__12_ XI11_7/XI0/XI0_5/d_12_ DECAP_INV_G11
XG2170 XI11_7/XI0/XI0_5/d__11_ XI11_7/XI0/XI0_5/d_11_ DECAP_INV_G11
XG2171 XI11_7/XI0/XI0_5/d__10_ XI11_7/XI0/XI0_5/d_10_ DECAP_INV_G11
XG2172 XI11_7/XI0/XI0_5/d__9_ XI11_7/XI0/XI0_5/d_9_ DECAP_INV_G11
XG2173 XI11_7/XI0/XI0_5/d__8_ XI11_7/XI0/XI0_5/d_8_ DECAP_INV_G11
XG2174 XI11_7/XI0/XI0_5/d__7_ XI11_7/XI0/XI0_5/d_7_ DECAP_INV_G11
XG2175 XI11_7/XI0/XI0_5/d__6_ XI11_7/XI0/XI0_5/d_6_ DECAP_INV_G11
XG2176 XI11_7/XI0/XI0_5/d__5_ XI11_7/XI0/XI0_5/d_5_ DECAP_INV_G11
XG2177 XI11_7/XI0/XI0_5/d__4_ XI11_7/XI0/XI0_5/d_4_ DECAP_INV_G11
XG2178 XI11_7/XI0/XI0_5/d__3_ XI11_7/XI0/XI0_5/d_3_ DECAP_INV_G11
XG2179 XI11_7/XI0/XI0_5/d__2_ XI11_7/XI0/XI0_5/d_2_ DECAP_INV_G11
XG2180 XI11_7/XI0/XI0_5/d__1_ XI11_7/XI0/XI0_5/d_1_ DECAP_INV_G11
XG2181 XI11_7/XI0/XI0_5/d__0_ XI11_7/XI0/XI0_5/d_0_ DECAP_INV_G11
XG2182 XI11_7/XI0/XI0_5/d_15_ XI11_7/XI0/XI0_5/d__15_ DECAP_INV_G11
XG2183 XI11_7/XI0/XI0_5/d_14_ XI11_7/XI0/XI0_5/d__14_ DECAP_INV_G11
XG2184 XI11_7/XI0/XI0_5/d_13_ XI11_7/XI0/XI0_5/d__13_ DECAP_INV_G11
XG2185 XI11_7/XI0/XI0_5/d_12_ XI11_7/XI0/XI0_5/d__12_ DECAP_INV_G11
XG2186 XI11_7/XI0/XI0_5/d_11_ XI11_7/XI0/XI0_5/d__11_ DECAP_INV_G11
XG2187 XI11_7/XI0/XI0_5/d_10_ XI11_7/XI0/XI0_5/d__10_ DECAP_INV_G11
XG2188 XI11_7/XI0/XI0_5/d_9_ XI11_7/XI0/XI0_5/d__9_ DECAP_INV_G11
XG2189 XI11_7/XI0/XI0_5/d_8_ XI11_7/XI0/XI0_5/d__8_ DECAP_INV_G11
XG2190 XI11_7/XI0/XI0_5/d_7_ XI11_7/XI0/XI0_5/d__7_ DECAP_INV_G11
XG2191 XI11_7/XI0/XI0_5/d_6_ XI11_7/XI0/XI0_5/d__6_ DECAP_INV_G11
XG2192 XI11_7/XI0/XI0_5/d_5_ XI11_7/XI0/XI0_5/d__5_ DECAP_INV_G11
XG2193 XI11_7/XI0/XI0_5/d_4_ XI11_7/XI0/XI0_5/d__4_ DECAP_INV_G11
XG2194 XI11_7/XI0/XI0_5/d_3_ XI11_7/XI0/XI0_5/d__3_ DECAP_INV_G11
XG2195 XI11_7/XI0/XI0_5/d_2_ XI11_7/XI0/XI0_5/d__2_ DECAP_INV_G11
XG2196 XI11_7/XI0/XI0_5/d_1_ XI11_7/XI0/XI0_5/d__1_ DECAP_INV_G11
XG2197 XI11_7/XI0/XI0_5/d_0_ XI11_7/XI0/XI0_5/d__0_ DECAP_INV_G11
XG2198 XI11_7/XI0/XI0_4/d__15_ XI11_7/XI0/XI0_4/d_15_ DECAP_INV_G11
XG2199 XI11_7/XI0/XI0_4/d__14_ XI11_7/XI0/XI0_4/d_14_ DECAP_INV_G11
XG2200 XI11_7/XI0/XI0_4/d__13_ XI11_7/XI0/XI0_4/d_13_ DECAP_INV_G11
XG2201 XI11_7/XI0/XI0_4/d__12_ XI11_7/XI0/XI0_4/d_12_ DECAP_INV_G11
XG2202 XI11_7/XI0/XI0_4/d__11_ XI11_7/XI0/XI0_4/d_11_ DECAP_INV_G11
XG2203 XI11_7/XI0/XI0_4/d__10_ XI11_7/XI0/XI0_4/d_10_ DECAP_INV_G11
XG2204 XI11_7/XI0/XI0_4/d__9_ XI11_7/XI0/XI0_4/d_9_ DECAP_INV_G11
XG2205 XI11_7/XI0/XI0_4/d__8_ XI11_7/XI0/XI0_4/d_8_ DECAP_INV_G11
XG2206 XI11_7/XI0/XI0_4/d__7_ XI11_7/XI0/XI0_4/d_7_ DECAP_INV_G11
XG2207 XI11_7/XI0/XI0_4/d__6_ XI11_7/XI0/XI0_4/d_6_ DECAP_INV_G11
XG2208 XI11_7/XI0/XI0_4/d__5_ XI11_7/XI0/XI0_4/d_5_ DECAP_INV_G11
XG2209 XI11_7/XI0/XI0_4/d__4_ XI11_7/XI0/XI0_4/d_4_ DECAP_INV_G11
XG2210 XI11_7/XI0/XI0_4/d__3_ XI11_7/XI0/XI0_4/d_3_ DECAP_INV_G11
XG2211 XI11_7/XI0/XI0_4/d__2_ XI11_7/XI0/XI0_4/d_2_ DECAP_INV_G11
XG2212 XI11_7/XI0/XI0_4/d__1_ XI11_7/XI0/XI0_4/d_1_ DECAP_INV_G11
XG2213 XI11_7/XI0/XI0_4/d__0_ XI11_7/XI0/XI0_4/d_0_ DECAP_INV_G11
XG2214 XI11_7/XI0/XI0_4/d_15_ XI11_7/XI0/XI0_4/d__15_ DECAP_INV_G11
XG2215 XI11_7/XI0/XI0_4/d_14_ XI11_7/XI0/XI0_4/d__14_ DECAP_INV_G11
XG2216 XI11_7/XI0/XI0_4/d_13_ XI11_7/XI0/XI0_4/d__13_ DECAP_INV_G11
XG2217 XI11_7/XI0/XI0_4/d_12_ XI11_7/XI0/XI0_4/d__12_ DECAP_INV_G11
XG2218 XI11_7/XI0/XI0_4/d_11_ XI11_7/XI0/XI0_4/d__11_ DECAP_INV_G11
XG2219 XI11_7/XI0/XI0_4/d_10_ XI11_7/XI0/XI0_4/d__10_ DECAP_INV_G11
XG2220 XI11_7/XI0/XI0_4/d_9_ XI11_7/XI0/XI0_4/d__9_ DECAP_INV_G11
XG2221 XI11_7/XI0/XI0_4/d_8_ XI11_7/XI0/XI0_4/d__8_ DECAP_INV_G11
XG2222 XI11_7/XI0/XI0_4/d_7_ XI11_7/XI0/XI0_4/d__7_ DECAP_INV_G11
XG2223 XI11_7/XI0/XI0_4/d_6_ XI11_7/XI0/XI0_4/d__6_ DECAP_INV_G11
XG2224 XI11_7/XI0/XI0_4/d_5_ XI11_7/XI0/XI0_4/d__5_ DECAP_INV_G11
XG2225 XI11_7/XI0/XI0_4/d_4_ XI11_7/XI0/XI0_4/d__4_ DECAP_INV_G11
XG2226 XI11_7/XI0/XI0_4/d_3_ XI11_7/XI0/XI0_4/d__3_ DECAP_INV_G11
XG2227 XI11_7/XI0/XI0_4/d_2_ XI11_7/XI0/XI0_4/d__2_ DECAP_INV_G11
XG2228 XI11_7/XI0/XI0_4/d_1_ XI11_7/XI0/XI0_4/d__1_ DECAP_INV_G11
XG2229 XI11_7/XI0/XI0_4/d_0_ XI11_7/XI0/XI0_4/d__0_ DECAP_INV_G11
XG2230 XI11_7/XI0/XI0_3/d__15_ XI11_7/XI0/XI0_3/d_15_ DECAP_INV_G11
XG2231 XI11_7/XI0/XI0_3/d__14_ XI11_7/XI0/XI0_3/d_14_ DECAP_INV_G11
XG2232 XI11_7/XI0/XI0_3/d__13_ XI11_7/XI0/XI0_3/d_13_ DECAP_INV_G11
XG2233 XI11_7/XI0/XI0_3/d__12_ XI11_7/XI0/XI0_3/d_12_ DECAP_INV_G11
XG2234 XI11_7/XI0/XI0_3/d__11_ XI11_7/XI0/XI0_3/d_11_ DECAP_INV_G11
XG2235 XI11_7/XI0/XI0_3/d__10_ XI11_7/XI0/XI0_3/d_10_ DECAP_INV_G11
XG2236 XI11_7/XI0/XI0_3/d__9_ XI11_7/XI0/XI0_3/d_9_ DECAP_INV_G11
XG2237 XI11_7/XI0/XI0_3/d__8_ XI11_7/XI0/XI0_3/d_8_ DECAP_INV_G11
XG2238 XI11_7/XI0/XI0_3/d__7_ XI11_7/XI0/XI0_3/d_7_ DECAP_INV_G11
XG2239 XI11_7/XI0/XI0_3/d__6_ XI11_7/XI0/XI0_3/d_6_ DECAP_INV_G11
XG2240 XI11_7/XI0/XI0_3/d__5_ XI11_7/XI0/XI0_3/d_5_ DECAP_INV_G11
XG2241 XI11_7/XI0/XI0_3/d__4_ XI11_7/XI0/XI0_3/d_4_ DECAP_INV_G11
XG2242 XI11_7/XI0/XI0_3/d__3_ XI11_7/XI0/XI0_3/d_3_ DECAP_INV_G11
XG2243 XI11_7/XI0/XI0_3/d__2_ XI11_7/XI0/XI0_3/d_2_ DECAP_INV_G11
XG2244 XI11_7/XI0/XI0_3/d__1_ XI11_7/XI0/XI0_3/d_1_ DECAP_INV_G11
XG2245 XI11_7/XI0/XI0_3/d__0_ XI11_7/XI0/XI0_3/d_0_ DECAP_INV_G11
XG2246 XI11_7/XI0/XI0_3/d_15_ XI11_7/XI0/XI0_3/d__15_ DECAP_INV_G11
XG2247 XI11_7/XI0/XI0_3/d_14_ XI11_7/XI0/XI0_3/d__14_ DECAP_INV_G11
XG2248 XI11_7/XI0/XI0_3/d_13_ XI11_7/XI0/XI0_3/d__13_ DECAP_INV_G11
XG2249 XI11_7/XI0/XI0_3/d_12_ XI11_7/XI0/XI0_3/d__12_ DECAP_INV_G11
XG2250 XI11_7/XI0/XI0_3/d_11_ XI11_7/XI0/XI0_3/d__11_ DECAP_INV_G11
XG2251 XI11_7/XI0/XI0_3/d_10_ XI11_7/XI0/XI0_3/d__10_ DECAP_INV_G11
XG2252 XI11_7/XI0/XI0_3/d_9_ XI11_7/XI0/XI0_3/d__9_ DECAP_INV_G11
XG2253 XI11_7/XI0/XI0_3/d_8_ XI11_7/XI0/XI0_3/d__8_ DECAP_INV_G11
XG2254 XI11_7/XI0/XI0_3/d_7_ XI11_7/XI0/XI0_3/d__7_ DECAP_INV_G11
XG2255 XI11_7/XI0/XI0_3/d_6_ XI11_7/XI0/XI0_3/d__6_ DECAP_INV_G11
XG2256 XI11_7/XI0/XI0_3/d_5_ XI11_7/XI0/XI0_3/d__5_ DECAP_INV_G11
XG2257 XI11_7/XI0/XI0_3/d_4_ XI11_7/XI0/XI0_3/d__4_ DECAP_INV_G11
XG2258 XI11_7/XI0/XI0_3/d_3_ XI11_7/XI0/XI0_3/d__3_ DECAP_INV_G11
XG2259 XI11_7/XI0/XI0_3/d_2_ XI11_7/XI0/XI0_3/d__2_ DECAP_INV_G11
XG2260 XI11_7/XI0/XI0_3/d_1_ XI11_7/XI0/XI0_3/d__1_ DECAP_INV_G11
XG2261 XI11_7/XI0/XI0_3/d_0_ XI11_7/XI0/XI0_3/d__0_ DECAP_INV_G11
XG2262 XI11_7/XI0/XI0_2/d__15_ XI11_7/XI0/XI0_2/d_15_ DECAP_INV_G11
XG2263 XI11_7/XI0/XI0_2/d__14_ XI11_7/XI0/XI0_2/d_14_ DECAP_INV_G11
XG2264 XI11_7/XI0/XI0_2/d__13_ XI11_7/XI0/XI0_2/d_13_ DECAP_INV_G11
XG2265 XI11_7/XI0/XI0_2/d__12_ XI11_7/XI0/XI0_2/d_12_ DECAP_INV_G11
XG2266 XI11_7/XI0/XI0_2/d__11_ XI11_7/XI0/XI0_2/d_11_ DECAP_INV_G11
XG2267 XI11_7/XI0/XI0_2/d__10_ XI11_7/XI0/XI0_2/d_10_ DECAP_INV_G11
XG2268 XI11_7/XI0/XI0_2/d__9_ XI11_7/XI0/XI0_2/d_9_ DECAP_INV_G11
XG2269 XI11_7/XI0/XI0_2/d__8_ XI11_7/XI0/XI0_2/d_8_ DECAP_INV_G11
XG2270 XI11_7/XI0/XI0_2/d__7_ XI11_7/XI0/XI0_2/d_7_ DECAP_INV_G11
XG2271 XI11_7/XI0/XI0_2/d__6_ XI11_7/XI0/XI0_2/d_6_ DECAP_INV_G11
XG2272 XI11_7/XI0/XI0_2/d__5_ XI11_7/XI0/XI0_2/d_5_ DECAP_INV_G11
XG2273 XI11_7/XI0/XI0_2/d__4_ XI11_7/XI0/XI0_2/d_4_ DECAP_INV_G11
XG2274 XI11_7/XI0/XI0_2/d__3_ XI11_7/XI0/XI0_2/d_3_ DECAP_INV_G11
XG2275 XI11_7/XI0/XI0_2/d__2_ XI11_7/XI0/XI0_2/d_2_ DECAP_INV_G11
XG2276 XI11_7/XI0/XI0_2/d__1_ XI11_7/XI0/XI0_2/d_1_ DECAP_INV_G11
XG2277 XI11_7/XI0/XI0_2/d__0_ XI11_7/XI0/XI0_2/d_0_ DECAP_INV_G11
XG2278 XI11_7/XI0/XI0_2/d_15_ XI11_7/XI0/XI0_2/d__15_ DECAP_INV_G11
XG2279 XI11_7/XI0/XI0_2/d_14_ XI11_7/XI0/XI0_2/d__14_ DECAP_INV_G11
XG2280 XI11_7/XI0/XI0_2/d_13_ XI11_7/XI0/XI0_2/d__13_ DECAP_INV_G11
XG2281 XI11_7/XI0/XI0_2/d_12_ XI11_7/XI0/XI0_2/d__12_ DECAP_INV_G11
XG2282 XI11_7/XI0/XI0_2/d_11_ XI11_7/XI0/XI0_2/d__11_ DECAP_INV_G11
XG2283 XI11_7/XI0/XI0_2/d_10_ XI11_7/XI0/XI0_2/d__10_ DECAP_INV_G11
XG2284 XI11_7/XI0/XI0_2/d_9_ XI11_7/XI0/XI0_2/d__9_ DECAP_INV_G11
XG2285 XI11_7/XI0/XI0_2/d_8_ XI11_7/XI0/XI0_2/d__8_ DECAP_INV_G11
XG2286 XI11_7/XI0/XI0_2/d_7_ XI11_7/XI0/XI0_2/d__7_ DECAP_INV_G11
XG2287 XI11_7/XI0/XI0_2/d_6_ XI11_7/XI0/XI0_2/d__6_ DECAP_INV_G11
XG2288 XI11_7/XI0/XI0_2/d_5_ XI11_7/XI0/XI0_2/d__5_ DECAP_INV_G11
XG2289 XI11_7/XI0/XI0_2/d_4_ XI11_7/XI0/XI0_2/d__4_ DECAP_INV_G11
XG2290 XI11_7/XI0/XI0_2/d_3_ XI11_7/XI0/XI0_2/d__3_ DECAP_INV_G11
XG2291 XI11_7/XI0/XI0_2/d_2_ XI11_7/XI0/XI0_2/d__2_ DECAP_INV_G11
XG2292 XI11_7/XI0/XI0_2/d_1_ XI11_7/XI0/XI0_2/d__1_ DECAP_INV_G11
XG2293 XI11_7/XI0/XI0_2/d_0_ XI11_7/XI0/XI0_2/d__0_ DECAP_INV_G11
XG2294 XI11_7/XI0/XI0_1/d__15_ XI11_7/XI0/XI0_1/d_15_ DECAP_INV_G11
XG2295 XI11_7/XI0/XI0_1/d__14_ XI11_7/XI0/XI0_1/d_14_ DECAP_INV_G11
XG2296 XI11_7/XI0/XI0_1/d__13_ XI11_7/XI0/XI0_1/d_13_ DECAP_INV_G11
XG2297 XI11_7/XI0/XI0_1/d__12_ XI11_7/XI0/XI0_1/d_12_ DECAP_INV_G11
XG2298 XI11_7/XI0/XI0_1/d__11_ XI11_7/XI0/XI0_1/d_11_ DECAP_INV_G11
XG2299 XI11_7/XI0/XI0_1/d__10_ XI11_7/XI0/XI0_1/d_10_ DECAP_INV_G11
XG2300 XI11_7/XI0/XI0_1/d__9_ XI11_7/XI0/XI0_1/d_9_ DECAP_INV_G11
XG2301 XI11_7/XI0/XI0_1/d__8_ XI11_7/XI0/XI0_1/d_8_ DECAP_INV_G11
XG2302 XI11_7/XI0/XI0_1/d__7_ XI11_7/XI0/XI0_1/d_7_ DECAP_INV_G11
XG2303 XI11_7/XI0/XI0_1/d__6_ XI11_7/XI0/XI0_1/d_6_ DECAP_INV_G11
XG2304 XI11_7/XI0/XI0_1/d__5_ XI11_7/XI0/XI0_1/d_5_ DECAP_INV_G11
XG2305 XI11_7/XI0/XI0_1/d__4_ XI11_7/XI0/XI0_1/d_4_ DECAP_INV_G11
XG2306 XI11_7/XI0/XI0_1/d__3_ XI11_7/XI0/XI0_1/d_3_ DECAP_INV_G11
XG2307 XI11_7/XI0/XI0_1/d__2_ XI11_7/XI0/XI0_1/d_2_ DECAP_INV_G11
XG2308 XI11_7/XI0/XI0_1/d__1_ XI11_7/XI0/XI0_1/d_1_ DECAP_INV_G11
XG2309 XI11_7/XI0/XI0_1/d__0_ XI11_7/XI0/XI0_1/d_0_ DECAP_INV_G11
XG2310 XI11_7/XI0/XI0_1/d_15_ XI11_7/XI0/XI0_1/d__15_ DECAP_INV_G11
XG2311 XI11_7/XI0/XI0_1/d_14_ XI11_7/XI0/XI0_1/d__14_ DECAP_INV_G11
XG2312 XI11_7/XI0/XI0_1/d_13_ XI11_7/XI0/XI0_1/d__13_ DECAP_INV_G11
XG2313 XI11_7/XI0/XI0_1/d_12_ XI11_7/XI0/XI0_1/d__12_ DECAP_INV_G11
XG2314 XI11_7/XI0/XI0_1/d_11_ XI11_7/XI0/XI0_1/d__11_ DECAP_INV_G11
XG2315 XI11_7/XI0/XI0_1/d_10_ XI11_7/XI0/XI0_1/d__10_ DECAP_INV_G11
XG2316 XI11_7/XI0/XI0_1/d_9_ XI11_7/XI0/XI0_1/d__9_ DECAP_INV_G11
XG2317 XI11_7/XI0/XI0_1/d_8_ XI11_7/XI0/XI0_1/d__8_ DECAP_INV_G11
XG2318 XI11_7/XI0/XI0_1/d_7_ XI11_7/XI0/XI0_1/d__7_ DECAP_INV_G11
XG2319 XI11_7/XI0/XI0_1/d_6_ XI11_7/XI0/XI0_1/d__6_ DECAP_INV_G11
XG2320 XI11_7/XI0/XI0_1/d_5_ XI11_7/XI0/XI0_1/d__5_ DECAP_INV_G11
XG2321 XI11_7/XI0/XI0_1/d_4_ XI11_7/XI0/XI0_1/d__4_ DECAP_INV_G11
XG2322 XI11_7/XI0/XI0_1/d_3_ XI11_7/XI0/XI0_1/d__3_ DECAP_INV_G11
XG2323 XI11_7/XI0/XI0_1/d_2_ XI11_7/XI0/XI0_1/d__2_ DECAP_INV_G11
XG2324 XI11_7/XI0/XI0_1/d_1_ XI11_7/XI0/XI0_1/d__1_ DECAP_INV_G11
XG2325 XI11_7/XI0/XI0_1/d_0_ XI11_7/XI0/XI0_1/d__0_ DECAP_INV_G11
XG2326 XI11_7/XI0/XI0_0/d__15_ XI11_7/XI0/XI0_0/d_15_ DECAP_INV_G11
XG2327 XI11_7/XI0/XI0_0/d__14_ XI11_7/XI0/XI0_0/d_14_ DECAP_INV_G11
XG2328 XI11_7/XI0/XI0_0/d__13_ XI11_7/XI0/XI0_0/d_13_ DECAP_INV_G11
XG2329 XI11_7/XI0/XI0_0/d__12_ XI11_7/XI0/XI0_0/d_12_ DECAP_INV_G11
XG2330 XI11_7/XI0/XI0_0/d__11_ XI11_7/XI0/XI0_0/d_11_ DECAP_INV_G11
XG2331 XI11_7/XI0/XI0_0/d__10_ XI11_7/XI0/XI0_0/d_10_ DECAP_INV_G11
XG2332 XI11_7/XI0/XI0_0/d__9_ XI11_7/XI0/XI0_0/d_9_ DECAP_INV_G11
XG2333 XI11_7/XI0/XI0_0/d__8_ XI11_7/XI0/XI0_0/d_8_ DECAP_INV_G11
XG2334 XI11_7/XI0/XI0_0/d__7_ XI11_7/XI0/XI0_0/d_7_ DECAP_INV_G11
XG2335 XI11_7/XI0/XI0_0/d__6_ XI11_7/XI0/XI0_0/d_6_ DECAP_INV_G11
XG2336 XI11_7/XI0/XI0_0/d__5_ XI11_7/XI0/XI0_0/d_5_ DECAP_INV_G11
XG2337 XI11_7/XI0/XI0_0/d__4_ XI11_7/XI0/XI0_0/d_4_ DECAP_INV_G11
XG2338 XI11_7/XI0/XI0_0/d__3_ XI11_7/XI0/XI0_0/d_3_ DECAP_INV_G11
XG2339 XI11_7/XI0/XI0_0/d__2_ XI11_7/XI0/XI0_0/d_2_ DECAP_INV_G11
XG2340 XI11_7/XI0/XI0_0/d__1_ XI11_7/XI0/XI0_0/d_1_ DECAP_INV_G11
XG2341 XI11_7/XI0/XI0_0/d__0_ XI11_7/XI0/XI0_0/d_0_ DECAP_INV_G11
XG2342 XI11_7/XI0/XI0_0/d_15_ XI11_7/XI0/XI0_0/d__15_ DECAP_INV_G11
XG2343 XI11_7/XI0/XI0_0/d_14_ XI11_7/XI0/XI0_0/d__14_ DECAP_INV_G11
XG2344 XI11_7/XI0/XI0_0/d_13_ XI11_7/XI0/XI0_0/d__13_ DECAP_INV_G11
XG2345 XI11_7/XI0/XI0_0/d_12_ XI11_7/XI0/XI0_0/d__12_ DECAP_INV_G11
XG2346 XI11_7/XI0/XI0_0/d_11_ XI11_7/XI0/XI0_0/d__11_ DECAP_INV_G11
XG2347 XI11_7/XI0/XI0_0/d_10_ XI11_7/XI0/XI0_0/d__10_ DECAP_INV_G11
XG2348 XI11_7/XI0/XI0_0/d_9_ XI11_7/XI0/XI0_0/d__9_ DECAP_INV_G11
XG2349 XI11_7/XI0/XI0_0/d_8_ XI11_7/XI0/XI0_0/d__8_ DECAP_INV_G11
XG2350 XI11_7/XI0/XI0_0/d_7_ XI11_7/XI0/XI0_0/d__7_ DECAP_INV_G11
XG2351 XI11_7/XI0/XI0_0/d_6_ XI11_7/XI0/XI0_0/d__6_ DECAP_INV_G11
XG2352 XI11_7/XI0/XI0_0/d_5_ XI11_7/XI0/XI0_0/d__5_ DECAP_INV_G11
XG2353 XI11_7/XI0/XI0_0/d_4_ XI11_7/XI0/XI0_0/d__4_ DECAP_INV_G11
XG2354 XI11_7/XI0/XI0_0/d_3_ XI11_7/XI0/XI0_0/d__3_ DECAP_INV_G11
XG2355 XI11_7/XI0/XI0_0/d_2_ XI11_7/XI0/XI0_0/d__2_ DECAP_INV_G11
XG2356 XI11_7/XI0/XI0_0/d_1_ XI11_7/XI0/XI0_0/d__1_ DECAP_INV_G11
XG2357 XI11_7/XI0/XI0_0/d_0_ XI11_7/XI0/XI0_0/d__0_ DECAP_INV_G11
XG2358 XI11_6/XI3/net17 XI11_6/XI3/net5 DECAP_INV_G7
XG2359 XI11_6/XI3/net5 XI11_6/preck DECAP_INV_G8
XG2360 sck_bar XI11_6/XI3/net018 DECAP_INV_G9
XG2361 XI11_6/XI3/net018 XI11_6/XI3/net012 DECAP_INV_G9
XG2362 XI11_6/XI3/net014 XI11_6/XI3/net7 DECAP_INV_G9
XG2363 XI11_6/XI3/net012 XI11_6/XI3/net014 DECAP_INV_G9
XG2364 XI11_6/XI4/net063 XI11_6/XI4/net0112 DECAP_INV_G10
XG2365 XI11_6/XI4/net26 XI11_6/XI4/net089 DECAP_INV_G10
XG2366 XI11_6/XI4/data_out XI11_6/XI4/data_out_ DECAP_INV_G10
XG2367 XI11_6/XI4/net20 XI11_6/XI4/net0103 DECAP_INV_G10
XG2368 XI11_6/net12 XI11_6/XI4/net32 DECAP_INV_G7
XG2369 XI11_6/net9 XI11_6/XI4/net52 DECAP_INV_G7
XG2370 XI11_6/XI4/data_out_ XI11_6/XI4/data_out DECAP_INV_G10
XG2371 XI11_6/XI0/XI0_63/d__15_ XI11_6/XI0/XI0_63/d_15_ DECAP_INV_G11
XG2372 XI11_6/XI0/XI0_63/d__14_ XI11_6/XI0/XI0_63/d_14_ DECAP_INV_G11
XG2373 XI11_6/XI0/XI0_63/d__13_ XI11_6/XI0/XI0_63/d_13_ DECAP_INV_G11
XG2374 XI11_6/XI0/XI0_63/d__12_ XI11_6/XI0/XI0_63/d_12_ DECAP_INV_G11
XG2375 XI11_6/XI0/XI0_63/d__11_ XI11_6/XI0/XI0_63/d_11_ DECAP_INV_G11
XG2376 XI11_6/XI0/XI0_63/d__10_ XI11_6/XI0/XI0_63/d_10_ DECAP_INV_G11
XG2377 XI11_6/XI0/XI0_63/d__9_ XI11_6/XI0/XI0_63/d_9_ DECAP_INV_G11
XG2378 XI11_6/XI0/XI0_63/d__8_ XI11_6/XI0/XI0_63/d_8_ DECAP_INV_G11
XG2379 XI11_6/XI0/XI0_63/d__7_ XI11_6/XI0/XI0_63/d_7_ DECAP_INV_G11
XG2380 XI11_6/XI0/XI0_63/d__6_ XI11_6/XI0/XI0_63/d_6_ DECAP_INV_G11
XG2381 XI11_6/XI0/XI0_63/d__5_ XI11_6/XI0/XI0_63/d_5_ DECAP_INV_G11
XG2382 XI11_6/XI0/XI0_63/d__4_ XI11_6/XI0/XI0_63/d_4_ DECAP_INV_G11
XG2383 XI11_6/XI0/XI0_63/d__3_ XI11_6/XI0/XI0_63/d_3_ DECAP_INV_G11
XG2384 XI11_6/XI0/XI0_63/d__2_ XI11_6/XI0/XI0_63/d_2_ DECAP_INV_G11
XG2385 XI11_6/XI0/XI0_63/d__1_ XI11_6/XI0/XI0_63/d_1_ DECAP_INV_G11
XG2386 XI11_6/XI0/XI0_63/d__0_ XI11_6/XI0/XI0_63/d_0_ DECAP_INV_G11
XG2387 XI11_6/XI0/XI0_63/d_15_ XI11_6/XI0/XI0_63/d__15_ DECAP_INV_G11
XG2388 XI11_6/XI0/XI0_63/d_14_ XI11_6/XI0/XI0_63/d__14_ DECAP_INV_G11
XG2389 XI11_6/XI0/XI0_63/d_13_ XI11_6/XI0/XI0_63/d__13_ DECAP_INV_G11
XG2390 XI11_6/XI0/XI0_63/d_12_ XI11_6/XI0/XI0_63/d__12_ DECAP_INV_G11
XG2391 XI11_6/XI0/XI0_63/d_11_ XI11_6/XI0/XI0_63/d__11_ DECAP_INV_G11
XG2392 XI11_6/XI0/XI0_63/d_10_ XI11_6/XI0/XI0_63/d__10_ DECAP_INV_G11
XG2393 XI11_6/XI0/XI0_63/d_9_ XI11_6/XI0/XI0_63/d__9_ DECAP_INV_G11
XG2394 XI11_6/XI0/XI0_63/d_8_ XI11_6/XI0/XI0_63/d__8_ DECAP_INV_G11
XG2395 XI11_6/XI0/XI0_63/d_7_ XI11_6/XI0/XI0_63/d__7_ DECAP_INV_G11
XG2396 XI11_6/XI0/XI0_63/d_6_ XI11_6/XI0/XI0_63/d__6_ DECAP_INV_G11
XG2397 XI11_6/XI0/XI0_63/d_5_ XI11_6/XI0/XI0_63/d__5_ DECAP_INV_G11
XG2398 XI11_6/XI0/XI0_63/d_4_ XI11_6/XI0/XI0_63/d__4_ DECAP_INV_G11
XG2399 XI11_6/XI0/XI0_63/d_3_ XI11_6/XI0/XI0_63/d__3_ DECAP_INV_G11
XG2400 XI11_6/XI0/XI0_63/d_2_ XI11_6/XI0/XI0_63/d__2_ DECAP_INV_G11
XG2401 XI11_6/XI0/XI0_63/d_1_ XI11_6/XI0/XI0_63/d__1_ DECAP_INV_G11
XG2402 XI11_6/XI0/XI0_63/d_0_ XI11_6/XI0/XI0_63/d__0_ DECAP_INV_G11
XG2403 XI11_6/XI0/XI0_62/d__15_ XI11_6/XI0/XI0_62/d_15_ DECAP_INV_G11
XG2404 XI11_6/XI0/XI0_62/d__14_ XI11_6/XI0/XI0_62/d_14_ DECAP_INV_G11
XG2405 XI11_6/XI0/XI0_62/d__13_ XI11_6/XI0/XI0_62/d_13_ DECAP_INV_G11
XG2406 XI11_6/XI0/XI0_62/d__12_ XI11_6/XI0/XI0_62/d_12_ DECAP_INV_G11
XG2407 XI11_6/XI0/XI0_62/d__11_ XI11_6/XI0/XI0_62/d_11_ DECAP_INV_G11
XG2408 XI11_6/XI0/XI0_62/d__10_ XI11_6/XI0/XI0_62/d_10_ DECAP_INV_G11
XG2409 XI11_6/XI0/XI0_62/d__9_ XI11_6/XI0/XI0_62/d_9_ DECAP_INV_G11
XG2410 XI11_6/XI0/XI0_62/d__8_ XI11_6/XI0/XI0_62/d_8_ DECAP_INV_G11
XG2411 XI11_6/XI0/XI0_62/d__7_ XI11_6/XI0/XI0_62/d_7_ DECAP_INV_G11
XG2412 XI11_6/XI0/XI0_62/d__6_ XI11_6/XI0/XI0_62/d_6_ DECAP_INV_G11
XG2413 XI11_6/XI0/XI0_62/d__5_ XI11_6/XI0/XI0_62/d_5_ DECAP_INV_G11
XG2414 XI11_6/XI0/XI0_62/d__4_ XI11_6/XI0/XI0_62/d_4_ DECAP_INV_G11
XG2415 XI11_6/XI0/XI0_62/d__3_ XI11_6/XI0/XI0_62/d_3_ DECAP_INV_G11
XG2416 XI11_6/XI0/XI0_62/d__2_ XI11_6/XI0/XI0_62/d_2_ DECAP_INV_G11
XG2417 XI11_6/XI0/XI0_62/d__1_ XI11_6/XI0/XI0_62/d_1_ DECAP_INV_G11
XG2418 XI11_6/XI0/XI0_62/d__0_ XI11_6/XI0/XI0_62/d_0_ DECAP_INV_G11
XG2419 XI11_6/XI0/XI0_62/d_15_ XI11_6/XI0/XI0_62/d__15_ DECAP_INV_G11
XG2420 XI11_6/XI0/XI0_62/d_14_ XI11_6/XI0/XI0_62/d__14_ DECAP_INV_G11
XG2421 XI11_6/XI0/XI0_62/d_13_ XI11_6/XI0/XI0_62/d__13_ DECAP_INV_G11
XG2422 XI11_6/XI0/XI0_62/d_12_ XI11_6/XI0/XI0_62/d__12_ DECAP_INV_G11
XG2423 XI11_6/XI0/XI0_62/d_11_ XI11_6/XI0/XI0_62/d__11_ DECAP_INV_G11
XG2424 XI11_6/XI0/XI0_62/d_10_ XI11_6/XI0/XI0_62/d__10_ DECAP_INV_G11
XG2425 XI11_6/XI0/XI0_62/d_9_ XI11_6/XI0/XI0_62/d__9_ DECAP_INV_G11
XG2426 XI11_6/XI0/XI0_62/d_8_ XI11_6/XI0/XI0_62/d__8_ DECAP_INV_G11
XG2427 XI11_6/XI0/XI0_62/d_7_ XI11_6/XI0/XI0_62/d__7_ DECAP_INV_G11
XG2428 XI11_6/XI0/XI0_62/d_6_ XI11_6/XI0/XI0_62/d__6_ DECAP_INV_G11
XG2429 XI11_6/XI0/XI0_62/d_5_ XI11_6/XI0/XI0_62/d__5_ DECAP_INV_G11
XG2430 XI11_6/XI0/XI0_62/d_4_ XI11_6/XI0/XI0_62/d__4_ DECAP_INV_G11
XG2431 XI11_6/XI0/XI0_62/d_3_ XI11_6/XI0/XI0_62/d__3_ DECAP_INV_G11
XG2432 XI11_6/XI0/XI0_62/d_2_ XI11_6/XI0/XI0_62/d__2_ DECAP_INV_G11
XG2433 XI11_6/XI0/XI0_62/d_1_ XI11_6/XI0/XI0_62/d__1_ DECAP_INV_G11
XG2434 XI11_6/XI0/XI0_62/d_0_ XI11_6/XI0/XI0_62/d__0_ DECAP_INV_G11
XG2435 XI11_6/XI0/XI0_61/d__15_ XI11_6/XI0/XI0_61/d_15_ DECAP_INV_G11
XG2436 XI11_6/XI0/XI0_61/d__14_ XI11_6/XI0/XI0_61/d_14_ DECAP_INV_G11
XG2437 XI11_6/XI0/XI0_61/d__13_ XI11_6/XI0/XI0_61/d_13_ DECAP_INV_G11
XG2438 XI11_6/XI0/XI0_61/d__12_ XI11_6/XI0/XI0_61/d_12_ DECAP_INV_G11
XG2439 XI11_6/XI0/XI0_61/d__11_ XI11_6/XI0/XI0_61/d_11_ DECAP_INV_G11
XG2440 XI11_6/XI0/XI0_61/d__10_ XI11_6/XI0/XI0_61/d_10_ DECAP_INV_G11
XG2441 XI11_6/XI0/XI0_61/d__9_ XI11_6/XI0/XI0_61/d_9_ DECAP_INV_G11
XG2442 XI11_6/XI0/XI0_61/d__8_ XI11_6/XI0/XI0_61/d_8_ DECAP_INV_G11
XG2443 XI11_6/XI0/XI0_61/d__7_ XI11_6/XI0/XI0_61/d_7_ DECAP_INV_G11
XG2444 XI11_6/XI0/XI0_61/d__6_ XI11_6/XI0/XI0_61/d_6_ DECAP_INV_G11
XG2445 XI11_6/XI0/XI0_61/d__5_ XI11_6/XI0/XI0_61/d_5_ DECAP_INV_G11
XG2446 XI11_6/XI0/XI0_61/d__4_ XI11_6/XI0/XI0_61/d_4_ DECAP_INV_G11
XG2447 XI11_6/XI0/XI0_61/d__3_ XI11_6/XI0/XI0_61/d_3_ DECAP_INV_G11
XG2448 XI11_6/XI0/XI0_61/d__2_ XI11_6/XI0/XI0_61/d_2_ DECAP_INV_G11
XG2449 XI11_6/XI0/XI0_61/d__1_ XI11_6/XI0/XI0_61/d_1_ DECAP_INV_G11
XG2450 XI11_6/XI0/XI0_61/d__0_ XI11_6/XI0/XI0_61/d_0_ DECAP_INV_G11
XG2451 XI11_6/XI0/XI0_61/d_15_ XI11_6/XI0/XI0_61/d__15_ DECAP_INV_G11
XG2452 XI11_6/XI0/XI0_61/d_14_ XI11_6/XI0/XI0_61/d__14_ DECAP_INV_G11
XG2453 XI11_6/XI0/XI0_61/d_13_ XI11_6/XI0/XI0_61/d__13_ DECAP_INV_G11
XG2454 XI11_6/XI0/XI0_61/d_12_ XI11_6/XI0/XI0_61/d__12_ DECAP_INV_G11
XG2455 XI11_6/XI0/XI0_61/d_11_ XI11_6/XI0/XI0_61/d__11_ DECAP_INV_G11
XG2456 XI11_6/XI0/XI0_61/d_10_ XI11_6/XI0/XI0_61/d__10_ DECAP_INV_G11
XG2457 XI11_6/XI0/XI0_61/d_9_ XI11_6/XI0/XI0_61/d__9_ DECAP_INV_G11
XG2458 XI11_6/XI0/XI0_61/d_8_ XI11_6/XI0/XI0_61/d__8_ DECAP_INV_G11
XG2459 XI11_6/XI0/XI0_61/d_7_ XI11_6/XI0/XI0_61/d__7_ DECAP_INV_G11
XG2460 XI11_6/XI0/XI0_61/d_6_ XI11_6/XI0/XI0_61/d__6_ DECAP_INV_G11
XG2461 XI11_6/XI0/XI0_61/d_5_ XI11_6/XI0/XI0_61/d__5_ DECAP_INV_G11
XG2462 XI11_6/XI0/XI0_61/d_4_ XI11_6/XI0/XI0_61/d__4_ DECAP_INV_G11
XG2463 XI11_6/XI0/XI0_61/d_3_ XI11_6/XI0/XI0_61/d__3_ DECAP_INV_G11
XG2464 XI11_6/XI0/XI0_61/d_2_ XI11_6/XI0/XI0_61/d__2_ DECAP_INV_G11
XG2465 XI11_6/XI0/XI0_61/d_1_ XI11_6/XI0/XI0_61/d__1_ DECAP_INV_G11
XG2466 XI11_6/XI0/XI0_61/d_0_ XI11_6/XI0/XI0_61/d__0_ DECAP_INV_G11
XG2467 XI11_6/XI0/XI0_60/d__15_ XI11_6/XI0/XI0_60/d_15_ DECAP_INV_G11
XG2468 XI11_6/XI0/XI0_60/d__14_ XI11_6/XI0/XI0_60/d_14_ DECAP_INV_G11
XG2469 XI11_6/XI0/XI0_60/d__13_ XI11_6/XI0/XI0_60/d_13_ DECAP_INV_G11
XG2470 XI11_6/XI0/XI0_60/d__12_ XI11_6/XI0/XI0_60/d_12_ DECAP_INV_G11
XG2471 XI11_6/XI0/XI0_60/d__11_ XI11_6/XI0/XI0_60/d_11_ DECAP_INV_G11
XG2472 XI11_6/XI0/XI0_60/d__10_ XI11_6/XI0/XI0_60/d_10_ DECAP_INV_G11
XG2473 XI11_6/XI0/XI0_60/d__9_ XI11_6/XI0/XI0_60/d_9_ DECAP_INV_G11
XG2474 XI11_6/XI0/XI0_60/d__8_ XI11_6/XI0/XI0_60/d_8_ DECAP_INV_G11
XG2475 XI11_6/XI0/XI0_60/d__7_ XI11_6/XI0/XI0_60/d_7_ DECAP_INV_G11
XG2476 XI11_6/XI0/XI0_60/d__6_ XI11_6/XI0/XI0_60/d_6_ DECAP_INV_G11
XG2477 XI11_6/XI0/XI0_60/d__5_ XI11_6/XI0/XI0_60/d_5_ DECAP_INV_G11
XG2478 XI11_6/XI0/XI0_60/d__4_ XI11_6/XI0/XI0_60/d_4_ DECAP_INV_G11
XG2479 XI11_6/XI0/XI0_60/d__3_ XI11_6/XI0/XI0_60/d_3_ DECAP_INV_G11
XG2480 XI11_6/XI0/XI0_60/d__2_ XI11_6/XI0/XI0_60/d_2_ DECAP_INV_G11
XG2481 XI11_6/XI0/XI0_60/d__1_ XI11_6/XI0/XI0_60/d_1_ DECAP_INV_G11
XG2482 XI11_6/XI0/XI0_60/d__0_ XI11_6/XI0/XI0_60/d_0_ DECAP_INV_G11
XG2483 XI11_6/XI0/XI0_60/d_15_ XI11_6/XI0/XI0_60/d__15_ DECAP_INV_G11
XG2484 XI11_6/XI0/XI0_60/d_14_ XI11_6/XI0/XI0_60/d__14_ DECAP_INV_G11
XG2485 XI11_6/XI0/XI0_60/d_13_ XI11_6/XI0/XI0_60/d__13_ DECAP_INV_G11
XG2486 XI11_6/XI0/XI0_60/d_12_ XI11_6/XI0/XI0_60/d__12_ DECAP_INV_G11
XG2487 XI11_6/XI0/XI0_60/d_11_ XI11_6/XI0/XI0_60/d__11_ DECAP_INV_G11
XG2488 XI11_6/XI0/XI0_60/d_10_ XI11_6/XI0/XI0_60/d__10_ DECAP_INV_G11
XG2489 XI11_6/XI0/XI0_60/d_9_ XI11_6/XI0/XI0_60/d__9_ DECAP_INV_G11
XG2490 XI11_6/XI0/XI0_60/d_8_ XI11_6/XI0/XI0_60/d__8_ DECAP_INV_G11
XG2491 XI11_6/XI0/XI0_60/d_7_ XI11_6/XI0/XI0_60/d__7_ DECAP_INV_G11
XG2492 XI11_6/XI0/XI0_60/d_6_ XI11_6/XI0/XI0_60/d__6_ DECAP_INV_G11
XG2493 XI11_6/XI0/XI0_60/d_5_ XI11_6/XI0/XI0_60/d__5_ DECAP_INV_G11
XG2494 XI11_6/XI0/XI0_60/d_4_ XI11_6/XI0/XI0_60/d__4_ DECAP_INV_G11
XG2495 XI11_6/XI0/XI0_60/d_3_ XI11_6/XI0/XI0_60/d__3_ DECAP_INV_G11
XG2496 XI11_6/XI0/XI0_60/d_2_ XI11_6/XI0/XI0_60/d__2_ DECAP_INV_G11
XG2497 XI11_6/XI0/XI0_60/d_1_ XI11_6/XI0/XI0_60/d__1_ DECAP_INV_G11
XG2498 XI11_6/XI0/XI0_60/d_0_ XI11_6/XI0/XI0_60/d__0_ DECAP_INV_G11
XG2499 XI11_6/XI0/XI0_59/d__15_ XI11_6/XI0/XI0_59/d_15_ DECAP_INV_G11
XG2500 XI11_6/XI0/XI0_59/d__14_ XI11_6/XI0/XI0_59/d_14_ DECAP_INV_G11
XG2501 XI11_6/XI0/XI0_59/d__13_ XI11_6/XI0/XI0_59/d_13_ DECAP_INV_G11
XG2502 XI11_6/XI0/XI0_59/d__12_ XI11_6/XI0/XI0_59/d_12_ DECAP_INV_G11
XG2503 XI11_6/XI0/XI0_59/d__11_ XI11_6/XI0/XI0_59/d_11_ DECAP_INV_G11
XG2504 XI11_6/XI0/XI0_59/d__10_ XI11_6/XI0/XI0_59/d_10_ DECAP_INV_G11
XG2505 XI11_6/XI0/XI0_59/d__9_ XI11_6/XI0/XI0_59/d_9_ DECAP_INV_G11
XG2506 XI11_6/XI0/XI0_59/d__8_ XI11_6/XI0/XI0_59/d_8_ DECAP_INV_G11
XG2507 XI11_6/XI0/XI0_59/d__7_ XI11_6/XI0/XI0_59/d_7_ DECAP_INV_G11
XG2508 XI11_6/XI0/XI0_59/d__6_ XI11_6/XI0/XI0_59/d_6_ DECAP_INV_G11
XG2509 XI11_6/XI0/XI0_59/d__5_ XI11_6/XI0/XI0_59/d_5_ DECAP_INV_G11
XG2510 XI11_6/XI0/XI0_59/d__4_ XI11_6/XI0/XI0_59/d_4_ DECAP_INV_G11
XG2511 XI11_6/XI0/XI0_59/d__3_ XI11_6/XI0/XI0_59/d_3_ DECAP_INV_G11
XG2512 XI11_6/XI0/XI0_59/d__2_ XI11_6/XI0/XI0_59/d_2_ DECAP_INV_G11
XG2513 XI11_6/XI0/XI0_59/d__1_ XI11_6/XI0/XI0_59/d_1_ DECAP_INV_G11
XG2514 XI11_6/XI0/XI0_59/d__0_ XI11_6/XI0/XI0_59/d_0_ DECAP_INV_G11
XG2515 XI11_6/XI0/XI0_59/d_15_ XI11_6/XI0/XI0_59/d__15_ DECAP_INV_G11
XG2516 XI11_6/XI0/XI0_59/d_14_ XI11_6/XI0/XI0_59/d__14_ DECAP_INV_G11
XG2517 XI11_6/XI0/XI0_59/d_13_ XI11_6/XI0/XI0_59/d__13_ DECAP_INV_G11
XG2518 XI11_6/XI0/XI0_59/d_12_ XI11_6/XI0/XI0_59/d__12_ DECAP_INV_G11
XG2519 XI11_6/XI0/XI0_59/d_11_ XI11_6/XI0/XI0_59/d__11_ DECAP_INV_G11
XG2520 XI11_6/XI0/XI0_59/d_10_ XI11_6/XI0/XI0_59/d__10_ DECAP_INV_G11
XG2521 XI11_6/XI0/XI0_59/d_9_ XI11_6/XI0/XI0_59/d__9_ DECAP_INV_G11
XG2522 XI11_6/XI0/XI0_59/d_8_ XI11_6/XI0/XI0_59/d__8_ DECAP_INV_G11
XG2523 XI11_6/XI0/XI0_59/d_7_ XI11_6/XI0/XI0_59/d__7_ DECAP_INV_G11
XG2524 XI11_6/XI0/XI0_59/d_6_ XI11_6/XI0/XI0_59/d__6_ DECAP_INV_G11
XG2525 XI11_6/XI0/XI0_59/d_5_ XI11_6/XI0/XI0_59/d__5_ DECAP_INV_G11
XG2526 XI11_6/XI0/XI0_59/d_4_ XI11_6/XI0/XI0_59/d__4_ DECAP_INV_G11
XG2527 XI11_6/XI0/XI0_59/d_3_ XI11_6/XI0/XI0_59/d__3_ DECAP_INV_G11
XG2528 XI11_6/XI0/XI0_59/d_2_ XI11_6/XI0/XI0_59/d__2_ DECAP_INV_G11
XG2529 XI11_6/XI0/XI0_59/d_1_ XI11_6/XI0/XI0_59/d__1_ DECAP_INV_G11
XG2530 XI11_6/XI0/XI0_59/d_0_ XI11_6/XI0/XI0_59/d__0_ DECAP_INV_G11
XG2531 XI11_6/XI0/XI0_58/d__15_ XI11_6/XI0/XI0_58/d_15_ DECAP_INV_G11
XG2532 XI11_6/XI0/XI0_58/d__14_ XI11_6/XI0/XI0_58/d_14_ DECAP_INV_G11
XG2533 XI11_6/XI0/XI0_58/d__13_ XI11_6/XI0/XI0_58/d_13_ DECAP_INV_G11
XG2534 XI11_6/XI0/XI0_58/d__12_ XI11_6/XI0/XI0_58/d_12_ DECAP_INV_G11
XG2535 XI11_6/XI0/XI0_58/d__11_ XI11_6/XI0/XI0_58/d_11_ DECAP_INV_G11
XG2536 XI11_6/XI0/XI0_58/d__10_ XI11_6/XI0/XI0_58/d_10_ DECAP_INV_G11
XG2537 XI11_6/XI0/XI0_58/d__9_ XI11_6/XI0/XI0_58/d_9_ DECAP_INV_G11
XG2538 XI11_6/XI0/XI0_58/d__8_ XI11_6/XI0/XI0_58/d_8_ DECAP_INV_G11
XG2539 XI11_6/XI0/XI0_58/d__7_ XI11_6/XI0/XI0_58/d_7_ DECAP_INV_G11
XG2540 XI11_6/XI0/XI0_58/d__6_ XI11_6/XI0/XI0_58/d_6_ DECAP_INV_G11
XG2541 XI11_6/XI0/XI0_58/d__5_ XI11_6/XI0/XI0_58/d_5_ DECAP_INV_G11
XG2542 XI11_6/XI0/XI0_58/d__4_ XI11_6/XI0/XI0_58/d_4_ DECAP_INV_G11
XG2543 XI11_6/XI0/XI0_58/d__3_ XI11_6/XI0/XI0_58/d_3_ DECAP_INV_G11
XG2544 XI11_6/XI0/XI0_58/d__2_ XI11_6/XI0/XI0_58/d_2_ DECAP_INV_G11
XG2545 XI11_6/XI0/XI0_58/d__1_ XI11_6/XI0/XI0_58/d_1_ DECAP_INV_G11
XG2546 XI11_6/XI0/XI0_58/d__0_ XI11_6/XI0/XI0_58/d_0_ DECAP_INV_G11
XG2547 XI11_6/XI0/XI0_58/d_15_ XI11_6/XI0/XI0_58/d__15_ DECAP_INV_G11
XG2548 XI11_6/XI0/XI0_58/d_14_ XI11_6/XI0/XI0_58/d__14_ DECAP_INV_G11
XG2549 XI11_6/XI0/XI0_58/d_13_ XI11_6/XI0/XI0_58/d__13_ DECAP_INV_G11
XG2550 XI11_6/XI0/XI0_58/d_12_ XI11_6/XI0/XI0_58/d__12_ DECAP_INV_G11
XG2551 XI11_6/XI0/XI0_58/d_11_ XI11_6/XI0/XI0_58/d__11_ DECAP_INV_G11
XG2552 XI11_6/XI0/XI0_58/d_10_ XI11_6/XI0/XI0_58/d__10_ DECAP_INV_G11
XG2553 XI11_6/XI0/XI0_58/d_9_ XI11_6/XI0/XI0_58/d__9_ DECAP_INV_G11
XG2554 XI11_6/XI0/XI0_58/d_8_ XI11_6/XI0/XI0_58/d__8_ DECAP_INV_G11
XG2555 XI11_6/XI0/XI0_58/d_7_ XI11_6/XI0/XI0_58/d__7_ DECAP_INV_G11
XG2556 XI11_6/XI0/XI0_58/d_6_ XI11_6/XI0/XI0_58/d__6_ DECAP_INV_G11
XG2557 XI11_6/XI0/XI0_58/d_5_ XI11_6/XI0/XI0_58/d__5_ DECAP_INV_G11
XG2558 XI11_6/XI0/XI0_58/d_4_ XI11_6/XI0/XI0_58/d__4_ DECAP_INV_G11
XG2559 XI11_6/XI0/XI0_58/d_3_ XI11_6/XI0/XI0_58/d__3_ DECAP_INV_G11
XG2560 XI11_6/XI0/XI0_58/d_2_ XI11_6/XI0/XI0_58/d__2_ DECAP_INV_G11
XG2561 XI11_6/XI0/XI0_58/d_1_ XI11_6/XI0/XI0_58/d__1_ DECAP_INV_G11
XG2562 XI11_6/XI0/XI0_58/d_0_ XI11_6/XI0/XI0_58/d__0_ DECAP_INV_G11
XG2563 XI11_6/XI0/XI0_57/d__15_ XI11_6/XI0/XI0_57/d_15_ DECAP_INV_G11
XG2564 XI11_6/XI0/XI0_57/d__14_ XI11_6/XI0/XI0_57/d_14_ DECAP_INV_G11
XG2565 XI11_6/XI0/XI0_57/d__13_ XI11_6/XI0/XI0_57/d_13_ DECAP_INV_G11
XG2566 XI11_6/XI0/XI0_57/d__12_ XI11_6/XI0/XI0_57/d_12_ DECAP_INV_G11
XG2567 XI11_6/XI0/XI0_57/d__11_ XI11_6/XI0/XI0_57/d_11_ DECAP_INV_G11
XG2568 XI11_6/XI0/XI0_57/d__10_ XI11_6/XI0/XI0_57/d_10_ DECAP_INV_G11
XG2569 XI11_6/XI0/XI0_57/d__9_ XI11_6/XI0/XI0_57/d_9_ DECAP_INV_G11
XG2570 XI11_6/XI0/XI0_57/d__8_ XI11_6/XI0/XI0_57/d_8_ DECAP_INV_G11
XG2571 XI11_6/XI0/XI0_57/d__7_ XI11_6/XI0/XI0_57/d_7_ DECAP_INV_G11
XG2572 XI11_6/XI0/XI0_57/d__6_ XI11_6/XI0/XI0_57/d_6_ DECAP_INV_G11
XG2573 XI11_6/XI0/XI0_57/d__5_ XI11_6/XI0/XI0_57/d_5_ DECAP_INV_G11
XG2574 XI11_6/XI0/XI0_57/d__4_ XI11_6/XI0/XI0_57/d_4_ DECAP_INV_G11
XG2575 XI11_6/XI0/XI0_57/d__3_ XI11_6/XI0/XI0_57/d_3_ DECAP_INV_G11
XG2576 XI11_6/XI0/XI0_57/d__2_ XI11_6/XI0/XI0_57/d_2_ DECAP_INV_G11
XG2577 XI11_6/XI0/XI0_57/d__1_ XI11_6/XI0/XI0_57/d_1_ DECAP_INV_G11
XG2578 XI11_6/XI0/XI0_57/d__0_ XI11_6/XI0/XI0_57/d_0_ DECAP_INV_G11
XG2579 XI11_6/XI0/XI0_57/d_15_ XI11_6/XI0/XI0_57/d__15_ DECAP_INV_G11
XG2580 XI11_6/XI0/XI0_57/d_14_ XI11_6/XI0/XI0_57/d__14_ DECAP_INV_G11
XG2581 XI11_6/XI0/XI0_57/d_13_ XI11_6/XI0/XI0_57/d__13_ DECAP_INV_G11
XG2582 XI11_6/XI0/XI0_57/d_12_ XI11_6/XI0/XI0_57/d__12_ DECAP_INV_G11
XG2583 XI11_6/XI0/XI0_57/d_11_ XI11_6/XI0/XI0_57/d__11_ DECAP_INV_G11
XG2584 XI11_6/XI0/XI0_57/d_10_ XI11_6/XI0/XI0_57/d__10_ DECAP_INV_G11
XG2585 XI11_6/XI0/XI0_57/d_9_ XI11_6/XI0/XI0_57/d__9_ DECAP_INV_G11
XG2586 XI11_6/XI0/XI0_57/d_8_ XI11_6/XI0/XI0_57/d__8_ DECAP_INV_G11
XG2587 XI11_6/XI0/XI0_57/d_7_ XI11_6/XI0/XI0_57/d__7_ DECAP_INV_G11
XG2588 XI11_6/XI0/XI0_57/d_6_ XI11_6/XI0/XI0_57/d__6_ DECAP_INV_G11
XG2589 XI11_6/XI0/XI0_57/d_5_ XI11_6/XI0/XI0_57/d__5_ DECAP_INV_G11
XG2590 XI11_6/XI0/XI0_57/d_4_ XI11_6/XI0/XI0_57/d__4_ DECAP_INV_G11
XG2591 XI11_6/XI0/XI0_57/d_3_ XI11_6/XI0/XI0_57/d__3_ DECAP_INV_G11
XG2592 XI11_6/XI0/XI0_57/d_2_ XI11_6/XI0/XI0_57/d__2_ DECAP_INV_G11
XG2593 XI11_6/XI0/XI0_57/d_1_ XI11_6/XI0/XI0_57/d__1_ DECAP_INV_G11
XG2594 XI11_6/XI0/XI0_57/d_0_ XI11_6/XI0/XI0_57/d__0_ DECAP_INV_G11
XG2595 XI11_6/XI0/XI0_56/d__15_ XI11_6/XI0/XI0_56/d_15_ DECAP_INV_G11
XG2596 XI11_6/XI0/XI0_56/d__14_ XI11_6/XI0/XI0_56/d_14_ DECAP_INV_G11
XG2597 XI11_6/XI0/XI0_56/d__13_ XI11_6/XI0/XI0_56/d_13_ DECAP_INV_G11
XG2598 XI11_6/XI0/XI0_56/d__12_ XI11_6/XI0/XI0_56/d_12_ DECAP_INV_G11
XG2599 XI11_6/XI0/XI0_56/d__11_ XI11_6/XI0/XI0_56/d_11_ DECAP_INV_G11
XG2600 XI11_6/XI0/XI0_56/d__10_ XI11_6/XI0/XI0_56/d_10_ DECAP_INV_G11
XG2601 XI11_6/XI0/XI0_56/d__9_ XI11_6/XI0/XI0_56/d_9_ DECAP_INV_G11
XG2602 XI11_6/XI0/XI0_56/d__8_ XI11_6/XI0/XI0_56/d_8_ DECAP_INV_G11
XG2603 XI11_6/XI0/XI0_56/d__7_ XI11_6/XI0/XI0_56/d_7_ DECAP_INV_G11
XG2604 XI11_6/XI0/XI0_56/d__6_ XI11_6/XI0/XI0_56/d_6_ DECAP_INV_G11
XG2605 XI11_6/XI0/XI0_56/d__5_ XI11_6/XI0/XI0_56/d_5_ DECAP_INV_G11
XG2606 XI11_6/XI0/XI0_56/d__4_ XI11_6/XI0/XI0_56/d_4_ DECAP_INV_G11
XG2607 XI11_6/XI0/XI0_56/d__3_ XI11_6/XI0/XI0_56/d_3_ DECAP_INV_G11
XG2608 XI11_6/XI0/XI0_56/d__2_ XI11_6/XI0/XI0_56/d_2_ DECAP_INV_G11
XG2609 XI11_6/XI0/XI0_56/d__1_ XI11_6/XI0/XI0_56/d_1_ DECAP_INV_G11
XG2610 XI11_6/XI0/XI0_56/d__0_ XI11_6/XI0/XI0_56/d_0_ DECAP_INV_G11
XG2611 XI11_6/XI0/XI0_56/d_15_ XI11_6/XI0/XI0_56/d__15_ DECAP_INV_G11
XG2612 XI11_6/XI0/XI0_56/d_14_ XI11_6/XI0/XI0_56/d__14_ DECAP_INV_G11
XG2613 XI11_6/XI0/XI0_56/d_13_ XI11_6/XI0/XI0_56/d__13_ DECAP_INV_G11
XG2614 XI11_6/XI0/XI0_56/d_12_ XI11_6/XI0/XI0_56/d__12_ DECAP_INV_G11
XG2615 XI11_6/XI0/XI0_56/d_11_ XI11_6/XI0/XI0_56/d__11_ DECAP_INV_G11
XG2616 XI11_6/XI0/XI0_56/d_10_ XI11_6/XI0/XI0_56/d__10_ DECAP_INV_G11
XG2617 XI11_6/XI0/XI0_56/d_9_ XI11_6/XI0/XI0_56/d__9_ DECAP_INV_G11
XG2618 XI11_6/XI0/XI0_56/d_8_ XI11_6/XI0/XI0_56/d__8_ DECAP_INV_G11
XG2619 XI11_6/XI0/XI0_56/d_7_ XI11_6/XI0/XI0_56/d__7_ DECAP_INV_G11
XG2620 XI11_6/XI0/XI0_56/d_6_ XI11_6/XI0/XI0_56/d__6_ DECAP_INV_G11
XG2621 XI11_6/XI0/XI0_56/d_5_ XI11_6/XI0/XI0_56/d__5_ DECAP_INV_G11
XG2622 XI11_6/XI0/XI0_56/d_4_ XI11_6/XI0/XI0_56/d__4_ DECAP_INV_G11
XG2623 XI11_6/XI0/XI0_56/d_3_ XI11_6/XI0/XI0_56/d__3_ DECAP_INV_G11
XG2624 XI11_6/XI0/XI0_56/d_2_ XI11_6/XI0/XI0_56/d__2_ DECAP_INV_G11
XG2625 XI11_6/XI0/XI0_56/d_1_ XI11_6/XI0/XI0_56/d__1_ DECAP_INV_G11
XG2626 XI11_6/XI0/XI0_56/d_0_ XI11_6/XI0/XI0_56/d__0_ DECAP_INV_G11
XG2627 XI11_6/XI0/XI0_55/d__15_ XI11_6/XI0/XI0_55/d_15_ DECAP_INV_G11
XG2628 XI11_6/XI0/XI0_55/d__14_ XI11_6/XI0/XI0_55/d_14_ DECAP_INV_G11
XG2629 XI11_6/XI0/XI0_55/d__13_ XI11_6/XI0/XI0_55/d_13_ DECAP_INV_G11
XG2630 XI11_6/XI0/XI0_55/d__12_ XI11_6/XI0/XI0_55/d_12_ DECAP_INV_G11
XG2631 XI11_6/XI0/XI0_55/d__11_ XI11_6/XI0/XI0_55/d_11_ DECAP_INV_G11
XG2632 XI11_6/XI0/XI0_55/d__10_ XI11_6/XI0/XI0_55/d_10_ DECAP_INV_G11
XG2633 XI11_6/XI0/XI0_55/d__9_ XI11_6/XI0/XI0_55/d_9_ DECAP_INV_G11
XG2634 XI11_6/XI0/XI0_55/d__8_ XI11_6/XI0/XI0_55/d_8_ DECAP_INV_G11
XG2635 XI11_6/XI0/XI0_55/d__7_ XI11_6/XI0/XI0_55/d_7_ DECAP_INV_G11
XG2636 XI11_6/XI0/XI0_55/d__6_ XI11_6/XI0/XI0_55/d_6_ DECAP_INV_G11
XG2637 XI11_6/XI0/XI0_55/d__5_ XI11_6/XI0/XI0_55/d_5_ DECAP_INV_G11
XG2638 XI11_6/XI0/XI0_55/d__4_ XI11_6/XI0/XI0_55/d_4_ DECAP_INV_G11
XG2639 XI11_6/XI0/XI0_55/d__3_ XI11_6/XI0/XI0_55/d_3_ DECAP_INV_G11
XG2640 XI11_6/XI0/XI0_55/d__2_ XI11_6/XI0/XI0_55/d_2_ DECAP_INV_G11
XG2641 XI11_6/XI0/XI0_55/d__1_ XI11_6/XI0/XI0_55/d_1_ DECAP_INV_G11
XG2642 XI11_6/XI0/XI0_55/d__0_ XI11_6/XI0/XI0_55/d_0_ DECAP_INV_G11
XG2643 XI11_6/XI0/XI0_55/d_15_ XI11_6/XI0/XI0_55/d__15_ DECAP_INV_G11
XG2644 XI11_6/XI0/XI0_55/d_14_ XI11_6/XI0/XI0_55/d__14_ DECAP_INV_G11
XG2645 XI11_6/XI0/XI0_55/d_13_ XI11_6/XI0/XI0_55/d__13_ DECAP_INV_G11
XG2646 XI11_6/XI0/XI0_55/d_12_ XI11_6/XI0/XI0_55/d__12_ DECAP_INV_G11
XG2647 XI11_6/XI0/XI0_55/d_11_ XI11_6/XI0/XI0_55/d__11_ DECAP_INV_G11
XG2648 XI11_6/XI0/XI0_55/d_10_ XI11_6/XI0/XI0_55/d__10_ DECAP_INV_G11
XG2649 XI11_6/XI0/XI0_55/d_9_ XI11_6/XI0/XI0_55/d__9_ DECAP_INV_G11
XG2650 XI11_6/XI0/XI0_55/d_8_ XI11_6/XI0/XI0_55/d__8_ DECAP_INV_G11
XG2651 XI11_6/XI0/XI0_55/d_7_ XI11_6/XI0/XI0_55/d__7_ DECAP_INV_G11
XG2652 XI11_6/XI0/XI0_55/d_6_ XI11_6/XI0/XI0_55/d__6_ DECAP_INV_G11
XG2653 XI11_6/XI0/XI0_55/d_5_ XI11_6/XI0/XI0_55/d__5_ DECAP_INV_G11
XG2654 XI11_6/XI0/XI0_55/d_4_ XI11_6/XI0/XI0_55/d__4_ DECAP_INV_G11
XG2655 XI11_6/XI0/XI0_55/d_3_ XI11_6/XI0/XI0_55/d__3_ DECAP_INV_G11
XG2656 XI11_6/XI0/XI0_55/d_2_ XI11_6/XI0/XI0_55/d__2_ DECAP_INV_G11
XG2657 XI11_6/XI0/XI0_55/d_1_ XI11_6/XI0/XI0_55/d__1_ DECAP_INV_G11
XG2658 XI11_6/XI0/XI0_55/d_0_ XI11_6/XI0/XI0_55/d__0_ DECAP_INV_G11
XG2659 XI11_6/XI0/XI0_54/d__15_ XI11_6/XI0/XI0_54/d_15_ DECAP_INV_G11
XG2660 XI11_6/XI0/XI0_54/d__14_ XI11_6/XI0/XI0_54/d_14_ DECAP_INV_G11
XG2661 XI11_6/XI0/XI0_54/d__13_ XI11_6/XI0/XI0_54/d_13_ DECAP_INV_G11
XG2662 XI11_6/XI0/XI0_54/d__12_ XI11_6/XI0/XI0_54/d_12_ DECAP_INV_G11
XG2663 XI11_6/XI0/XI0_54/d__11_ XI11_6/XI0/XI0_54/d_11_ DECAP_INV_G11
XG2664 XI11_6/XI0/XI0_54/d__10_ XI11_6/XI0/XI0_54/d_10_ DECAP_INV_G11
XG2665 XI11_6/XI0/XI0_54/d__9_ XI11_6/XI0/XI0_54/d_9_ DECAP_INV_G11
XG2666 XI11_6/XI0/XI0_54/d__8_ XI11_6/XI0/XI0_54/d_8_ DECAP_INV_G11
XG2667 XI11_6/XI0/XI0_54/d__7_ XI11_6/XI0/XI0_54/d_7_ DECAP_INV_G11
XG2668 XI11_6/XI0/XI0_54/d__6_ XI11_6/XI0/XI0_54/d_6_ DECAP_INV_G11
XG2669 XI11_6/XI0/XI0_54/d__5_ XI11_6/XI0/XI0_54/d_5_ DECAP_INV_G11
XG2670 XI11_6/XI0/XI0_54/d__4_ XI11_6/XI0/XI0_54/d_4_ DECAP_INV_G11
XG2671 XI11_6/XI0/XI0_54/d__3_ XI11_6/XI0/XI0_54/d_3_ DECAP_INV_G11
XG2672 XI11_6/XI0/XI0_54/d__2_ XI11_6/XI0/XI0_54/d_2_ DECAP_INV_G11
XG2673 XI11_6/XI0/XI0_54/d__1_ XI11_6/XI0/XI0_54/d_1_ DECAP_INV_G11
XG2674 XI11_6/XI0/XI0_54/d__0_ XI11_6/XI0/XI0_54/d_0_ DECAP_INV_G11
XG2675 XI11_6/XI0/XI0_54/d_15_ XI11_6/XI0/XI0_54/d__15_ DECAP_INV_G11
XG2676 XI11_6/XI0/XI0_54/d_14_ XI11_6/XI0/XI0_54/d__14_ DECAP_INV_G11
XG2677 XI11_6/XI0/XI0_54/d_13_ XI11_6/XI0/XI0_54/d__13_ DECAP_INV_G11
XG2678 XI11_6/XI0/XI0_54/d_12_ XI11_6/XI0/XI0_54/d__12_ DECAP_INV_G11
XG2679 XI11_6/XI0/XI0_54/d_11_ XI11_6/XI0/XI0_54/d__11_ DECAP_INV_G11
XG2680 XI11_6/XI0/XI0_54/d_10_ XI11_6/XI0/XI0_54/d__10_ DECAP_INV_G11
XG2681 XI11_6/XI0/XI0_54/d_9_ XI11_6/XI0/XI0_54/d__9_ DECAP_INV_G11
XG2682 XI11_6/XI0/XI0_54/d_8_ XI11_6/XI0/XI0_54/d__8_ DECAP_INV_G11
XG2683 XI11_6/XI0/XI0_54/d_7_ XI11_6/XI0/XI0_54/d__7_ DECAP_INV_G11
XG2684 XI11_6/XI0/XI0_54/d_6_ XI11_6/XI0/XI0_54/d__6_ DECAP_INV_G11
XG2685 XI11_6/XI0/XI0_54/d_5_ XI11_6/XI0/XI0_54/d__5_ DECAP_INV_G11
XG2686 XI11_6/XI0/XI0_54/d_4_ XI11_6/XI0/XI0_54/d__4_ DECAP_INV_G11
XG2687 XI11_6/XI0/XI0_54/d_3_ XI11_6/XI0/XI0_54/d__3_ DECAP_INV_G11
XG2688 XI11_6/XI0/XI0_54/d_2_ XI11_6/XI0/XI0_54/d__2_ DECAP_INV_G11
XG2689 XI11_6/XI0/XI0_54/d_1_ XI11_6/XI0/XI0_54/d__1_ DECAP_INV_G11
XG2690 XI11_6/XI0/XI0_54/d_0_ XI11_6/XI0/XI0_54/d__0_ DECAP_INV_G11
XG2691 XI11_6/XI0/XI0_53/d__15_ XI11_6/XI0/XI0_53/d_15_ DECAP_INV_G11
XG2692 XI11_6/XI0/XI0_53/d__14_ XI11_6/XI0/XI0_53/d_14_ DECAP_INV_G11
XG2693 XI11_6/XI0/XI0_53/d__13_ XI11_6/XI0/XI0_53/d_13_ DECAP_INV_G11
XG2694 XI11_6/XI0/XI0_53/d__12_ XI11_6/XI0/XI0_53/d_12_ DECAP_INV_G11
XG2695 XI11_6/XI0/XI0_53/d__11_ XI11_6/XI0/XI0_53/d_11_ DECAP_INV_G11
XG2696 XI11_6/XI0/XI0_53/d__10_ XI11_6/XI0/XI0_53/d_10_ DECAP_INV_G11
XG2697 XI11_6/XI0/XI0_53/d__9_ XI11_6/XI0/XI0_53/d_9_ DECAP_INV_G11
XG2698 XI11_6/XI0/XI0_53/d__8_ XI11_6/XI0/XI0_53/d_8_ DECAP_INV_G11
XG2699 XI11_6/XI0/XI0_53/d__7_ XI11_6/XI0/XI0_53/d_7_ DECAP_INV_G11
XG2700 XI11_6/XI0/XI0_53/d__6_ XI11_6/XI0/XI0_53/d_6_ DECAP_INV_G11
XG2701 XI11_6/XI0/XI0_53/d__5_ XI11_6/XI0/XI0_53/d_5_ DECAP_INV_G11
XG2702 XI11_6/XI0/XI0_53/d__4_ XI11_6/XI0/XI0_53/d_4_ DECAP_INV_G11
XG2703 XI11_6/XI0/XI0_53/d__3_ XI11_6/XI0/XI0_53/d_3_ DECAP_INV_G11
XG2704 XI11_6/XI0/XI0_53/d__2_ XI11_6/XI0/XI0_53/d_2_ DECAP_INV_G11
XG2705 XI11_6/XI0/XI0_53/d__1_ XI11_6/XI0/XI0_53/d_1_ DECAP_INV_G11
XG2706 XI11_6/XI0/XI0_53/d__0_ XI11_6/XI0/XI0_53/d_0_ DECAP_INV_G11
XG2707 XI11_6/XI0/XI0_53/d_15_ XI11_6/XI0/XI0_53/d__15_ DECAP_INV_G11
XG2708 XI11_6/XI0/XI0_53/d_14_ XI11_6/XI0/XI0_53/d__14_ DECAP_INV_G11
XG2709 XI11_6/XI0/XI0_53/d_13_ XI11_6/XI0/XI0_53/d__13_ DECAP_INV_G11
XG2710 XI11_6/XI0/XI0_53/d_12_ XI11_6/XI0/XI0_53/d__12_ DECAP_INV_G11
XG2711 XI11_6/XI0/XI0_53/d_11_ XI11_6/XI0/XI0_53/d__11_ DECAP_INV_G11
XG2712 XI11_6/XI0/XI0_53/d_10_ XI11_6/XI0/XI0_53/d__10_ DECAP_INV_G11
XG2713 XI11_6/XI0/XI0_53/d_9_ XI11_6/XI0/XI0_53/d__9_ DECAP_INV_G11
XG2714 XI11_6/XI0/XI0_53/d_8_ XI11_6/XI0/XI0_53/d__8_ DECAP_INV_G11
XG2715 XI11_6/XI0/XI0_53/d_7_ XI11_6/XI0/XI0_53/d__7_ DECAP_INV_G11
XG2716 XI11_6/XI0/XI0_53/d_6_ XI11_6/XI0/XI0_53/d__6_ DECAP_INV_G11
XG2717 XI11_6/XI0/XI0_53/d_5_ XI11_6/XI0/XI0_53/d__5_ DECAP_INV_G11
XG2718 XI11_6/XI0/XI0_53/d_4_ XI11_6/XI0/XI0_53/d__4_ DECAP_INV_G11
XG2719 XI11_6/XI0/XI0_53/d_3_ XI11_6/XI0/XI0_53/d__3_ DECAP_INV_G11
XG2720 XI11_6/XI0/XI0_53/d_2_ XI11_6/XI0/XI0_53/d__2_ DECAP_INV_G11
XG2721 XI11_6/XI0/XI0_53/d_1_ XI11_6/XI0/XI0_53/d__1_ DECAP_INV_G11
XG2722 XI11_6/XI0/XI0_53/d_0_ XI11_6/XI0/XI0_53/d__0_ DECAP_INV_G11
XG2723 XI11_6/XI0/XI0_52/d__15_ XI11_6/XI0/XI0_52/d_15_ DECAP_INV_G11
XG2724 XI11_6/XI0/XI0_52/d__14_ XI11_6/XI0/XI0_52/d_14_ DECAP_INV_G11
XG2725 XI11_6/XI0/XI0_52/d__13_ XI11_6/XI0/XI0_52/d_13_ DECAP_INV_G11
XG2726 XI11_6/XI0/XI0_52/d__12_ XI11_6/XI0/XI0_52/d_12_ DECAP_INV_G11
XG2727 XI11_6/XI0/XI0_52/d__11_ XI11_6/XI0/XI0_52/d_11_ DECAP_INV_G11
XG2728 XI11_6/XI0/XI0_52/d__10_ XI11_6/XI0/XI0_52/d_10_ DECAP_INV_G11
XG2729 XI11_6/XI0/XI0_52/d__9_ XI11_6/XI0/XI0_52/d_9_ DECAP_INV_G11
XG2730 XI11_6/XI0/XI0_52/d__8_ XI11_6/XI0/XI0_52/d_8_ DECAP_INV_G11
XG2731 XI11_6/XI0/XI0_52/d__7_ XI11_6/XI0/XI0_52/d_7_ DECAP_INV_G11
XG2732 XI11_6/XI0/XI0_52/d__6_ XI11_6/XI0/XI0_52/d_6_ DECAP_INV_G11
XG2733 XI11_6/XI0/XI0_52/d__5_ XI11_6/XI0/XI0_52/d_5_ DECAP_INV_G11
XG2734 XI11_6/XI0/XI0_52/d__4_ XI11_6/XI0/XI0_52/d_4_ DECAP_INV_G11
XG2735 XI11_6/XI0/XI0_52/d__3_ XI11_6/XI0/XI0_52/d_3_ DECAP_INV_G11
XG2736 XI11_6/XI0/XI0_52/d__2_ XI11_6/XI0/XI0_52/d_2_ DECAP_INV_G11
XG2737 XI11_6/XI0/XI0_52/d__1_ XI11_6/XI0/XI0_52/d_1_ DECAP_INV_G11
XG2738 XI11_6/XI0/XI0_52/d__0_ XI11_6/XI0/XI0_52/d_0_ DECAP_INV_G11
XG2739 XI11_6/XI0/XI0_52/d_15_ XI11_6/XI0/XI0_52/d__15_ DECAP_INV_G11
XG2740 XI11_6/XI0/XI0_52/d_14_ XI11_6/XI0/XI0_52/d__14_ DECAP_INV_G11
XG2741 XI11_6/XI0/XI0_52/d_13_ XI11_6/XI0/XI0_52/d__13_ DECAP_INV_G11
XG2742 XI11_6/XI0/XI0_52/d_12_ XI11_6/XI0/XI0_52/d__12_ DECAP_INV_G11
XG2743 XI11_6/XI0/XI0_52/d_11_ XI11_6/XI0/XI0_52/d__11_ DECAP_INV_G11
XG2744 XI11_6/XI0/XI0_52/d_10_ XI11_6/XI0/XI0_52/d__10_ DECAP_INV_G11
XG2745 XI11_6/XI0/XI0_52/d_9_ XI11_6/XI0/XI0_52/d__9_ DECAP_INV_G11
XG2746 XI11_6/XI0/XI0_52/d_8_ XI11_6/XI0/XI0_52/d__8_ DECAP_INV_G11
XG2747 XI11_6/XI0/XI0_52/d_7_ XI11_6/XI0/XI0_52/d__7_ DECAP_INV_G11
XG2748 XI11_6/XI0/XI0_52/d_6_ XI11_6/XI0/XI0_52/d__6_ DECAP_INV_G11
XG2749 XI11_6/XI0/XI0_52/d_5_ XI11_6/XI0/XI0_52/d__5_ DECAP_INV_G11
XG2750 XI11_6/XI0/XI0_52/d_4_ XI11_6/XI0/XI0_52/d__4_ DECAP_INV_G11
XG2751 XI11_6/XI0/XI0_52/d_3_ XI11_6/XI0/XI0_52/d__3_ DECAP_INV_G11
XG2752 XI11_6/XI0/XI0_52/d_2_ XI11_6/XI0/XI0_52/d__2_ DECAP_INV_G11
XG2753 XI11_6/XI0/XI0_52/d_1_ XI11_6/XI0/XI0_52/d__1_ DECAP_INV_G11
XG2754 XI11_6/XI0/XI0_52/d_0_ XI11_6/XI0/XI0_52/d__0_ DECAP_INV_G11
XG2755 XI11_6/XI0/XI0_51/d__15_ XI11_6/XI0/XI0_51/d_15_ DECAP_INV_G11
XG2756 XI11_6/XI0/XI0_51/d__14_ XI11_6/XI0/XI0_51/d_14_ DECAP_INV_G11
XG2757 XI11_6/XI0/XI0_51/d__13_ XI11_6/XI0/XI0_51/d_13_ DECAP_INV_G11
XG2758 XI11_6/XI0/XI0_51/d__12_ XI11_6/XI0/XI0_51/d_12_ DECAP_INV_G11
XG2759 XI11_6/XI0/XI0_51/d__11_ XI11_6/XI0/XI0_51/d_11_ DECAP_INV_G11
XG2760 XI11_6/XI0/XI0_51/d__10_ XI11_6/XI0/XI0_51/d_10_ DECAP_INV_G11
XG2761 XI11_6/XI0/XI0_51/d__9_ XI11_6/XI0/XI0_51/d_9_ DECAP_INV_G11
XG2762 XI11_6/XI0/XI0_51/d__8_ XI11_6/XI0/XI0_51/d_8_ DECAP_INV_G11
XG2763 XI11_6/XI0/XI0_51/d__7_ XI11_6/XI0/XI0_51/d_7_ DECAP_INV_G11
XG2764 XI11_6/XI0/XI0_51/d__6_ XI11_6/XI0/XI0_51/d_6_ DECAP_INV_G11
XG2765 XI11_6/XI0/XI0_51/d__5_ XI11_6/XI0/XI0_51/d_5_ DECAP_INV_G11
XG2766 XI11_6/XI0/XI0_51/d__4_ XI11_6/XI0/XI0_51/d_4_ DECAP_INV_G11
XG2767 XI11_6/XI0/XI0_51/d__3_ XI11_6/XI0/XI0_51/d_3_ DECAP_INV_G11
XG2768 XI11_6/XI0/XI0_51/d__2_ XI11_6/XI0/XI0_51/d_2_ DECAP_INV_G11
XG2769 XI11_6/XI0/XI0_51/d__1_ XI11_6/XI0/XI0_51/d_1_ DECAP_INV_G11
XG2770 XI11_6/XI0/XI0_51/d__0_ XI11_6/XI0/XI0_51/d_0_ DECAP_INV_G11
XG2771 XI11_6/XI0/XI0_51/d_15_ XI11_6/XI0/XI0_51/d__15_ DECAP_INV_G11
XG2772 XI11_6/XI0/XI0_51/d_14_ XI11_6/XI0/XI0_51/d__14_ DECAP_INV_G11
XG2773 XI11_6/XI0/XI0_51/d_13_ XI11_6/XI0/XI0_51/d__13_ DECAP_INV_G11
XG2774 XI11_6/XI0/XI0_51/d_12_ XI11_6/XI0/XI0_51/d__12_ DECAP_INV_G11
XG2775 XI11_6/XI0/XI0_51/d_11_ XI11_6/XI0/XI0_51/d__11_ DECAP_INV_G11
XG2776 XI11_6/XI0/XI0_51/d_10_ XI11_6/XI0/XI0_51/d__10_ DECAP_INV_G11
XG2777 XI11_6/XI0/XI0_51/d_9_ XI11_6/XI0/XI0_51/d__9_ DECAP_INV_G11
XG2778 XI11_6/XI0/XI0_51/d_8_ XI11_6/XI0/XI0_51/d__8_ DECAP_INV_G11
XG2779 XI11_6/XI0/XI0_51/d_7_ XI11_6/XI0/XI0_51/d__7_ DECAP_INV_G11
XG2780 XI11_6/XI0/XI0_51/d_6_ XI11_6/XI0/XI0_51/d__6_ DECAP_INV_G11
XG2781 XI11_6/XI0/XI0_51/d_5_ XI11_6/XI0/XI0_51/d__5_ DECAP_INV_G11
XG2782 XI11_6/XI0/XI0_51/d_4_ XI11_6/XI0/XI0_51/d__4_ DECAP_INV_G11
XG2783 XI11_6/XI0/XI0_51/d_3_ XI11_6/XI0/XI0_51/d__3_ DECAP_INV_G11
XG2784 XI11_6/XI0/XI0_51/d_2_ XI11_6/XI0/XI0_51/d__2_ DECAP_INV_G11
XG2785 XI11_6/XI0/XI0_51/d_1_ XI11_6/XI0/XI0_51/d__1_ DECAP_INV_G11
XG2786 XI11_6/XI0/XI0_51/d_0_ XI11_6/XI0/XI0_51/d__0_ DECAP_INV_G11
XG2787 XI11_6/XI0/XI0_50/d__15_ XI11_6/XI0/XI0_50/d_15_ DECAP_INV_G11
XG2788 XI11_6/XI0/XI0_50/d__14_ XI11_6/XI0/XI0_50/d_14_ DECAP_INV_G11
XG2789 XI11_6/XI0/XI0_50/d__13_ XI11_6/XI0/XI0_50/d_13_ DECAP_INV_G11
XG2790 XI11_6/XI0/XI0_50/d__12_ XI11_6/XI0/XI0_50/d_12_ DECAP_INV_G11
XG2791 XI11_6/XI0/XI0_50/d__11_ XI11_6/XI0/XI0_50/d_11_ DECAP_INV_G11
XG2792 XI11_6/XI0/XI0_50/d__10_ XI11_6/XI0/XI0_50/d_10_ DECAP_INV_G11
XG2793 XI11_6/XI0/XI0_50/d__9_ XI11_6/XI0/XI0_50/d_9_ DECAP_INV_G11
XG2794 XI11_6/XI0/XI0_50/d__8_ XI11_6/XI0/XI0_50/d_8_ DECAP_INV_G11
XG2795 XI11_6/XI0/XI0_50/d__7_ XI11_6/XI0/XI0_50/d_7_ DECAP_INV_G11
XG2796 XI11_6/XI0/XI0_50/d__6_ XI11_6/XI0/XI0_50/d_6_ DECAP_INV_G11
XG2797 XI11_6/XI0/XI0_50/d__5_ XI11_6/XI0/XI0_50/d_5_ DECAP_INV_G11
XG2798 XI11_6/XI0/XI0_50/d__4_ XI11_6/XI0/XI0_50/d_4_ DECAP_INV_G11
XG2799 XI11_6/XI0/XI0_50/d__3_ XI11_6/XI0/XI0_50/d_3_ DECAP_INV_G11
XG2800 XI11_6/XI0/XI0_50/d__2_ XI11_6/XI0/XI0_50/d_2_ DECAP_INV_G11
XG2801 XI11_6/XI0/XI0_50/d__1_ XI11_6/XI0/XI0_50/d_1_ DECAP_INV_G11
XG2802 XI11_6/XI0/XI0_50/d__0_ XI11_6/XI0/XI0_50/d_0_ DECAP_INV_G11
XG2803 XI11_6/XI0/XI0_50/d_15_ XI11_6/XI0/XI0_50/d__15_ DECAP_INV_G11
XG2804 XI11_6/XI0/XI0_50/d_14_ XI11_6/XI0/XI0_50/d__14_ DECAP_INV_G11
XG2805 XI11_6/XI0/XI0_50/d_13_ XI11_6/XI0/XI0_50/d__13_ DECAP_INV_G11
XG2806 XI11_6/XI0/XI0_50/d_12_ XI11_6/XI0/XI0_50/d__12_ DECAP_INV_G11
XG2807 XI11_6/XI0/XI0_50/d_11_ XI11_6/XI0/XI0_50/d__11_ DECAP_INV_G11
XG2808 XI11_6/XI0/XI0_50/d_10_ XI11_6/XI0/XI0_50/d__10_ DECAP_INV_G11
XG2809 XI11_6/XI0/XI0_50/d_9_ XI11_6/XI0/XI0_50/d__9_ DECAP_INV_G11
XG2810 XI11_6/XI0/XI0_50/d_8_ XI11_6/XI0/XI0_50/d__8_ DECAP_INV_G11
XG2811 XI11_6/XI0/XI0_50/d_7_ XI11_6/XI0/XI0_50/d__7_ DECAP_INV_G11
XG2812 XI11_6/XI0/XI0_50/d_6_ XI11_6/XI0/XI0_50/d__6_ DECAP_INV_G11
XG2813 XI11_6/XI0/XI0_50/d_5_ XI11_6/XI0/XI0_50/d__5_ DECAP_INV_G11
XG2814 XI11_6/XI0/XI0_50/d_4_ XI11_6/XI0/XI0_50/d__4_ DECAP_INV_G11
XG2815 XI11_6/XI0/XI0_50/d_3_ XI11_6/XI0/XI0_50/d__3_ DECAP_INV_G11
XG2816 XI11_6/XI0/XI0_50/d_2_ XI11_6/XI0/XI0_50/d__2_ DECAP_INV_G11
XG2817 XI11_6/XI0/XI0_50/d_1_ XI11_6/XI0/XI0_50/d__1_ DECAP_INV_G11
XG2818 XI11_6/XI0/XI0_50/d_0_ XI11_6/XI0/XI0_50/d__0_ DECAP_INV_G11
XG2819 XI11_6/XI0/XI0_49/d__15_ XI11_6/XI0/XI0_49/d_15_ DECAP_INV_G11
XG2820 XI11_6/XI0/XI0_49/d__14_ XI11_6/XI0/XI0_49/d_14_ DECAP_INV_G11
XG2821 XI11_6/XI0/XI0_49/d__13_ XI11_6/XI0/XI0_49/d_13_ DECAP_INV_G11
XG2822 XI11_6/XI0/XI0_49/d__12_ XI11_6/XI0/XI0_49/d_12_ DECAP_INV_G11
XG2823 XI11_6/XI0/XI0_49/d__11_ XI11_6/XI0/XI0_49/d_11_ DECAP_INV_G11
XG2824 XI11_6/XI0/XI0_49/d__10_ XI11_6/XI0/XI0_49/d_10_ DECAP_INV_G11
XG2825 XI11_6/XI0/XI0_49/d__9_ XI11_6/XI0/XI0_49/d_9_ DECAP_INV_G11
XG2826 XI11_6/XI0/XI0_49/d__8_ XI11_6/XI0/XI0_49/d_8_ DECAP_INV_G11
XG2827 XI11_6/XI0/XI0_49/d__7_ XI11_6/XI0/XI0_49/d_7_ DECAP_INV_G11
XG2828 XI11_6/XI0/XI0_49/d__6_ XI11_6/XI0/XI0_49/d_6_ DECAP_INV_G11
XG2829 XI11_6/XI0/XI0_49/d__5_ XI11_6/XI0/XI0_49/d_5_ DECAP_INV_G11
XG2830 XI11_6/XI0/XI0_49/d__4_ XI11_6/XI0/XI0_49/d_4_ DECAP_INV_G11
XG2831 XI11_6/XI0/XI0_49/d__3_ XI11_6/XI0/XI0_49/d_3_ DECAP_INV_G11
XG2832 XI11_6/XI0/XI0_49/d__2_ XI11_6/XI0/XI0_49/d_2_ DECAP_INV_G11
XG2833 XI11_6/XI0/XI0_49/d__1_ XI11_6/XI0/XI0_49/d_1_ DECAP_INV_G11
XG2834 XI11_6/XI0/XI0_49/d__0_ XI11_6/XI0/XI0_49/d_0_ DECAP_INV_G11
XG2835 XI11_6/XI0/XI0_49/d_15_ XI11_6/XI0/XI0_49/d__15_ DECAP_INV_G11
XG2836 XI11_6/XI0/XI0_49/d_14_ XI11_6/XI0/XI0_49/d__14_ DECAP_INV_G11
XG2837 XI11_6/XI0/XI0_49/d_13_ XI11_6/XI0/XI0_49/d__13_ DECAP_INV_G11
XG2838 XI11_6/XI0/XI0_49/d_12_ XI11_6/XI0/XI0_49/d__12_ DECAP_INV_G11
XG2839 XI11_6/XI0/XI0_49/d_11_ XI11_6/XI0/XI0_49/d__11_ DECAP_INV_G11
XG2840 XI11_6/XI0/XI0_49/d_10_ XI11_6/XI0/XI0_49/d__10_ DECAP_INV_G11
XG2841 XI11_6/XI0/XI0_49/d_9_ XI11_6/XI0/XI0_49/d__9_ DECAP_INV_G11
XG2842 XI11_6/XI0/XI0_49/d_8_ XI11_6/XI0/XI0_49/d__8_ DECAP_INV_G11
XG2843 XI11_6/XI0/XI0_49/d_7_ XI11_6/XI0/XI0_49/d__7_ DECAP_INV_G11
XG2844 XI11_6/XI0/XI0_49/d_6_ XI11_6/XI0/XI0_49/d__6_ DECAP_INV_G11
XG2845 XI11_6/XI0/XI0_49/d_5_ XI11_6/XI0/XI0_49/d__5_ DECAP_INV_G11
XG2846 XI11_6/XI0/XI0_49/d_4_ XI11_6/XI0/XI0_49/d__4_ DECAP_INV_G11
XG2847 XI11_6/XI0/XI0_49/d_3_ XI11_6/XI0/XI0_49/d__3_ DECAP_INV_G11
XG2848 XI11_6/XI0/XI0_49/d_2_ XI11_6/XI0/XI0_49/d__2_ DECAP_INV_G11
XG2849 XI11_6/XI0/XI0_49/d_1_ XI11_6/XI0/XI0_49/d__1_ DECAP_INV_G11
XG2850 XI11_6/XI0/XI0_49/d_0_ XI11_6/XI0/XI0_49/d__0_ DECAP_INV_G11
XG2851 XI11_6/XI0/XI0_48/d__15_ XI11_6/XI0/XI0_48/d_15_ DECAP_INV_G11
XG2852 XI11_6/XI0/XI0_48/d__14_ XI11_6/XI0/XI0_48/d_14_ DECAP_INV_G11
XG2853 XI11_6/XI0/XI0_48/d__13_ XI11_6/XI0/XI0_48/d_13_ DECAP_INV_G11
XG2854 XI11_6/XI0/XI0_48/d__12_ XI11_6/XI0/XI0_48/d_12_ DECAP_INV_G11
XG2855 XI11_6/XI0/XI0_48/d__11_ XI11_6/XI0/XI0_48/d_11_ DECAP_INV_G11
XG2856 XI11_6/XI0/XI0_48/d__10_ XI11_6/XI0/XI0_48/d_10_ DECAP_INV_G11
XG2857 XI11_6/XI0/XI0_48/d__9_ XI11_6/XI0/XI0_48/d_9_ DECAP_INV_G11
XG2858 XI11_6/XI0/XI0_48/d__8_ XI11_6/XI0/XI0_48/d_8_ DECAP_INV_G11
XG2859 XI11_6/XI0/XI0_48/d__7_ XI11_6/XI0/XI0_48/d_7_ DECAP_INV_G11
XG2860 XI11_6/XI0/XI0_48/d__6_ XI11_6/XI0/XI0_48/d_6_ DECAP_INV_G11
XG2861 XI11_6/XI0/XI0_48/d__5_ XI11_6/XI0/XI0_48/d_5_ DECAP_INV_G11
XG2862 XI11_6/XI0/XI0_48/d__4_ XI11_6/XI0/XI0_48/d_4_ DECAP_INV_G11
XG2863 XI11_6/XI0/XI0_48/d__3_ XI11_6/XI0/XI0_48/d_3_ DECAP_INV_G11
XG2864 XI11_6/XI0/XI0_48/d__2_ XI11_6/XI0/XI0_48/d_2_ DECAP_INV_G11
XG2865 XI11_6/XI0/XI0_48/d__1_ XI11_6/XI0/XI0_48/d_1_ DECAP_INV_G11
XG2866 XI11_6/XI0/XI0_48/d__0_ XI11_6/XI0/XI0_48/d_0_ DECAP_INV_G11
XG2867 XI11_6/XI0/XI0_48/d_15_ XI11_6/XI0/XI0_48/d__15_ DECAP_INV_G11
XG2868 XI11_6/XI0/XI0_48/d_14_ XI11_6/XI0/XI0_48/d__14_ DECAP_INV_G11
XG2869 XI11_6/XI0/XI0_48/d_13_ XI11_6/XI0/XI0_48/d__13_ DECAP_INV_G11
XG2870 XI11_6/XI0/XI0_48/d_12_ XI11_6/XI0/XI0_48/d__12_ DECAP_INV_G11
XG2871 XI11_6/XI0/XI0_48/d_11_ XI11_6/XI0/XI0_48/d__11_ DECAP_INV_G11
XG2872 XI11_6/XI0/XI0_48/d_10_ XI11_6/XI0/XI0_48/d__10_ DECAP_INV_G11
XG2873 XI11_6/XI0/XI0_48/d_9_ XI11_6/XI0/XI0_48/d__9_ DECAP_INV_G11
XG2874 XI11_6/XI0/XI0_48/d_8_ XI11_6/XI0/XI0_48/d__8_ DECAP_INV_G11
XG2875 XI11_6/XI0/XI0_48/d_7_ XI11_6/XI0/XI0_48/d__7_ DECAP_INV_G11
XG2876 XI11_6/XI0/XI0_48/d_6_ XI11_6/XI0/XI0_48/d__6_ DECAP_INV_G11
XG2877 XI11_6/XI0/XI0_48/d_5_ XI11_6/XI0/XI0_48/d__5_ DECAP_INV_G11
XG2878 XI11_6/XI0/XI0_48/d_4_ XI11_6/XI0/XI0_48/d__4_ DECAP_INV_G11
XG2879 XI11_6/XI0/XI0_48/d_3_ XI11_6/XI0/XI0_48/d__3_ DECAP_INV_G11
XG2880 XI11_6/XI0/XI0_48/d_2_ XI11_6/XI0/XI0_48/d__2_ DECAP_INV_G11
XG2881 XI11_6/XI0/XI0_48/d_1_ XI11_6/XI0/XI0_48/d__1_ DECAP_INV_G11
XG2882 XI11_6/XI0/XI0_48/d_0_ XI11_6/XI0/XI0_48/d__0_ DECAP_INV_G11
XG2883 XI11_6/XI0/XI0_47/d__15_ XI11_6/XI0/XI0_47/d_15_ DECAP_INV_G11
XG2884 XI11_6/XI0/XI0_47/d__14_ XI11_6/XI0/XI0_47/d_14_ DECAP_INV_G11
XG2885 XI11_6/XI0/XI0_47/d__13_ XI11_6/XI0/XI0_47/d_13_ DECAP_INV_G11
XG2886 XI11_6/XI0/XI0_47/d__12_ XI11_6/XI0/XI0_47/d_12_ DECAP_INV_G11
XG2887 XI11_6/XI0/XI0_47/d__11_ XI11_6/XI0/XI0_47/d_11_ DECAP_INV_G11
XG2888 XI11_6/XI0/XI0_47/d__10_ XI11_6/XI0/XI0_47/d_10_ DECAP_INV_G11
XG2889 XI11_6/XI0/XI0_47/d__9_ XI11_6/XI0/XI0_47/d_9_ DECAP_INV_G11
XG2890 XI11_6/XI0/XI0_47/d__8_ XI11_6/XI0/XI0_47/d_8_ DECAP_INV_G11
XG2891 XI11_6/XI0/XI0_47/d__7_ XI11_6/XI0/XI0_47/d_7_ DECAP_INV_G11
XG2892 XI11_6/XI0/XI0_47/d__6_ XI11_6/XI0/XI0_47/d_6_ DECAP_INV_G11
XG2893 XI11_6/XI0/XI0_47/d__5_ XI11_6/XI0/XI0_47/d_5_ DECAP_INV_G11
XG2894 XI11_6/XI0/XI0_47/d__4_ XI11_6/XI0/XI0_47/d_4_ DECAP_INV_G11
XG2895 XI11_6/XI0/XI0_47/d__3_ XI11_6/XI0/XI0_47/d_3_ DECAP_INV_G11
XG2896 XI11_6/XI0/XI0_47/d__2_ XI11_6/XI0/XI0_47/d_2_ DECAP_INV_G11
XG2897 XI11_6/XI0/XI0_47/d__1_ XI11_6/XI0/XI0_47/d_1_ DECAP_INV_G11
XG2898 XI11_6/XI0/XI0_47/d__0_ XI11_6/XI0/XI0_47/d_0_ DECAP_INV_G11
XG2899 XI11_6/XI0/XI0_47/d_15_ XI11_6/XI0/XI0_47/d__15_ DECAP_INV_G11
XG2900 XI11_6/XI0/XI0_47/d_14_ XI11_6/XI0/XI0_47/d__14_ DECAP_INV_G11
XG2901 XI11_6/XI0/XI0_47/d_13_ XI11_6/XI0/XI0_47/d__13_ DECAP_INV_G11
XG2902 XI11_6/XI0/XI0_47/d_12_ XI11_6/XI0/XI0_47/d__12_ DECAP_INV_G11
XG2903 XI11_6/XI0/XI0_47/d_11_ XI11_6/XI0/XI0_47/d__11_ DECAP_INV_G11
XG2904 XI11_6/XI0/XI0_47/d_10_ XI11_6/XI0/XI0_47/d__10_ DECAP_INV_G11
XG2905 XI11_6/XI0/XI0_47/d_9_ XI11_6/XI0/XI0_47/d__9_ DECAP_INV_G11
XG2906 XI11_6/XI0/XI0_47/d_8_ XI11_6/XI0/XI0_47/d__8_ DECAP_INV_G11
XG2907 XI11_6/XI0/XI0_47/d_7_ XI11_6/XI0/XI0_47/d__7_ DECAP_INV_G11
XG2908 XI11_6/XI0/XI0_47/d_6_ XI11_6/XI0/XI0_47/d__6_ DECAP_INV_G11
XG2909 XI11_6/XI0/XI0_47/d_5_ XI11_6/XI0/XI0_47/d__5_ DECAP_INV_G11
XG2910 XI11_6/XI0/XI0_47/d_4_ XI11_6/XI0/XI0_47/d__4_ DECAP_INV_G11
XG2911 XI11_6/XI0/XI0_47/d_3_ XI11_6/XI0/XI0_47/d__3_ DECAP_INV_G11
XG2912 XI11_6/XI0/XI0_47/d_2_ XI11_6/XI0/XI0_47/d__2_ DECAP_INV_G11
XG2913 XI11_6/XI0/XI0_47/d_1_ XI11_6/XI0/XI0_47/d__1_ DECAP_INV_G11
XG2914 XI11_6/XI0/XI0_47/d_0_ XI11_6/XI0/XI0_47/d__0_ DECAP_INV_G11
XG2915 XI11_6/XI0/XI0_46/d__15_ XI11_6/XI0/XI0_46/d_15_ DECAP_INV_G11
XG2916 XI11_6/XI0/XI0_46/d__14_ XI11_6/XI0/XI0_46/d_14_ DECAP_INV_G11
XG2917 XI11_6/XI0/XI0_46/d__13_ XI11_6/XI0/XI0_46/d_13_ DECAP_INV_G11
XG2918 XI11_6/XI0/XI0_46/d__12_ XI11_6/XI0/XI0_46/d_12_ DECAP_INV_G11
XG2919 XI11_6/XI0/XI0_46/d__11_ XI11_6/XI0/XI0_46/d_11_ DECAP_INV_G11
XG2920 XI11_6/XI0/XI0_46/d__10_ XI11_6/XI0/XI0_46/d_10_ DECAP_INV_G11
XG2921 XI11_6/XI0/XI0_46/d__9_ XI11_6/XI0/XI0_46/d_9_ DECAP_INV_G11
XG2922 XI11_6/XI0/XI0_46/d__8_ XI11_6/XI0/XI0_46/d_8_ DECAP_INV_G11
XG2923 XI11_6/XI0/XI0_46/d__7_ XI11_6/XI0/XI0_46/d_7_ DECAP_INV_G11
XG2924 XI11_6/XI0/XI0_46/d__6_ XI11_6/XI0/XI0_46/d_6_ DECAP_INV_G11
XG2925 XI11_6/XI0/XI0_46/d__5_ XI11_6/XI0/XI0_46/d_5_ DECAP_INV_G11
XG2926 XI11_6/XI0/XI0_46/d__4_ XI11_6/XI0/XI0_46/d_4_ DECAP_INV_G11
XG2927 XI11_6/XI0/XI0_46/d__3_ XI11_6/XI0/XI0_46/d_3_ DECAP_INV_G11
XG2928 XI11_6/XI0/XI0_46/d__2_ XI11_6/XI0/XI0_46/d_2_ DECAP_INV_G11
XG2929 XI11_6/XI0/XI0_46/d__1_ XI11_6/XI0/XI0_46/d_1_ DECAP_INV_G11
XG2930 XI11_6/XI0/XI0_46/d__0_ XI11_6/XI0/XI0_46/d_0_ DECAP_INV_G11
XG2931 XI11_6/XI0/XI0_46/d_15_ XI11_6/XI0/XI0_46/d__15_ DECAP_INV_G11
XG2932 XI11_6/XI0/XI0_46/d_14_ XI11_6/XI0/XI0_46/d__14_ DECAP_INV_G11
XG2933 XI11_6/XI0/XI0_46/d_13_ XI11_6/XI0/XI0_46/d__13_ DECAP_INV_G11
XG2934 XI11_6/XI0/XI0_46/d_12_ XI11_6/XI0/XI0_46/d__12_ DECAP_INV_G11
XG2935 XI11_6/XI0/XI0_46/d_11_ XI11_6/XI0/XI0_46/d__11_ DECAP_INV_G11
XG2936 XI11_6/XI0/XI0_46/d_10_ XI11_6/XI0/XI0_46/d__10_ DECAP_INV_G11
XG2937 XI11_6/XI0/XI0_46/d_9_ XI11_6/XI0/XI0_46/d__9_ DECAP_INV_G11
XG2938 XI11_6/XI0/XI0_46/d_8_ XI11_6/XI0/XI0_46/d__8_ DECAP_INV_G11
XG2939 XI11_6/XI0/XI0_46/d_7_ XI11_6/XI0/XI0_46/d__7_ DECAP_INV_G11
XG2940 XI11_6/XI0/XI0_46/d_6_ XI11_6/XI0/XI0_46/d__6_ DECAP_INV_G11
XG2941 XI11_6/XI0/XI0_46/d_5_ XI11_6/XI0/XI0_46/d__5_ DECAP_INV_G11
XG2942 XI11_6/XI0/XI0_46/d_4_ XI11_6/XI0/XI0_46/d__4_ DECAP_INV_G11
XG2943 XI11_6/XI0/XI0_46/d_3_ XI11_6/XI0/XI0_46/d__3_ DECAP_INV_G11
XG2944 XI11_6/XI0/XI0_46/d_2_ XI11_6/XI0/XI0_46/d__2_ DECAP_INV_G11
XG2945 XI11_6/XI0/XI0_46/d_1_ XI11_6/XI0/XI0_46/d__1_ DECAP_INV_G11
XG2946 XI11_6/XI0/XI0_46/d_0_ XI11_6/XI0/XI0_46/d__0_ DECAP_INV_G11
XG2947 XI11_6/XI0/XI0_45/d__15_ XI11_6/XI0/XI0_45/d_15_ DECAP_INV_G11
XG2948 XI11_6/XI0/XI0_45/d__14_ XI11_6/XI0/XI0_45/d_14_ DECAP_INV_G11
XG2949 XI11_6/XI0/XI0_45/d__13_ XI11_6/XI0/XI0_45/d_13_ DECAP_INV_G11
XG2950 XI11_6/XI0/XI0_45/d__12_ XI11_6/XI0/XI0_45/d_12_ DECAP_INV_G11
XG2951 XI11_6/XI0/XI0_45/d__11_ XI11_6/XI0/XI0_45/d_11_ DECAP_INV_G11
XG2952 XI11_6/XI0/XI0_45/d__10_ XI11_6/XI0/XI0_45/d_10_ DECAP_INV_G11
XG2953 XI11_6/XI0/XI0_45/d__9_ XI11_6/XI0/XI0_45/d_9_ DECAP_INV_G11
XG2954 XI11_6/XI0/XI0_45/d__8_ XI11_6/XI0/XI0_45/d_8_ DECAP_INV_G11
XG2955 XI11_6/XI0/XI0_45/d__7_ XI11_6/XI0/XI0_45/d_7_ DECAP_INV_G11
XG2956 XI11_6/XI0/XI0_45/d__6_ XI11_6/XI0/XI0_45/d_6_ DECAP_INV_G11
XG2957 XI11_6/XI0/XI0_45/d__5_ XI11_6/XI0/XI0_45/d_5_ DECAP_INV_G11
XG2958 XI11_6/XI0/XI0_45/d__4_ XI11_6/XI0/XI0_45/d_4_ DECAP_INV_G11
XG2959 XI11_6/XI0/XI0_45/d__3_ XI11_6/XI0/XI0_45/d_3_ DECAP_INV_G11
XG2960 XI11_6/XI0/XI0_45/d__2_ XI11_6/XI0/XI0_45/d_2_ DECAP_INV_G11
XG2961 XI11_6/XI0/XI0_45/d__1_ XI11_6/XI0/XI0_45/d_1_ DECAP_INV_G11
XG2962 XI11_6/XI0/XI0_45/d__0_ XI11_6/XI0/XI0_45/d_0_ DECAP_INV_G11
XG2963 XI11_6/XI0/XI0_45/d_15_ XI11_6/XI0/XI0_45/d__15_ DECAP_INV_G11
XG2964 XI11_6/XI0/XI0_45/d_14_ XI11_6/XI0/XI0_45/d__14_ DECAP_INV_G11
XG2965 XI11_6/XI0/XI0_45/d_13_ XI11_6/XI0/XI0_45/d__13_ DECAP_INV_G11
XG2966 XI11_6/XI0/XI0_45/d_12_ XI11_6/XI0/XI0_45/d__12_ DECAP_INV_G11
XG2967 XI11_6/XI0/XI0_45/d_11_ XI11_6/XI0/XI0_45/d__11_ DECAP_INV_G11
XG2968 XI11_6/XI0/XI0_45/d_10_ XI11_6/XI0/XI0_45/d__10_ DECAP_INV_G11
XG2969 XI11_6/XI0/XI0_45/d_9_ XI11_6/XI0/XI0_45/d__9_ DECAP_INV_G11
XG2970 XI11_6/XI0/XI0_45/d_8_ XI11_6/XI0/XI0_45/d__8_ DECAP_INV_G11
XG2971 XI11_6/XI0/XI0_45/d_7_ XI11_6/XI0/XI0_45/d__7_ DECAP_INV_G11
XG2972 XI11_6/XI0/XI0_45/d_6_ XI11_6/XI0/XI0_45/d__6_ DECAP_INV_G11
XG2973 XI11_6/XI0/XI0_45/d_5_ XI11_6/XI0/XI0_45/d__5_ DECAP_INV_G11
XG2974 XI11_6/XI0/XI0_45/d_4_ XI11_6/XI0/XI0_45/d__4_ DECAP_INV_G11
XG2975 XI11_6/XI0/XI0_45/d_3_ XI11_6/XI0/XI0_45/d__3_ DECAP_INV_G11
XG2976 XI11_6/XI0/XI0_45/d_2_ XI11_6/XI0/XI0_45/d__2_ DECAP_INV_G11
XG2977 XI11_6/XI0/XI0_45/d_1_ XI11_6/XI0/XI0_45/d__1_ DECAP_INV_G11
XG2978 XI11_6/XI0/XI0_45/d_0_ XI11_6/XI0/XI0_45/d__0_ DECAP_INV_G11
XG2979 XI11_6/XI0/XI0_44/d__15_ XI11_6/XI0/XI0_44/d_15_ DECAP_INV_G11
XG2980 XI11_6/XI0/XI0_44/d__14_ XI11_6/XI0/XI0_44/d_14_ DECAP_INV_G11
XG2981 XI11_6/XI0/XI0_44/d__13_ XI11_6/XI0/XI0_44/d_13_ DECAP_INV_G11
XG2982 XI11_6/XI0/XI0_44/d__12_ XI11_6/XI0/XI0_44/d_12_ DECAP_INV_G11
XG2983 XI11_6/XI0/XI0_44/d__11_ XI11_6/XI0/XI0_44/d_11_ DECAP_INV_G11
XG2984 XI11_6/XI0/XI0_44/d__10_ XI11_6/XI0/XI0_44/d_10_ DECAP_INV_G11
XG2985 XI11_6/XI0/XI0_44/d__9_ XI11_6/XI0/XI0_44/d_9_ DECAP_INV_G11
XG2986 XI11_6/XI0/XI0_44/d__8_ XI11_6/XI0/XI0_44/d_8_ DECAP_INV_G11
XG2987 XI11_6/XI0/XI0_44/d__7_ XI11_6/XI0/XI0_44/d_7_ DECAP_INV_G11
XG2988 XI11_6/XI0/XI0_44/d__6_ XI11_6/XI0/XI0_44/d_6_ DECAP_INV_G11
XG2989 XI11_6/XI0/XI0_44/d__5_ XI11_6/XI0/XI0_44/d_5_ DECAP_INV_G11
XG2990 XI11_6/XI0/XI0_44/d__4_ XI11_6/XI0/XI0_44/d_4_ DECAP_INV_G11
XG2991 XI11_6/XI0/XI0_44/d__3_ XI11_6/XI0/XI0_44/d_3_ DECAP_INV_G11
XG2992 XI11_6/XI0/XI0_44/d__2_ XI11_6/XI0/XI0_44/d_2_ DECAP_INV_G11
XG2993 XI11_6/XI0/XI0_44/d__1_ XI11_6/XI0/XI0_44/d_1_ DECAP_INV_G11
XG2994 XI11_6/XI0/XI0_44/d__0_ XI11_6/XI0/XI0_44/d_0_ DECAP_INV_G11
XG2995 XI11_6/XI0/XI0_44/d_15_ XI11_6/XI0/XI0_44/d__15_ DECAP_INV_G11
XG2996 XI11_6/XI0/XI0_44/d_14_ XI11_6/XI0/XI0_44/d__14_ DECAP_INV_G11
XG2997 XI11_6/XI0/XI0_44/d_13_ XI11_6/XI0/XI0_44/d__13_ DECAP_INV_G11
XG2998 XI11_6/XI0/XI0_44/d_12_ XI11_6/XI0/XI0_44/d__12_ DECAP_INV_G11
XG2999 XI11_6/XI0/XI0_44/d_11_ XI11_6/XI0/XI0_44/d__11_ DECAP_INV_G11
XG3000 XI11_6/XI0/XI0_44/d_10_ XI11_6/XI0/XI0_44/d__10_ DECAP_INV_G11
XG3001 XI11_6/XI0/XI0_44/d_9_ XI11_6/XI0/XI0_44/d__9_ DECAP_INV_G11
XG3002 XI11_6/XI0/XI0_44/d_8_ XI11_6/XI0/XI0_44/d__8_ DECAP_INV_G11
XG3003 XI11_6/XI0/XI0_44/d_7_ XI11_6/XI0/XI0_44/d__7_ DECAP_INV_G11
XG3004 XI11_6/XI0/XI0_44/d_6_ XI11_6/XI0/XI0_44/d__6_ DECAP_INV_G11
XG3005 XI11_6/XI0/XI0_44/d_5_ XI11_6/XI0/XI0_44/d__5_ DECAP_INV_G11
XG3006 XI11_6/XI0/XI0_44/d_4_ XI11_6/XI0/XI0_44/d__4_ DECAP_INV_G11
XG3007 XI11_6/XI0/XI0_44/d_3_ XI11_6/XI0/XI0_44/d__3_ DECAP_INV_G11
XG3008 XI11_6/XI0/XI0_44/d_2_ XI11_6/XI0/XI0_44/d__2_ DECAP_INV_G11
XG3009 XI11_6/XI0/XI0_44/d_1_ XI11_6/XI0/XI0_44/d__1_ DECAP_INV_G11
XG3010 XI11_6/XI0/XI0_44/d_0_ XI11_6/XI0/XI0_44/d__0_ DECAP_INV_G11
XG3011 XI11_6/XI0/XI0_43/d__15_ XI11_6/XI0/XI0_43/d_15_ DECAP_INV_G11
XG3012 XI11_6/XI0/XI0_43/d__14_ XI11_6/XI0/XI0_43/d_14_ DECAP_INV_G11
XG3013 XI11_6/XI0/XI0_43/d__13_ XI11_6/XI0/XI0_43/d_13_ DECAP_INV_G11
XG3014 XI11_6/XI0/XI0_43/d__12_ XI11_6/XI0/XI0_43/d_12_ DECAP_INV_G11
XG3015 XI11_6/XI0/XI0_43/d__11_ XI11_6/XI0/XI0_43/d_11_ DECAP_INV_G11
XG3016 XI11_6/XI0/XI0_43/d__10_ XI11_6/XI0/XI0_43/d_10_ DECAP_INV_G11
XG3017 XI11_6/XI0/XI0_43/d__9_ XI11_6/XI0/XI0_43/d_9_ DECAP_INV_G11
XG3018 XI11_6/XI0/XI0_43/d__8_ XI11_6/XI0/XI0_43/d_8_ DECAP_INV_G11
XG3019 XI11_6/XI0/XI0_43/d__7_ XI11_6/XI0/XI0_43/d_7_ DECAP_INV_G11
XG3020 XI11_6/XI0/XI0_43/d__6_ XI11_6/XI0/XI0_43/d_6_ DECAP_INV_G11
XG3021 XI11_6/XI0/XI0_43/d__5_ XI11_6/XI0/XI0_43/d_5_ DECAP_INV_G11
XG3022 XI11_6/XI0/XI0_43/d__4_ XI11_6/XI0/XI0_43/d_4_ DECAP_INV_G11
XG3023 XI11_6/XI0/XI0_43/d__3_ XI11_6/XI0/XI0_43/d_3_ DECAP_INV_G11
XG3024 XI11_6/XI0/XI0_43/d__2_ XI11_6/XI0/XI0_43/d_2_ DECAP_INV_G11
XG3025 XI11_6/XI0/XI0_43/d__1_ XI11_6/XI0/XI0_43/d_1_ DECAP_INV_G11
XG3026 XI11_6/XI0/XI0_43/d__0_ XI11_6/XI0/XI0_43/d_0_ DECAP_INV_G11
XG3027 XI11_6/XI0/XI0_43/d_15_ XI11_6/XI0/XI0_43/d__15_ DECAP_INV_G11
XG3028 XI11_6/XI0/XI0_43/d_14_ XI11_6/XI0/XI0_43/d__14_ DECAP_INV_G11
XG3029 XI11_6/XI0/XI0_43/d_13_ XI11_6/XI0/XI0_43/d__13_ DECAP_INV_G11
XG3030 XI11_6/XI0/XI0_43/d_12_ XI11_6/XI0/XI0_43/d__12_ DECAP_INV_G11
XG3031 XI11_6/XI0/XI0_43/d_11_ XI11_6/XI0/XI0_43/d__11_ DECAP_INV_G11
XG3032 XI11_6/XI0/XI0_43/d_10_ XI11_6/XI0/XI0_43/d__10_ DECAP_INV_G11
XG3033 XI11_6/XI0/XI0_43/d_9_ XI11_6/XI0/XI0_43/d__9_ DECAP_INV_G11
XG3034 XI11_6/XI0/XI0_43/d_8_ XI11_6/XI0/XI0_43/d__8_ DECAP_INV_G11
XG3035 XI11_6/XI0/XI0_43/d_7_ XI11_6/XI0/XI0_43/d__7_ DECAP_INV_G11
XG3036 XI11_6/XI0/XI0_43/d_6_ XI11_6/XI0/XI0_43/d__6_ DECAP_INV_G11
XG3037 XI11_6/XI0/XI0_43/d_5_ XI11_6/XI0/XI0_43/d__5_ DECAP_INV_G11
XG3038 XI11_6/XI0/XI0_43/d_4_ XI11_6/XI0/XI0_43/d__4_ DECAP_INV_G11
XG3039 XI11_6/XI0/XI0_43/d_3_ XI11_6/XI0/XI0_43/d__3_ DECAP_INV_G11
XG3040 XI11_6/XI0/XI0_43/d_2_ XI11_6/XI0/XI0_43/d__2_ DECAP_INV_G11
XG3041 XI11_6/XI0/XI0_43/d_1_ XI11_6/XI0/XI0_43/d__1_ DECAP_INV_G11
XG3042 XI11_6/XI0/XI0_43/d_0_ XI11_6/XI0/XI0_43/d__0_ DECAP_INV_G11
XG3043 XI11_6/XI0/XI0_42/d__15_ XI11_6/XI0/XI0_42/d_15_ DECAP_INV_G11
XG3044 XI11_6/XI0/XI0_42/d__14_ XI11_6/XI0/XI0_42/d_14_ DECAP_INV_G11
XG3045 XI11_6/XI0/XI0_42/d__13_ XI11_6/XI0/XI0_42/d_13_ DECAP_INV_G11
XG3046 XI11_6/XI0/XI0_42/d__12_ XI11_6/XI0/XI0_42/d_12_ DECAP_INV_G11
XG3047 XI11_6/XI0/XI0_42/d__11_ XI11_6/XI0/XI0_42/d_11_ DECAP_INV_G11
XG3048 XI11_6/XI0/XI0_42/d__10_ XI11_6/XI0/XI0_42/d_10_ DECAP_INV_G11
XG3049 XI11_6/XI0/XI0_42/d__9_ XI11_6/XI0/XI0_42/d_9_ DECAP_INV_G11
XG3050 XI11_6/XI0/XI0_42/d__8_ XI11_6/XI0/XI0_42/d_8_ DECAP_INV_G11
XG3051 XI11_6/XI0/XI0_42/d__7_ XI11_6/XI0/XI0_42/d_7_ DECAP_INV_G11
XG3052 XI11_6/XI0/XI0_42/d__6_ XI11_6/XI0/XI0_42/d_6_ DECAP_INV_G11
XG3053 XI11_6/XI0/XI0_42/d__5_ XI11_6/XI0/XI0_42/d_5_ DECAP_INV_G11
XG3054 XI11_6/XI0/XI0_42/d__4_ XI11_6/XI0/XI0_42/d_4_ DECAP_INV_G11
XG3055 XI11_6/XI0/XI0_42/d__3_ XI11_6/XI0/XI0_42/d_3_ DECAP_INV_G11
XG3056 XI11_6/XI0/XI0_42/d__2_ XI11_6/XI0/XI0_42/d_2_ DECAP_INV_G11
XG3057 XI11_6/XI0/XI0_42/d__1_ XI11_6/XI0/XI0_42/d_1_ DECAP_INV_G11
XG3058 XI11_6/XI0/XI0_42/d__0_ XI11_6/XI0/XI0_42/d_0_ DECAP_INV_G11
XG3059 XI11_6/XI0/XI0_42/d_15_ XI11_6/XI0/XI0_42/d__15_ DECAP_INV_G11
XG3060 XI11_6/XI0/XI0_42/d_14_ XI11_6/XI0/XI0_42/d__14_ DECAP_INV_G11
XG3061 XI11_6/XI0/XI0_42/d_13_ XI11_6/XI0/XI0_42/d__13_ DECAP_INV_G11
XG3062 XI11_6/XI0/XI0_42/d_12_ XI11_6/XI0/XI0_42/d__12_ DECAP_INV_G11
XG3063 XI11_6/XI0/XI0_42/d_11_ XI11_6/XI0/XI0_42/d__11_ DECAP_INV_G11
XG3064 XI11_6/XI0/XI0_42/d_10_ XI11_6/XI0/XI0_42/d__10_ DECAP_INV_G11
XG3065 XI11_6/XI0/XI0_42/d_9_ XI11_6/XI0/XI0_42/d__9_ DECAP_INV_G11
XG3066 XI11_6/XI0/XI0_42/d_8_ XI11_6/XI0/XI0_42/d__8_ DECAP_INV_G11
XG3067 XI11_6/XI0/XI0_42/d_7_ XI11_6/XI0/XI0_42/d__7_ DECAP_INV_G11
XG3068 XI11_6/XI0/XI0_42/d_6_ XI11_6/XI0/XI0_42/d__6_ DECAP_INV_G11
XG3069 XI11_6/XI0/XI0_42/d_5_ XI11_6/XI0/XI0_42/d__5_ DECAP_INV_G11
XG3070 XI11_6/XI0/XI0_42/d_4_ XI11_6/XI0/XI0_42/d__4_ DECAP_INV_G11
XG3071 XI11_6/XI0/XI0_42/d_3_ XI11_6/XI0/XI0_42/d__3_ DECAP_INV_G11
XG3072 XI11_6/XI0/XI0_42/d_2_ XI11_6/XI0/XI0_42/d__2_ DECAP_INV_G11
XG3073 XI11_6/XI0/XI0_42/d_1_ XI11_6/XI0/XI0_42/d__1_ DECAP_INV_G11
XG3074 XI11_6/XI0/XI0_42/d_0_ XI11_6/XI0/XI0_42/d__0_ DECAP_INV_G11
XG3075 XI11_6/XI0/XI0_41/d__15_ XI11_6/XI0/XI0_41/d_15_ DECAP_INV_G11
XG3076 XI11_6/XI0/XI0_41/d__14_ XI11_6/XI0/XI0_41/d_14_ DECAP_INV_G11
XG3077 XI11_6/XI0/XI0_41/d__13_ XI11_6/XI0/XI0_41/d_13_ DECAP_INV_G11
XG3078 XI11_6/XI0/XI0_41/d__12_ XI11_6/XI0/XI0_41/d_12_ DECAP_INV_G11
XG3079 XI11_6/XI0/XI0_41/d__11_ XI11_6/XI0/XI0_41/d_11_ DECAP_INV_G11
XG3080 XI11_6/XI0/XI0_41/d__10_ XI11_6/XI0/XI0_41/d_10_ DECAP_INV_G11
XG3081 XI11_6/XI0/XI0_41/d__9_ XI11_6/XI0/XI0_41/d_9_ DECAP_INV_G11
XG3082 XI11_6/XI0/XI0_41/d__8_ XI11_6/XI0/XI0_41/d_8_ DECAP_INV_G11
XG3083 XI11_6/XI0/XI0_41/d__7_ XI11_6/XI0/XI0_41/d_7_ DECAP_INV_G11
XG3084 XI11_6/XI0/XI0_41/d__6_ XI11_6/XI0/XI0_41/d_6_ DECAP_INV_G11
XG3085 XI11_6/XI0/XI0_41/d__5_ XI11_6/XI0/XI0_41/d_5_ DECAP_INV_G11
XG3086 XI11_6/XI0/XI0_41/d__4_ XI11_6/XI0/XI0_41/d_4_ DECAP_INV_G11
XG3087 XI11_6/XI0/XI0_41/d__3_ XI11_6/XI0/XI0_41/d_3_ DECAP_INV_G11
XG3088 XI11_6/XI0/XI0_41/d__2_ XI11_6/XI0/XI0_41/d_2_ DECAP_INV_G11
XG3089 XI11_6/XI0/XI0_41/d__1_ XI11_6/XI0/XI0_41/d_1_ DECAP_INV_G11
XG3090 XI11_6/XI0/XI0_41/d__0_ XI11_6/XI0/XI0_41/d_0_ DECAP_INV_G11
XG3091 XI11_6/XI0/XI0_41/d_15_ XI11_6/XI0/XI0_41/d__15_ DECAP_INV_G11
XG3092 XI11_6/XI0/XI0_41/d_14_ XI11_6/XI0/XI0_41/d__14_ DECAP_INV_G11
XG3093 XI11_6/XI0/XI0_41/d_13_ XI11_6/XI0/XI0_41/d__13_ DECAP_INV_G11
XG3094 XI11_6/XI0/XI0_41/d_12_ XI11_6/XI0/XI0_41/d__12_ DECAP_INV_G11
XG3095 XI11_6/XI0/XI0_41/d_11_ XI11_6/XI0/XI0_41/d__11_ DECAP_INV_G11
XG3096 XI11_6/XI0/XI0_41/d_10_ XI11_6/XI0/XI0_41/d__10_ DECAP_INV_G11
XG3097 XI11_6/XI0/XI0_41/d_9_ XI11_6/XI0/XI0_41/d__9_ DECAP_INV_G11
XG3098 XI11_6/XI0/XI0_41/d_8_ XI11_6/XI0/XI0_41/d__8_ DECAP_INV_G11
XG3099 XI11_6/XI0/XI0_41/d_7_ XI11_6/XI0/XI0_41/d__7_ DECAP_INV_G11
XG3100 XI11_6/XI0/XI0_41/d_6_ XI11_6/XI0/XI0_41/d__6_ DECAP_INV_G11
XG3101 XI11_6/XI0/XI0_41/d_5_ XI11_6/XI0/XI0_41/d__5_ DECAP_INV_G11
XG3102 XI11_6/XI0/XI0_41/d_4_ XI11_6/XI0/XI0_41/d__4_ DECAP_INV_G11
XG3103 XI11_6/XI0/XI0_41/d_3_ XI11_6/XI0/XI0_41/d__3_ DECAP_INV_G11
XG3104 XI11_6/XI0/XI0_41/d_2_ XI11_6/XI0/XI0_41/d__2_ DECAP_INV_G11
XG3105 XI11_6/XI0/XI0_41/d_1_ XI11_6/XI0/XI0_41/d__1_ DECAP_INV_G11
XG3106 XI11_6/XI0/XI0_41/d_0_ XI11_6/XI0/XI0_41/d__0_ DECAP_INV_G11
XG3107 XI11_6/XI0/XI0_40/d__15_ XI11_6/XI0/XI0_40/d_15_ DECAP_INV_G11
XG3108 XI11_6/XI0/XI0_40/d__14_ XI11_6/XI0/XI0_40/d_14_ DECAP_INV_G11
XG3109 XI11_6/XI0/XI0_40/d__13_ XI11_6/XI0/XI0_40/d_13_ DECAP_INV_G11
XG3110 XI11_6/XI0/XI0_40/d__12_ XI11_6/XI0/XI0_40/d_12_ DECAP_INV_G11
XG3111 XI11_6/XI0/XI0_40/d__11_ XI11_6/XI0/XI0_40/d_11_ DECAP_INV_G11
XG3112 XI11_6/XI0/XI0_40/d__10_ XI11_6/XI0/XI0_40/d_10_ DECAP_INV_G11
XG3113 XI11_6/XI0/XI0_40/d__9_ XI11_6/XI0/XI0_40/d_9_ DECAP_INV_G11
XG3114 XI11_6/XI0/XI0_40/d__8_ XI11_6/XI0/XI0_40/d_8_ DECAP_INV_G11
XG3115 XI11_6/XI0/XI0_40/d__7_ XI11_6/XI0/XI0_40/d_7_ DECAP_INV_G11
XG3116 XI11_6/XI0/XI0_40/d__6_ XI11_6/XI0/XI0_40/d_6_ DECAP_INV_G11
XG3117 XI11_6/XI0/XI0_40/d__5_ XI11_6/XI0/XI0_40/d_5_ DECAP_INV_G11
XG3118 XI11_6/XI0/XI0_40/d__4_ XI11_6/XI0/XI0_40/d_4_ DECAP_INV_G11
XG3119 XI11_6/XI0/XI0_40/d__3_ XI11_6/XI0/XI0_40/d_3_ DECAP_INV_G11
XG3120 XI11_6/XI0/XI0_40/d__2_ XI11_6/XI0/XI0_40/d_2_ DECAP_INV_G11
XG3121 XI11_6/XI0/XI0_40/d__1_ XI11_6/XI0/XI0_40/d_1_ DECAP_INV_G11
XG3122 XI11_6/XI0/XI0_40/d__0_ XI11_6/XI0/XI0_40/d_0_ DECAP_INV_G11
XG3123 XI11_6/XI0/XI0_40/d_15_ XI11_6/XI0/XI0_40/d__15_ DECAP_INV_G11
XG3124 XI11_6/XI0/XI0_40/d_14_ XI11_6/XI0/XI0_40/d__14_ DECAP_INV_G11
XG3125 XI11_6/XI0/XI0_40/d_13_ XI11_6/XI0/XI0_40/d__13_ DECAP_INV_G11
XG3126 XI11_6/XI0/XI0_40/d_12_ XI11_6/XI0/XI0_40/d__12_ DECAP_INV_G11
XG3127 XI11_6/XI0/XI0_40/d_11_ XI11_6/XI0/XI0_40/d__11_ DECAP_INV_G11
XG3128 XI11_6/XI0/XI0_40/d_10_ XI11_6/XI0/XI0_40/d__10_ DECAP_INV_G11
XG3129 XI11_6/XI0/XI0_40/d_9_ XI11_6/XI0/XI0_40/d__9_ DECAP_INV_G11
XG3130 XI11_6/XI0/XI0_40/d_8_ XI11_6/XI0/XI0_40/d__8_ DECAP_INV_G11
XG3131 XI11_6/XI0/XI0_40/d_7_ XI11_6/XI0/XI0_40/d__7_ DECAP_INV_G11
XG3132 XI11_6/XI0/XI0_40/d_6_ XI11_6/XI0/XI0_40/d__6_ DECAP_INV_G11
XG3133 XI11_6/XI0/XI0_40/d_5_ XI11_6/XI0/XI0_40/d__5_ DECAP_INV_G11
XG3134 XI11_6/XI0/XI0_40/d_4_ XI11_6/XI0/XI0_40/d__4_ DECAP_INV_G11
XG3135 XI11_6/XI0/XI0_40/d_3_ XI11_6/XI0/XI0_40/d__3_ DECAP_INV_G11
XG3136 XI11_6/XI0/XI0_40/d_2_ XI11_6/XI0/XI0_40/d__2_ DECAP_INV_G11
XG3137 XI11_6/XI0/XI0_40/d_1_ XI11_6/XI0/XI0_40/d__1_ DECAP_INV_G11
XG3138 XI11_6/XI0/XI0_40/d_0_ XI11_6/XI0/XI0_40/d__0_ DECAP_INV_G11
XG3139 XI11_6/XI0/XI0_39/d__15_ XI11_6/XI0/XI0_39/d_15_ DECAP_INV_G11
XG3140 XI11_6/XI0/XI0_39/d__14_ XI11_6/XI0/XI0_39/d_14_ DECAP_INV_G11
XG3141 XI11_6/XI0/XI0_39/d__13_ XI11_6/XI0/XI0_39/d_13_ DECAP_INV_G11
XG3142 XI11_6/XI0/XI0_39/d__12_ XI11_6/XI0/XI0_39/d_12_ DECAP_INV_G11
XG3143 XI11_6/XI0/XI0_39/d__11_ XI11_6/XI0/XI0_39/d_11_ DECAP_INV_G11
XG3144 XI11_6/XI0/XI0_39/d__10_ XI11_6/XI0/XI0_39/d_10_ DECAP_INV_G11
XG3145 XI11_6/XI0/XI0_39/d__9_ XI11_6/XI0/XI0_39/d_9_ DECAP_INV_G11
XG3146 XI11_6/XI0/XI0_39/d__8_ XI11_6/XI0/XI0_39/d_8_ DECAP_INV_G11
XG3147 XI11_6/XI0/XI0_39/d__7_ XI11_6/XI0/XI0_39/d_7_ DECAP_INV_G11
XG3148 XI11_6/XI0/XI0_39/d__6_ XI11_6/XI0/XI0_39/d_6_ DECAP_INV_G11
XG3149 XI11_6/XI0/XI0_39/d__5_ XI11_6/XI0/XI0_39/d_5_ DECAP_INV_G11
XG3150 XI11_6/XI0/XI0_39/d__4_ XI11_6/XI0/XI0_39/d_4_ DECAP_INV_G11
XG3151 XI11_6/XI0/XI0_39/d__3_ XI11_6/XI0/XI0_39/d_3_ DECAP_INV_G11
XG3152 XI11_6/XI0/XI0_39/d__2_ XI11_6/XI0/XI0_39/d_2_ DECAP_INV_G11
XG3153 XI11_6/XI0/XI0_39/d__1_ XI11_6/XI0/XI0_39/d_1_ DECAP_INV_G11
XG3154 XI11_6/XI0/XI0_39/d__0_ XI11_6/XI0/XI0_39/d_0_ DECAP_INV_G11
XG3155 XI11_6/XI0/XI0_39/d_15_ XI11_6/XI0/XI0_39/d__15_ DECAP_INV_G11
XG3156 XI11_6/XI0/XI0_39/d_14_ XI11_6/XI0/XI0_39/d__14_ DECAP_INV_G11
XG3157 XI11_6/XI0/XI0_39/d_13_ XI11_6/XI0/XI0_39/d__13_ DECAP_INV_G11
XG3158 XI11_6/XI0/XI0_39/d_12_ XI11_6/XI0/XI0_39/d__12_ DECAP_INV_G11
XG3159 XI11_6/XI0/XI0_39/d_11_ XI11_6/XI0/XI0_39/d__11_ DECAP_INV_G11
XG3160 XI11_6/XI0/XI0_39/d_10_ XI11_6/XI0/XI0_39/d__10_ DECAP_INV_G11
XG3161 XI11_6/XI0/XI0_39/d_9_ XI11_6/XI0/XI0_39/d__9_ DECAP_INV_G11
XG3162 XI11_6/XI0/XI0_39/d_8_ XI11_6/XI0/XI0_39/d__8_ DECAP_INV_G11
XG3163 XI11_6/XI0/XI0_39/d_7_ XI11_6/XI0/XI0_39/d__7_ DECAP_INV_G11
XG3164 XI11_6/XI0/XI0_39/d_6_ XI11_6/XI0/XI0_39/d__6_ DECAP_INV_G11
XG3165 XI11_6/XI0/XI0_39/d_5_ XI11_6/XI0/XI0_39/d__5_ DECAP_INV_G11
XG3166 XI11_6/XI0/XI0_39/d_4_ XI11_6/XI0/XI0_39/d__4_ DECAP_INV_G11
XG3167 XI11_6/XI0/XI0_39/d_3_ XI11_6/XI0/XI0_39/d__3_ DECAP_INV_G11
XG3168 XI11_6/XI0/XI0_39/d_2_ XI11_6/XI0/XI0_39/d__2_ DECAP_INV_G11
XG3169 XI11_6/XI0/XI0_39/d_1_ XI11_6/XI0/XI0_39/d__1_ DECAP_INV_G11
XG3170 XI11_6/XI0/XI0_39/d_0_ XI11_6/XI0/XI0_39/d__0_ DECAP_INV_G11
XG3171 XI11_6/XI0/XI0_38/d__15_ XI11_6/XI0/XI0_38/d_15_ DECAP_INV_G11
XG3172 XI11_6/XI0/XI0_38/d__14_ XI11_6/XI0/XI0_38/d_14_ DECAP_INV_G11
XG3173 XI11_6/XI0/XI0_38/d__13_ XI11_6/XI0/XI0_38/d_13_ DECAP_INV_G11
XG3174 XI11_6/XI0/XI0_38/d__12_ XI11_6/XI0/XI0_38/d_12_ DECAP_INV_G11
XG3175 XI11_6/XI0/XI0_38/d__11_ XI11_6/XI0/XI0_38/d_11_ DECAP_INV_G11
XG3176 XI11_6/XI0/XI0_38/d__10_ XI11_6/XI0/XI0_38/d_10_ DECAP_INV_G11
XG3177 XI11_6/XI0/XI0_38/d__9_ XI11_6/XI0/XI0_38/d_9_ DECAP_INV_G11
XG3178 XI11_6/XI0/XI0_38/d__8_ XI11_6/XI0/XI0_38/d_8_ DECAP_INV_G11
XG3179 XI11_6/XI0/XI0_38/d__7_ XI11_6/XI0/XI0_38/d_7_ DECAP_INV_G11
XG3180 XI11_6/XI0/XI0_38/d__6_ XI11_6/XI0/XI0_38/d_6_ DECAP_INV_G11
XG3181 XI11_6/XI0/XI0_38/d__5_ XI11_6/XI0/XI0_38/d_5_ DECAP_INV_G11
XG3182 XI11_6/XI0/XI0_38/d__4_ XI11_6/XI0/XI0_38/d_4_ DECAP_INV_G11
XG3183 XI11_6/XI0/XI0_38/d__3_ XI11_6/XI0/XI0_38/d_3_ DECAP_INV_G11
XG3184 XI11_6/XI0/XI0_38/d__2_ XI11_6/XI0/XI0_38/d_2_ DECAP_INV_G11
XG3185 XI11_6/XI0/XI0_38/d__1_ XI11_6/XI0/XI0_38/d_1_ DECAP_INV_G11
XG3186 XI11_6/XI0/XI0_38/d__0_ XI11_6/XI0/XI0_38/d_0_ DECAP_INV_G11
XG3187 XI11_6/XI0/XI0_38/d_15_ XI11_6/XI0/XI0_38/d__15_ DECAP_INV_G11
XG3188 XI11_6/XI0/XI0_38/d_14_ XI11_6/XI0/XI0_38/d__14_ DECAP_INV_G11
XG3189 XI11_6/XI0/XI0_38/d_13_ XI11_6/XI0/XI0_38/d__13_ DECAP_INV_G11
XG3190 XI11_6/XI0/XI0_38/d_12_ XI11_6/XI0/XI0_38/d__12_ DECAP_INV_G11
XG3191 XI11_6/XI0/XI0_38/d_11_ XI11_6/XI0/XI0_38/d__11_ DECAP_INV_G11
XG3192 XI11_6/XI0/XI0_38/d_10_ XI11_6/XI0/XI0_38/d__10_ DECAP_INV_G11
XG3193 XI11_6/XI0/XI0_38/d_9_ XI11_6/XI0/XI0_38/d__9_ DECAP_INV_G11
XG3194 XI11_6/XI0/XI0_38/d_8_ XI11_6/XI0/XI0_38/d__8_ DECAP_INV_G11
XG3195 XI11_6/XI0/XI0_38/d_7_ XI11_6/XI0/XI0_38/d__7_ DECAP_INV_G11
XG3196 XI11_6/XI0/XI0_38/d_6_ XI11_6/XI0/XI0_38/d__6_ DECAP_INV_G11
XG3197 XI11_6/XI0/XI0_38/d_5_ XI11_6/XI0/XI0_38/d__5_ DECAP_INV_G11
XG3198 XI11_6/XI0/XI0_38/d_4_ XI11_6/XI0/XI0_38/d__4_ DECAP_INV_G11
XG3199 XI11_6/XI0/XI0_38/d_3_ XI11_6/XI0/XI0_38/d__3_ DECAP_INV_G11
XG3200 XI11_6/XI0/XI0_38/d_2_ XI11_6/XI0/XI0_38/d__2_ DECAP_INV_G11
XG3201 XI11_6/XI0/XI0_38/d_1_ XI11_6/XI0/XI0_38/d__1_ DECAP_INV_G11
XG3202 XI11_6/XI0/XI0_38/d_0_ XI11_6/XI0/XI0_38/d__0_ DECAP_INV_G11
XG3203 XI11_6/XI0/XI0_37/d__15_ XI11_6/XI0/XI0_37/d_15_ DECAP_INV_G11
XG3204 XI11_6/XI0/XI0_37/d__14_ XI11_6/XI0/XI0_37/d_14_ DECAP_INV_G11
XG3205 XI11_6/XI0/XI0_37/d__13_ XI11_6/XI0/XI0_37/d_13_ DECAP_INV_G11
XG3206 XI11_6/XI0/XI0_37/d__12_ XI11_6/XI0/XI0_37/d_12_ DECAP_INV_G11
XG3207 XI11_6/XI0/XI0_37/d__11_ XI11_6/XI0/XI0_37/d_11_ DECAP_INV_G11
XG3208 XI11_6/XI0/XI0_37/d__10_ XI11_6/XI0/XI0_37/d_10_ DECAP_INV_G11
XG3209 XI11_6/XI0/XI0_37/d__9_ XI11_6/XI0/XI0_37/d_9_ DECAP_INV_G11
XG3210 XI11_6/XI0/XI0_37/d__8_ XI11_6/XI0/XI0_37/d_8_ DECAP_INV_G11
XG3211 XI11_6/XI0/XI0_37/d__7_ XI11_6/XI0/XI0_37/d_7_ DECAP_INV_G11
XG3212 XI11_6/XI0/XI0_37/d__6_ XI11_6/XI0/XI0_37/d_6_ DECAP_INV_G11
XG3213 XI11_6/XI0/XI0_37/d__5_ XI11_6/XI0/XI0_37/d_5_ DECAP_INV_G11
XG3214 XI11_6/XI0/XI0_37/d__4_ XI11_6/XI0/XI0_37/d_4_ DECAP_INV_G11
XG3215 XI11_6/XI0/XI0_37/d__3_ XI11_6/XI0/XI0_37/d_3_ DECAP_INV_G11
XG3216 XI11_6/XI0/XI0_37/d__2_ XI11_6/XI0/XI0_37/d_2_ DECAP_INV_G11
XG3217 XI11_6/XI0/XI0_37/d__1_ XI11_6/XI0/XI0_37/d_1_ DECAP_INV_G11
XG3218 XI11_6/XI0/XI0_37/d__0_ XI11_6/XI0/XI0_37/d_0_ DECAP_INV_G11
XG3219 XI11_6/XI0/XI0_37/d_15_ XI11_6/XI0/XI0_37/d__15_ DECAP_INV_G11
XG3220 XI11_6/XI0/XI0_37/d_14_ XI11_6/XI0/XI0_37/d__14_ DECAP_INV_G11
XG3221 XI11_6/XI0/XI0_37/d_13_ XI11_6/XI0/XI0_37/d__13_ DECAP_INV_G11
XG3222 XI11_6/XI0/XI0_37/d_12_ XI11_6/XI0/XI0_37/d__12_ DECAP_INV_G11
XG3223 XI11_6/XI0/XI0_37/d_11_ XI11_6/XI0/XI0_37/d__11_ DECAP_INV_G11
XG3224 XI11_6/XI0/XI0_37/d_10_ XI11_6/XI0/XI0_37/d__10_ DECAP_INV_G11
XG3225 XI11_6/XI0/XI0_37/d_9_ XI11_6/XI0/XI0_37/d__9_ DECAP_INV_G11
XG3226 XI11_6/XI0/XI0_37/d_8_ XI11_6/XI0/XI0_37/d__8_ DECAP_INV_G11
XG3227 XI11_6/XI0/XI0_37/d_7_ XI11_6/XI0/XI0_37/d__7_ DECAP_INV_G11
XG3228 XI11_6/XI0/XI0_37/d_6_ XI11_6/XI0/XI0_37/d__6_ DECAP_INV_G11
XG3229 XI11_6/XI0/XI0_37/d_5_ XI11_6/XI0/XI0_37/d__5_ DECAP_INV_G11
XG3230 XI11_6/XI0/XI0_37/d_4_ XI11_6/XI0/XI0_37/d__4_ DECAP_INV_G11
XG3231 XI11_6/XI0/XI0_37/d_3_ XI11_6/XI0/XI0_37/d__3_ DECAP_INV_G11
XG3232 XI11_6/XI0/XI0_37/d_2_ XI11_6/XI0/XI0_37/d__2_ DECAP_INV_G11
XG3233 XI11_6/XI0/XI0_37/d_1_ XI11_6/XI0/XI0_37/d__1_ DECAP_INV_G11
XG3234 XI11_6/XI0/XI0_37/d_0_ XI11_6/XI0/XI0_37/d__0_ DECAP_INV_G11
XG3235 XI11_6/XI0/XI0_36/d__15_ XI11_6/XI0/XI0_36/d_15_ DECAP_INV_G11
XG3236 XI11_6/XI0/XI0_36/d__14_ XI11_6/XI0/XI0_36/d_14_ DECAP_INV_G11
XG3237 XI11_6/XI0/XI0_36/d__13_ XI11_6/XI0/XI0_36/d_13_ DECAP_INV_G11
XG3238 XI11_6/XI0/XI0_36/d__12_ XI11_6/XI0/XI0_36/d_12_ DECAP_INV_G11
XG3239 XI11_6/XI0/XI0_36/d__11_ XI11_6/XI0/XI0_36/d_11_ DECAP_INV_G11
XG3240 XI11_6/XI0/XI0_36/d__10_ XI11_6/XI0/XI0_36/d_10_ DECAP_INV_G11
XG3241 XI11_6/XI0/XI0_36/d__9_ XI11_6/XI0/XI0_36/d_9_ DECAP_INV_G11
XG3242 XI11_6/XI0/XI0_36/d__8_ XI11_6/XI0/XI0_36/d_8_ DECAP_INV_G11
XG3243 XI11_6/XI0/XI0_36/d__7_ XI11_6/XI0/XI0_36/d_7_ DECAP_INV_G11
XG3244 XI11_6/XI0/XI0_36/d__6_ XI11_6/XI0/XI0_36/d_6_ DECAP_INV_G11
XG3245 XI11_6/XI0/XI0_36/d__5_ XI11_6/XI0/XI0_36/d_5_ DECAP_INV_G11
XG3246 XI11_6/XI0/XI0_36/d__4_ XI11_6/XI0/XI0_36/d_4_ DECAP_INV_G11
XG3247 XI11_6/XI0/XI0_36/d__3_ XI11_6/XI0/XI0_36/d_3_ DECAP_INV_G11
XG3248 XI11_6/XI0/XI0_36/d__2_ XI11_6/XI0/XI0_36/d_2_ DECAP_INV_G11
XG3249 XI11_6/XI0/XI0_36/d__1_ XI11_6/XI0/XI0_36/d_1_ DECAP_INV_G11
XG3250 XI11_6/XI0/XI0_36/d__0_ XI11_6/XI0/XI0_36/d_0_ DECAP_INV_G11
XG3251 XI11_6/XI0/XI0_36/d_15_ XI11_6/XI0/XI0_36/d__15_ DECAP_INV_G11
XG3252 XI11_6/XI0/XI0_36/d_14_ XI11_6/XI0/XI0_36/d__14_ DECAP_INV_G11
XG3253 XI11_6/XI0/XI0_36/d_13_ XI11_6/XI0/XI0_36/d__13_ DECAP_INV_G11
XG3254 XI11_6/XI0/XI0_36/d_12_ XI11_6/XI0/XI0_36/d__12_ DECAP_INV_G11
XG3255 XI11_6/XI0/XI0_36/d_11_ XI11_6/XI0/XI0_36/d__11_ DECAP_INV_G11
XG3256 XI11_6/XI0/XI0_36/d_10_ XI11_6/XI0/XI0_36/d__10_ DECAP_INV_G11
XG3257 XI11_6/XI0/XI0_36/d_9_ XI11_6/XI0/XI0_36/d__9_ DECAP_INV_G11
XG3258 XI11_6/XI0/XI0_36/d_8_ XI11_6/XI0/XI0_36/d__8_ DECAP_INV_G11
XG3259 XI11_6/XI0/XI0_36/d_7_ XI11_6/XI0/XI0_36/d__7_ DECAP_INV_G11
XG3260 XI11_6/XI0/XI0_36/d_6_ XI11_6/XI0/XI0_36/d__6_ DECAP_INV_G11
XG3261 XI11_6/XI0/XI0_36/d_5_ XI11_6/XI0/XI0_36/d__5_ DECAP_INV_G11
XG3262 XI11_6/XI0/XI0_36/d_4_ XI11_6/XI0/XI0_36/d__4_ DECAP_INV_G11
XG3263 XI11_6/XI0/XI0_36/d_3_ XI11_6/XI0/XI0_36/d__3_ DECAP_INV_G11
XG3264 XI11_6/XI0/XI0_36/d_2_ XI11_6/XI0/XI0_36/d__2_ DECAP_INV_G11
XG3265 XI11_6/XI0/XI0_36/d_1_ XI11_6/XI0/XI0_36/d__1_ DECAP_INV_G11
XG3266 XI11_6/XI0/XI0_36/d_0_ XI11_6/XI0/XI0_36/d__0_ DECAP_INV_G11
XG3267 XI11_6/XI0/XI0_35/d__15_ XI11_6/XI0/XI0_35/d_15_ DECAP_INV_G11
XG3268 XI11_6/XI0/XI0_35/d__14_ XI11_6/XI0/XI0_35/d_14_ DECAP_INV_G11
XG3269 XI11_6/XI0/XI0_35/d__13_ XI11_6/XI0/XI0_35/d_13_ DECAP_INV_G11
XG3270 XI11_6/XI0/XI0_35/d__12_ XI11_6/XI0/XI0_35/d_12_ DECAP_INV_G11
XG3271 XI11_6/XI0/XI0_35/d__11_ XI11_6/XI0/XI0_35/d_11_ DECAP_INV_G11
XG3272 XI11_6/XI0/XI0_35/d__10_ XI11_6/XI0/XI0_35/d_10_ DECAP_INV_G11
XG3273 XI11_6/XI0/XI0_35/d__9_ XI11_6/XI0/XI0_35/d_9_ DECAP_INV_G11
XG3274 XI11_6/XI0/XI0_35/d__8_ XI11_6/XI0/XI0_35/d_8_ DECAP_INV_G11
XG3275 XI11_6/XI0/XI0_35/d__7_ XI11_6/XI0/XI0_35/d_7_ DECAP_INV_G11
XG3276 XI11_6/XI0/XI0_35/d__6_ XI11_6/XI0/XI0_35/d_6_ DECAP_INV_G11
XG3277 XI11_6/XI0/XI0_35/d__5_ XI11_6/XI0/XI0_35/d_5_ DECAP_INV_G11
XG3278 XI11_6/XI0/XI0_35/d__4_ XI11_6/XI0/XI0_35/d_4_ DECAP_INV_G11
XG3279 XI11_6/XI0/XI0_35/d__3_ XI11_6/XI0/XI0_35/d_3_ DECAP_INV_G11
XG3280 XI11_6/XI0/XI0_35/d__2_ XI11_6/XI0/XI0_35/d_2_ DECAP_INV_G11
XG3281 XI11_6/XI0/XI0_35/d__1_ XI11_6/XI0/XI0_35/d_1_ DECAP_INV_G11
XG3282 XI11_6/XI0/XI0_35/d__0_ XI11_6/XI0/XI0_35/d_0_ DECAP_INV_G11
XG3283 XI11_6/XI0/XI0_35/d_15_ XI11_6/XI0/XI0_35/d__15_ DECAP_INV_G11
XG3284 XI11_6/XI0/XI0_35/d_14_ XI11_6/XI0/XI0_35/d__14_ DECAP_INV_G11
XG3285 XI11_6/XI0/XI0_35/d_13_ XI11_6/XI0/XI0_35/d__13_ DECAP_INV_G11
XG3286 XI11_6/XI0/XI0_35/d_12_ XI11_6/XI0/XI0_35/d__12_ DECAP_INV_G11
XG3287 XI11_6/XI0/XI0_35/d_11_ XI11_6/XI0/XI0_35/d__11_ DECAP_INV_G11
XG3288 XI11_6/XI0/XI0_35/d_10_ XI11_6/XI0/XI0_35/d__10_ DECAP_INV_G11
XG3289 XI11_6/XI0/XI0_35/d_9_ XI11_6/XI0/XI0_35/d__9_ DECAP_INV_G11
XG3290 XI11_6/XI0/XI0_35/d_8_ XI11_6/XI0/XI0_35/d__8_ DECAP_INV_G11
XG3291 XI11_6/XI0/XI0_35/d_7_ XI11_6/XI0/XI0_35/d__7_ DECAP_INV_G11
XG3292 XI11_6/XI0/XI0_35/d_6_ XI11_6/XI0/XI0_35/d__6_ DECAP_INV_G11
XG3293 XI11_6/XI0/XI0_35/d_5_ XI11_6/XI0/XI0_35/d__5_ DECAP_INV_G11
XG3294 XI11_6/XI0/XI0_35/d_4_ XI11_6/XI0/XI0_35/d__4_ DECAP_INV_G11
XG3295 XI11_6/XI0/XI0_35/d_3_ XI11_6/XI0/XI0_35/d__3_ DECAP_INV_G11
XG3296 XI11_6/XI0/XI0_35/d_2_ XI11_6/XI0/XI0_35/d__2_ DECAP_INV_G11
XG3297 XI11_6/XI0/XI0_35/d_1_ XI11_6/XI0/XI0_35/d__1_ DECAP_INV_G11
XG3298 XI11_6/XI0/XI0_35/d_0_ XI11_6/XI0/XI0_35/d__0_ DECAP_INV_G11
XG3299 XI11_6/XI0/XI0_34/d__15_ XI11_6/XI0/XI0_34/d_15_ DECAP_INV_G11
XG3300 XI11_6/XI0/XI0_34/d__14_ XI11_6/XI0/XI0_34/d_14_ DECAP_INV_G11
XG3301 XI11_6/XI0/XI0_34/d__13_ XI11_6/XI0/XI0_34/d_13_ DECAP_INV_G11
XG3302 XI11_6/XI0/XI0_34/d__12_ XI11_6/XI0/XI0_34/d_12_ DECAP_INV_G11
XG3303 XI11_6/XI0/XI0_34/d__11_ XI11_6/XI0/XI0_34/d_11_ DECAP_INV_G11
XG3304 XI11_6/XI0/XI0_34/d__10_ XI11_6/XI0/XI0_34/d_10_ DECAP_INV_G11
XG3305 XI11_6/XI0/XI0_34/d__9_ XI11_6/XI0/XI0_34/d_9_ DECAP_INV_G11
XG3306 XI11_6/XI0/XI0_34/d__8_ XI11_6/XI0/XI0_34/d_8_ DECAP_INV_G11
XG3307 XI11_6/XI0/XI0_34/d__7_ XI11_6/XI0/XI0_34/d_7_ DECAP_INV_G11
XG3308 XI11_6/XI0/XI0_34/d__6_ XI11_6/XI0/XI0_34/d_6_ DECAP_INV_G11
XG3309 XI11_6/XI0/XI0_34/d__5_ XI11_6/XI0/XI0_34/d_5_ DECAP_INV_G11
XG3310 XI11_6/XI0/XI0_34/d__4_ XI11_6/XI0/XI0_34/d_4_ DECAP_INV_G11
XG3311 XI11_6/XI0/XI0_34/d__3_ XI11_6/XI0/XI0_34/d_3_ DECAP_INV_G11
XG3312 XI11_6/XI0/XI0_34/d__2_ XI11_6/XI0/XI0_34/d_2_ DECAP_INV_G11
XG3313 XI11_6/XI0/XI0_34/d__1_ XI11_6/XI0/XI0_34/d_1_ DECAP_INV_G11
XG3314 XI11_6/XI0/XI0_34/d__0_ XI11_6/XI0/XI0_34/d_0_ DECAP_INV_G11
XG3315 XI11_6/XI0/XI0_34/d_15_ XI11_6/XI0/XI0_34/d__15_ DECAP_INV_G11
XG3316 XI11_6/XI0/XI0_34/d_14_ XI11_6/XI0/XI0_34/d__14_ DECAP_INV_G11
XG3317 XI11_6/XI0/XI0_34/d_13_ XI11_6/XI0/XI0_34/d__13_ DECAP_INV_G11
XG3318 XI11_6/XI0/XI0_34/d_12_ XI11_6/XI0/XI0_34/d__12_ DECAP_INV_G11
XG3319 XI11_6/XI0/XI0_34/d_11_ XI11_6/XI0/XI0_34/d__11_ DECAP_INV_G11
XG3320 XI11_6/XI0/XI0_34/d_10_ XI11_6/XI0/XI0_34/d__10_ DECAP_INV_G11
XG3321 XI11_6/XI0/XI0_34/d_9_ XI11_6/XI0/XI0_34/d__9_ DECAP_INV_G11
XG3322 XI11_6/XI0/XI0_34/d_8_ XI11_6/XI0/XI0_34/d__8_ DECAP_INV_G11
XG3323 XI11_6/XI0/XI0_34/d_7_ XI11_6/XI0/XI0_34/d__7_ DECAP_INV_G11
XG3324 XI11_6/XI0/XI0_34/d_6_ XI11_6/XI0/XI0_34/d__6_ DECAP_INV_G11
XG3325 XI11_6/XI0/XI0_34/d_5_ XI11_6/XI0/XI0_34/d__5_ DECAP_INV_G11
XG3326 XI11_6/XI0/XI0_34/d_4_ XI11_6/XI0/XI0_34/d__4_ DECAP_INV_G11
XG3327 XI11_6/XI0/XI0_34/d_3_ XI11_6/XI0/XI0_34/d__3_ DECAP_INV_G11
XG3328 XI11_6/XI0/XI0_34/d_2_ XI11_6/XI0/XI0_34/d__2_ DECAP_INV_G11
XG3329 XI11_6/XI0/XI0_34/d_1_ XI11_6/XI0/XI0_34/d__1_ DECAP_INV_G11
XG3330 XI11_6/XI0/XI0_34/d_0_ XI11_6/XI0/XI0_34/d__0_ DECAP_INV_G11
XG3331 XI11_6/XI0/XI0_33/d__15_ XI11_6/XI0/XI0_33/d_15_ DECAP_INV_G11
XG3332 XI11_6/XI0/XI0_33/d__14_ XI11_6/XI0/XI0_33/d_14_ DECAP_INV_G11
XG3333 XI11_6/XI0/XI0_33/d__13_ XI11_6/XI0/XI0_33/d_13_ DECAP_INV_G11
XG3334 XI11_6/XI0/XI0_33/d__12_ XI11_6/XI0/XI0_33/d_12_ DECAP_INV_G11
XG3335 XI11_6/XI0/XI0_33/d__11_ XI11_6/XI0/XI0_33/d_11_ DECAP_INV_G11
XG3336 XI11_6/XI0/XI0_33/d__10_ XI11_6/XI0/XI0_33/d_10_ DECAP_INV_G11
XG3337 XI11_6/XI0/XI0_33/d__9_ XI11_6/XI0/XI0_33/d_9_ DECAP_INV_G11
XG3338 XI11_6/XI0/XI0_33/d__8_ XI11_6/XI0/XI0_33/d_8_ DECAP_INV_G11
XG3339 XI11_6/XI0/XI0_33/d__7_ XI11_6/XI0/XI0_33/d_7_ DECAP_INV_G11
XG3340 XI11_6/XI0/XI0_33/d__6_ XI11_6/XI0/XI0_33/d_6_ DECAP_INV_G11
XG3341 XI11_6/XI0/XI0_33/d__5_ XI11_6/XI0/XI0_33/d_5_ DECAP_INV_G11
XG3342 XI11_6/XI0/XI0_33/d__4_ XI11_6/XI0/XI0_33/d_4_ DECAP_INV_G11
XG3343 XI11_6/XI0/XI0_33/d__3_ XI11_6/XI0/XI0_33/d_3_ DECAP_INV_G11
XG3344 XI11_6/XI0/XI0_33/d__2_ XI11_6/XI0/XI0_33/d_2_ DECAP_INV_G11
XG3345 XI11_6/XI0/XI0_33/d__1_ XI11_6/XI0/XI0_33/d_1_ DECAP_INV_G11
XG3346 XI11_6/XI0/XI0_33/d__0_ XI11_6/XI0/XI0_33/d_0_ DECAP_INV_G11
XG3347 XI11_6/XI0/XI0_33/d_15_ XI11_6/XI0/XI0_33/d__15_ DECAP_INV_G11
XG3348 XI11_6/XI0/XI0_33/d_14_ XI11_6/XI0/XI0_33/d__14_ DECAP_INV_G11
XG3349 XI11_6/XI0/XI0_33/d_13_ XI11_6/XI0/XI0_33/d__13_ DECAP_INV_G11
XG3350 XI11_6/XI0/XI0_33/d_12_ XI11_6/XI0/XI0_33/d__12_ DECAP_INV_G11
XG3351 XI11_6/XI0/XI0_33/d_11_ XI11_6/XI0/XI0_33/d__11_ DECAP_INV_G11
XG3352 XI11_6/XI0/XI0_33/d_10_ XI11_6/XI0/XI0_33/d__10_ DECAP_INV_G11
XG3353 XI11_6/XI0/XI0_33/d_9_ XI11_6/XI0/XI0_33/d__9_ DECAP_INV_G11
XG3354 XI11_6/XI0/XI0_33/d_8_ XI11_6/XI0/XI0_33/d__8_ DECAP_INV_G11
XG3355 XI11_6/XI0/XI0_33/d_7_ XI11_6/XI0/XI0_33/d__7_ DECAP_INV_G11
XG3356 XI11_6/XI0/XI0_33/d_6_ XI11_6/XI0/XI0_33/d__6_ DECAP_INV_G11
XG3357 XI11_6/XI0/XI0_33/d_5_ XI11_6/XI0/XI0_33/d__5_ DECAP_INV_G11
XG3358 XI11_6/XI0/XI0_33/d_4_ XI11_6/XI0/XI0_33/d__4_ DECAP_INV_G11
XG3359 XI11_6/XI0/XI0_33/d_3_ XI11_6/XI0/XI0_33/d__3_ DECAP_INV_G11
XG3360 XI11_6/XI0/XI0_33/d_2_ XI11_6/XI0/XI0_33/d__2_ DECAP_INV_G11
XG3361 XI11_6/XI0/XI0_33/d_1_ XI11_6/XI0/XI0_33/d__1_ DECAP_INV_G11
XG3362 XI11_6/XI0/XI0_33/d_0_ XI11_6/XI0/XI0_33/d__0_ DECAP_INV_G11
XG3363 XI11_6/XI0/XI0_32/d__15_ XI11_6/XI0/XI0_32/d_15_ DECAP_INV_G11
XG3364 XI11_6/XI0/XI0_32/d__14_ XI11_6/XI0/XI0_32/d_14_ DECAP_INV_G11
XG3365 XI11_6/XI0/XI0_32/d__13_ XI11_6/XI0/XI0_32/d_13_ DECAP_INV_G11
XG3366 XI11_6/XI0/XI0_32/d__12_ XI11_6/XI0/XI0_32/d_12_ DECAP_INV_G11
XG3367 XI11_6/XI0/XI0_32/d__11_ XI11_6/XI0/XI0_32/d_11_ DECAP_INV_G11
XG3368 XI11_6/XI0/XI0_32/d__10_ XI11_6/XI0/XI0_32/d_10_ DECAP_INV_G11
XG3369 XI11_6/XI0/XI0_32/d__9_ XI11_6/XI0/XI0_32/d_9_ DECAP_INV_G11
XG3370 XI11_6/XI0/XI0_32/d__8_ XI11_6/XI0/XI0_32/d_8_ DECAP_INV_G11
XG3371 XI11_6/XI0/XI0_32/d__7_ XI11_6/XI0/XI0_32/d_7_ DECAP_INV_G11
XG3372 XI11_6/XI0/XI0_32/d__6_ XI11_6/XI0/XI0_32/d_6_ DECAP_INV_G11
XG3373 XI11_6/XI0/XI0_32/d__5_ XI11_6/XI0/XI0_32/d_5_ DECAP_INV_G11
XG3374 XI11_6/XI0/XI0_32/d__4_ XI11_6/XI0/XI0_32/d_4_ DECAP_INV_G11
XG3375 XI11_6/XI0/XI0_32/d__3_ XI11_6/XI0/XI0_32/d_3_ DECAP_INV_G11
XG3376 XI11_6/XI0/XI0_32/d__2_ XI11_6/XI0/XI0_32/d_2_ DECAP_INV_G11
XG3377 XI11_6/XI0/XI0_32/d__1_ XI11_6/XI0/XI0_32/d_1_ DECAP_INV_G11
XG3378 XI11_6/XI0/XI0_32/d__0_ XI11_6/XI0/XI0_32/d_0_ DECAP_INV_G11
XG3379 XI11_6/XI0/XI0_32/d_15_ XI11_6/XI0/XI0_32/d__15_ DECAP_INV_G11
XG3380 XI11_6/XI0/XI0_32/d_14_ XI11_6/XI0/XI0_32/d__14_ DECAP_INV_G11
XG3381 XI11_6/XI0/XI0_32/d_13_ XI11_6/XI0/XI0_32/d__13_ DECAP_INV_G11
XG3382 XI11_6/XI0/XI0_32/d_12_ XI11_6/XI0/XI0_32/d__12_ DECAP_INV_G11
XG3383 XI11_6/XI0/XI0_32/d_11_ XI11_6/XI0/XI0_32/d__11_ DECAP_INV_G11
XG3384 XI11_6/XI0/XI0_32/d_10_ XI11_6/XI0/XI0_32/d__10_ DECAP_INV_G11
XG3385 XI11_6/XI0/XI0_32/d_9_ XI11_6/XI0/XI0_32/d__9_ DECAP_INV_G11
XG3386 XI11_6/XI0/XI0_32/d_8_ XI11_6/XI0/XI0_32/d__8_ DECAP_INV_G11
XG3387 XI11_6/XI0/XI0_32/d_7_ XI11_6/XI0/XI0_32/d__7_ DECAP_INV_G11
XG3388 XI11_6/XI0/XI0_32/d_6_ XI11_6/XI0/XI0_32/d__6_ DECAP_INV_G11
XG3389 XI11_6/XI0/XI0_32/d_5_ XI11_6/XI0/XI0_32/d__5_ DECAP_INV_G11
XG3390 XI11_6/XI0/XI0_32/d_4_ XI11_6/XI0/XI0_32/d__4_ DECAP_INV_G11
XG3391 XI11_6/XI0/XI0_32/d_3_ XI11_6/XI0/XI0_32/d__3_ DECAP_INV_G11
XG3392 XI11_6/XI0/XI0_32/d_2_ XI11_6/XI0/XI0_32/d__2_ DECAP_INV_G11
XG3393 XI11_6/XI0/XI0_32/d_1_ XI11_6/XI0/XI0_32/d__1_ DECAP_INV_G11
XG3394 XI11_6/XI0/XI0_32/d_0_ XI11_6/XI0/XI0_32/d__0_ DECAP_INV_G11
XG3395 XI11_6/XI0/XI0_31/d__15_ XI11_6/XI0/XI0_31/d_15_ DECAP_INV_G11
XG3396 XI11_6/XI0/XI0_31/d__14_ XI11_6/XI0/XI0_31/d_14_ DECAP_INV_G11
XG3397 XI11_6/XI0/XI0_31/d__13_ XI11_6/XI0/XI0_31/d_13_ DECAP_INV_G11
XG3398 XI11_6/XI0/XI0_31/d__12_ XI11_6/XI0/XI0_31/d_12_ DECAP_INV_G11
XG3399 XI11_6/XI0/XI0_31/d__11_ XI11_6/XI0/XI0_31/d_11_ DECAP_INV_G11
XG3400 XI11_6/XI0/XI0_31/d__10_ XI11_6/XI0/XI0_31/d_10_ DECAP_INV_G11
XG3401 XI11_6/XI0/XI0_31/d__9_ XI11_6/XI0/XI0_31/d_9_ DECAP_INV_G11
XG3402 XI11_6/XI0/XI0_31/d__8_ XI11_6/XI0/XI0_31/d_8_ DECAP_INV_G11
XG3403 XI11_6/XI0/XI0_31/d__7_ XI11_6/XI0/XI0_31/d_7_ DECAP_INV_G11
XG3404 XI11_6/XI0/XI0_31/d__6_ XI11_6/XI0/XI0_31/d_6_ DECAP_INV_G11
XG3405 XI11_6/XI0/XI0_31/d__5_ XI11_6/XI0/XI0_31/d_5_ DECAP_INV_G11
XG3406 XI11_6/XI0/XI0_31/d__4_ XI11_6/XI0/XI0_31/d_4_ DECAP_INV_G11
XG3407 XI11_6/XI0/XI0_31/d__3_ XI11_6/XI0/XI0_31/d_3_ DECAP_INV_G11
XG3408 XI11_6/XI0/XI0_31/d__2_ XI11_6/XI0/XI0_31/d_2_ DECAP_INV_G11
XG3409 XI11_6/XI0/XI0_31/d__1_ XI11_6/XI0/XI0_31/d_1_ DECAP_INV_G11
XG3410 XI11_6/XI0/XI0_31/d__0_ XI11_6/XI0/XI0_31/d_0_ DECAP_INV_G11
XG3411 XI11_6/XI0/XI0_31/d_15_ XI11_6/XI0/XI0_31/d__15_ DECAP_INV_G11
XG3412 XI11_6/XI0/XI0_31/d_14_ XI11_6/XI0/XI0_31/d__14_ DECAP_INV_G11
XG3413 XI11_6/XI0/XI0_31/d_13_ XI11_6/XI0/XI0_31/d__13_ DECAP_INV_G11
XG3414 XI11_6/XI0/XI0_31/d_12_ XI11_6/XI0/XI0_31/d__12_ DECAP_INV_G11
XG3415 XI11_6/XI0/XI0_31/d_11_ XI11_6/XI0/XI0_31/d__11_ DECAP_INV_G11
XG3416 XI11_6/XI0/XI0_31/d_10_ XI11_6/XI0/XI0_31/d__10_ DECAP_INV_G11
XG3417 XI11_6/XI0/XI0_31/d_9_ XI11_6/XI0/XI0_31/d__9_ DECAP_INV_G11
XG3418 XI11_6/XI0/XI0_31/d_8_ XI11_6/XI0/XI0_31/d__8_ DECAP_INV_G11
XG3419 XI11_6/XI0/XI0_31/d_7_ XI11_6/XI0/XI0_31/d__7_ DECAP_INV_G11
XG3420 XI11_6/XI0/XI0_31/d_6_ XI11_6/XI0/XI0_31/d__6_ DECAP_INV_G11
XG3421 XI11_6/XI0/XI0_31/d_5_ XI11_6/XI0/XI0_31/d__5_ DECAP_INV_G11
XG3422 XI11_6/XI0/XI0_31/d_4_ XI11_6/XI0/XI0_31/d__4_ DECAP_INV_G11
XG3423 XI11_6/XI0/XI0_31/d_3_ XI11_6/XI0/XI0_31/d__3_ DECAP_INV_G11
XG3424 XI11_6/XI0/XI0_31/d_2_ XI11_6/XI0/XI0_31/d__2_ DECAP_INV_G11
XG3425 XI11_6/XI0/XI0_31/d_1_ XI11_6/XI0/XI0_31/d__1_ DECAP_INV_G11
XG3426 XI11_6/XI0/XI0_31/d_0_ XI11_6/XI0/XI0_31/d__0_ DECAP_INV_G11
XG3427 XI11_6/XI0/XI0_30/d__15_ XI11_6/XI0/XI0_30/d_15_ DECAP_INV_G11
XG3428 XI11_6/XI0/XI0_30/d__14_ XI11_6/XI0/XI0_30/d_14_ DECAP_INV_G11
XG3429 XI11_6/XI0/XI0_30/d__13_ XI11_6/XI0/XI0_30/d_13_ DECAP_INV_G11
XG3430 XI11_6/XI0/XI0_30/d__12_ XI11_6/XI0/XI0_30/d_12_ DECAP_INV_G11
XG3431 XI11_6/XI0/XI0_30/d__11_ XI11_6/XI0/XI0_30/d_11_ DECAP_INV_G11
XG3432 XI11_6/XI0/XI0_30/d__10_ XI11_6/XI0/XI0_30/d_10_ DECAP_INV_G11
XG3433 XI11_6/XI0/XI0_30/d__9_ XI11_6/XI0/XI0_30/d_9_ DECAP_INV_G11
XG3434 XI11_6/XI0/XI0_30/d__8_ XI11_6/XI0/XI0_30/d_8_ DECAP_INV_G11
XG3435 XI11_6/XI0/XI0_30/d__7_ XI11_6/XI0/XI0_30/d_7_ DECAP_INV_G11
XG3436 XI11_6/XI0/XI0_30/d__6_ XI11_6/XI0/XI0_30/d_6_ DECAP_INV_G11
XG3437 XI11_6/XI0/XI0_30/d__5_ XI11_6/XI0/XI0_30/d_5_ DECAP_INV_G11
XG3438 XI11_6/XI0/XI0_30/d__4_ XI11_6/XI0/XI0_30/d_4_ DECAP_INV_G11
XG3439 XI11_6/XI0/XI0_30/d__3_ XI11_6/XI0/XI0_30/d_3_ DECAP_INV_G11
XG3440 XI11_6/XI0/XI0_30/d__2_ XI11_6/XI0/XI0_30/d_2_ DECAP_INV_G11
XG3441 XI11_6/XI0/XI0_30/d__1_ XI11_6/XI0/XI0_30/d_1_ DECAP_INV_G11
XG3442 XI11_6/XI0/XI0_30/d__0_ XI11_6/XI0/XI0_30/d_0_ DECAP_INV_G11
XG3443 XI11_6/XI0/XI0_30/d_15_ XI11_6/XI0/XI0_30/d__15_ DECAP_INV_G11
XG3444 XI11_6/XI0/XI0_30/d_14_ XI11_6/XI0/XI0_30/d__14_ DECAP_INV_G11
XG3445 XI11_6/XI0/XI0_30/d_13_ XI11_6/XI0/XI0_30/d__13_ DECAP_INV_G11
XG3446 XI11_6/XI0/XI0_30/d_12_ XI11_6/XI0/XI0_30/d__12_ DECAP_INV_G11
XG3447 XI11_6/XI0/XI0_30/d_11_ XI11_6/XI0/XI0_30/d__11_ DECAP_INV_G11
XG3448 XI11_6/XI0/XI0_30/d_10_ XI11_6/XI0/XI0_30/d__10_ DECAP_INV_G11
XG3449 XI11_6/XI0/XI0_30/d_9_ XI11_6/XI0/XI0_30/d__9_ DECAP_INV_G11
XG3450 XI11_6/XI0/XI0_30/d_8_ XI11_6/XI0/XI0_30/d__8_ DECAP_INV_G11
XG3451 XI11_6/XI0/XI0_30/d_7_ XI11_6/XI0/XI0_30/d__7_ DECAP_INV_G11
XG3452 XI11_6/XI0/XI0_30/d_6_ XI11_6/XI0/XI0_30/d__6_ DECAP_INV_G11
XG3453 XI11_6/XI0/XI0_30/d_5_ XI11_6/XI0/XI0_30/d__5_ DECAP_INV_G11
XG3454 XI11_6/XI0/XI0_30/d_4_ XI11_6/XI0/XI0_30/d__4_ DECAP_INV_G11
XG3455 XI11_6/XI0/XI0_30/d_3_ XI11_6/XI0/XI0_30/d__3_ DECAP_INV_G11
XG3456 XI11_6/XI0/XI0_30/d_2_ XI11_6/XI0/XI0_30/d__2_ DECAP_INV_G11
XG3457 XI11_6/XI0/XI0_30/d_1_ XI11_6/XI0/XI0_30/d__1_ DECAP_INV_G11
XG3458 XI11_6/XI0/XI0_30/d_0_ XI11_6/XI0/XI0_30/d__0_ DECAP_INV_G11
XG3459 XI11_6/XI0/XI0_29/d__15_ XI11_6/XI0/XI0_29/d_15_ DECAP_INV_G11
XG3460 XI11_6/XI0/XI0_29/d__14_ XI11_6/XI0/XI0_29/d_14_ DECAP_INV_G11
XG3461 XI11_6/XI0/XI0_29/d__13_ XI11_6/XI0/XI0_29/d_13_ DECAP_INV_G11
XG3462 XI11_6/XI0/XI0_29/d__12_ XI11_6/XI0/XI0_29/d_12_ DECAP_INV_G11
XG3463 XI11_6/XI0/XI0_29/d__11_ XI11_6/XI0/XI0_29/d_11_ DECAP_INV_G11
XG3464 XI11_6/XI0/XI0_29/d__10_ XI11_6/XI0/XI0_29/d_10_ DECAP_INV_G11
XG3465 XI11_6/XI0/XI0_29/d__9_ XI11_6/XI0/XI0_29/d_9_ DECAP_INV_G11
XG3466 XI11_6/XI0/XI0_29/d__8_ XI11_6/XI0/XI0_29/d_8_ DECAP_INV_G11
XG3467 XI11_6/XI0/XI0_29/d__7_ XI11_6/XI0/XI0_29/d_7_ DECAP_INV_G11
XG3468 XI11_6/XI0/XI0_29/d__6_ XI11_6/XI0/XI0_29/d_6_ DECAP_INV_G11
XG3469 XI11_6/XI0/XI0_29/d__5_ XI11_6/XI0/XI0_29/d_5_ DECAP_INV_G11
XG3470 XI11_6/XI0/XI0_29/d__4_ XI11_6/XI0/XI0_29/d_4_ DECAP_INV_G11
XG3471 XI11_6/XI0/XI0_29/d__3_ XI11_6/XI0/XI0_29/d_3_ DECAP_INV_G11
XG3472 XI11_6/XI0/XI0_29/d__2_ XI11_6/XI0/XI0_29/d_2_ DECAP_INV_G11
XG3473 XI11_6/XI0/XI0_29/d__1_ XI11_6/XI0/XI0_29/d_1_ DECAP_INV_G11
XG3474 XI11_6/XI0/XI0_29/d__0_ XI11_6/XI0/XI0_29/d_0_ DECAP_INV_G11
XG3475 XI11_6/XI0/XI0_29/d_15_ XI11_6/XI0/XI0_29/d__15_ DECAP_INV_G11
XG3476 XI11_6/XI0/XI0_29/d_14_ XI11_6/XI0/XI0_29/d__14_ DECAP_INV_G11
XG3477 XI11_6/XI0/XI0_29/d_13_ XI11_6/XI0/XI0_29/d__13_ DECAP_INV_G11
XG3478 XI11_6/XI0/XI0_29/d_12_ XI11_6/XI0/XI0_29/d__12_ DECAP_INV_G11
XG3479 XI11_6/XI0/XI0_29/d_11_ XI11_6/XI0/XI0_29/d__11_ DECAP_INV_G11
XG3480 XI11_6/XI0/XI0_29/d_10_ XI11_6/XI0/XI0_29/d__10_ DECAP_INV_G11
XG3481 XI11_6/XI0/XI0_29/d_9_ XI11_6/XI0/XI0_29/d__9_ DECAP_INV_G11
XG3482 XI11_6/XI0/XI0_29/d_8_ XI11_6/XI0/XI0_29/d__8_ DECAP_INV_G11
XG3483 XI11_6/XI0/XI0_29/d_7_ XI11_6/XI0/XI0_29/d__7_ DECAP_INV_G11
XG3484 XI11_6/XI0/XI0_29/d_6_ XI11_6/XI0/XI0_29/d__6_ DECAP_INV_G11
XG3485 XI11_6/XI0/XI0_29/d_5_ XI11_6/XI0/XI0_29/d__5_ DECAP_INV_G11
XG3486 XI11_6/XI0/XI0_29/d_4_ XI11_6/XI0/XI0_29/d__4_ DECAP_INV_G11
XG3487 XI11_6/XI0/XI0_29/d_3_ XI11_6/XI0/XI0_29/d__3_ DECAP_INV_G11
XG3488 XI11_6/XI0/XI0_29/d_2_ XI11_6/XI0/XI0_29/d__2_ DECAP_INV_G11
XG3489 XI11_6/XI0/XI0_29/d_1_ XI11_6/XI0/XI0_29/d__1_ DECAP_INV_G11
XG3490 XI11_6/XI0/XI0_29/d_0_ XI11_6/XI0/XI0_29/d__0_ DECAP_INV_G11
XG3491 XI11_6/XI0/XI0_28/d__15_ XI11_6/XI0/XI0_28/d_15_ DECAP_INV_G11
XG3492 XI11_6/XI0/XI0_28/d__14_ XI11_6/XI0/XI0_28/d_14_ DECAP_INV_G11
XG3493 XI11_6/XI0/XI0_28/d__13_ XI11_6/XI0/XI0_28/d_13_ DECAP_INV_G11
XG3494 XI11_6/XI0/XI0_28/d__12_ XI11_6/XI0/XI0_28/d_12_ DECAP_INV_G11
XG3495 XI11_6/XI0/XI0_28/d__11_ XI11_6/XI0/XI0_28/d_11_ DECAP_INV_G11
XG3496 XI11_6/XI0/XI0_28/d__10_ XI11_6/XI0/XI0_28/d_10_ DECAP_INV_G11
XG3497 XI11_6/XI0/XI0_28/d__9_ XI11_6/XI0/XI0_28/d_9_ DECAP_INV_G11
XG3498 XI11_6/XI0/XI0_28/d__8_ XI11_6/XI0/XI0_28/d_8_ DECAP_INV_G11
XG3499 XI11_6/XI0/XI0_28/d__7_ XI11_6/XI0/XI0_28/d_7_ DECAP_INV_G11
XG3500 XI11_6/XI0/XI0_28/d__6_ XI11_6/XI0/XI0_28/d_6_ DECAP_INV_G11
XG3501 XI11_6/XI0/XI0_28/d__5_ XI11_6/XI0/XI0_28/d_5_ DECAP_INV_G11
XG3502 XI11_6/XI0/XI0_28/d__4_ XI11_6/XI0/XI0_28/d_4_ DECAP_INV_G11
XG3503 XI11_6/XI0/XI0_28/d__3_ XI11_6/XI0/XI0_28/d_3_ DECAP_INV_G11
XG3504 XI11_6/XI0/XI0_28/d__2_ XI11_6/XI0/XI0_28/d_2_ DECAP_INV_G11
XG3505 XI11_6/XI0/XI0_28/d__1_ XI11_6/XI0/XI0_28/d_1_ DECAP_INV_G11
XG3506 XI11_6/XI0/XI0_28/d__0_ XI11_6/XI0/XI0_28/d_0_ DECAP_INV_G11
XG3507 XI11_6/XI0/XI0_28/d_15_ XI11_6/XI0/XI0_28/d__15_ DECAP_INV_G11
XG3508 XI11_6/XI0/XI0_28/d_14_ XI11_6/XI0/XI0_28/d__14_ DECAP_INV_G11
XG3509 XI11_6/XI0/XI0_28/d_13_ XI11_6/XI0/XI0_28/d__13_ DECAP_INV_G11
XG3510 XI11_6/XI0/XI0_28/d_12_ XI11_6/XI0/XI0_28/d__12_ DECAP_INV_G11
XG3511 XI11_6/XI0/XI0_28/d_11_ XI11_6/XI0/XI0_28/d__11_ DECAP_INV_G11
XG3512 XI11_6/XI0/XI0_28/d_10_ XI11_6/XI0/XI0_28/d__10_ DECAP_INV_G11
XG3513 XI11_6/XI0/XI0_28/d_9_ XI11_6/XI0/XI0_28/d__9_ DECAP_INV_G11
XG3514 XI11_6/XI0/XI0_28/d_8_ XI11_6/XI0/XI0_28/d__8_ DECAP_INV_G11
XG3515 XI11_6/XI0/XI0_28/d_7_ XI11_6/XI0/XI0_28/d__7_ DECAP_INV_G11
XG3516 XI11_6/XI0/XI0_28/d_6_ XI11_6/XI0/XI0_28/d__6_ DECAP_INV_G11
XG3517 XI11_6/XI0/XI0_28/d_5_ XI11_6/XI0/XI0_28/d__5_ DECAP_INV_G11
XG3518 XI11_6/XI0/XI0_28/d_4_ XI11_6/XI0/XI0_28/d__4_ DECAP_INV_G11
XG3519 XI11_6/XI0/XI0_28/d_3_ XI11_6/XI0/XI0_28/d__3_ DECAP_INV_G11
XG3520 XI11_6/XI0/XI0_28/d_2_ XI11_6/XI0/XI0_28/d__2_ DECAP_INV_G11
XG3521 XI11_6/XI0/XI0_28/d_1_ XI11_6/XI0/XI0_28/d__1_ DECAP_INV_G11
XG3522 XI11_6/XI0/XI0_28/d_0_ XI11_6/XI0/XI0_28/d__0_ DECAP_INV_G11
XG3523 XI11_6/XI0/XI0_27/d__15_ XI11_6/XI0/XI0_27/d_15_ DECAP_INV_G11
XG3524 XI11_6/XI0/XI0_27/d__14_ XI11_6/XI0/XI0_27/d_14_ DECAP_INV_G11
XG3525 XI11_6/XI0/XI0_27/d__13_ XI11_6/XI0/XI0_27/d_13_ DECAP_INV_G11
XG3526 XI11_6/XI0/XI0_27/d__12_ XI11_6/XI0/XI0_27/d_12_ DECAP_INV_G11
XG3527 XI11_6/XI0/XI0_27/d__11_ XI11_6/XI0/XI0_27/d_11_ DECAP_INV_G11
XG3528 XI11_6/XI0/XI0_27/d__10_ XI11_6/XI0/XI0_27/d_10_ DECAP_INV_G11
XG3529 XI11_6/XI0/XI0_27/d__9_ XI11_6/XI0/XI0_27/d_9_ DECAP_INV_G11
XG3530 XI11_6/XI0/XI0_27/d__8_ XI11_6/XI0/XI0_27/d_8_ DECAP_INV_G11
XG3531 XI11_6/XI0/XI0_27/d__7_ XI11_6/XI0/XI0_27/d_7_ DECAP_INV_G11
XG3532 XI11_6/XI0/XI0_27/d__6_ XI11_6/XI0/XI0_27/d_6_ DECAP_INV_G11
XG3533 XI11_6/XI0/XI0_27/d__5_ XI11_6/XI0/XI0_27/d_5_ DECAP_INV_G11
XG3534 XI11_6/XI0/XI0_27/d__4_ XI11_6/XI0/XI0_27/d_4_ DECAP_INV_G11
XG3535 XI11_6/XI0/XI0_27/d__3_ XI11_6/XI0/XI0_27/d_3_ DECAP_INV_G11
XG3536 XI11_6/XI0/XI0_27/d__2_ XI11_6/XI0/XI0_27/d_2_ DECAP_INV_G11
XG3537 XI11_6/XI0/XI0_27/d__1_ XI11_6/XI0/XI0_27/d_1_ DECAP_INV_G11
XG3538 XI11_6/XI0/XI0_27/d__0_ XI11_6/XI0/XI0_27/d_0_ DECAP_INV_G11
XG3539 XI11_6/XI0/XI0_27/d_15_ XI11_6/XI0/XI0_27/d__15_ DECAP_INV_G11
XG3540 XI11_6/XI0/XI0_27/d_14_ XI11_6/XI0/XI0_27/d__14_ DECAP_INV_G11
XG3541 XI11_6/XI0/XI0_27/d_13_ XI11_6/XI0/XI0_27/d__13_ DECAP_INV_G11
XG3542 XI11_6/XI0/XI0_27/d_12_ XI11_6/XI0/XI0_27/d__12_ DECAP_INV_G11
XG3543 XI11_6/XI0/XI0_27/d_11_ XI11_6/XI0/XI0_27/d__11_ DECAP_INV_G11
XG3544 XI11_6/XI0/XI0_27/d_10_ XI11_6/XI0/XI0_27/d__10_ DECAP_INV_G11
XG3545 XI11_6/XI0/XI0_27/d_9_ XI11_6/XI0/XI0_27/d__9_ DECAP_INV_G11
XG3546 XI11_6/XI0/XI0_27/d_8_ XI11_6/XI0/XI0_27/d__8_ DECAP_INV_G11
XG3547 XI11_6/XI0/XI0_27/d_7_ XI11_6/XI0/XI0_27/d__7_ DECAP_INV_G11
XG3548 XI11_6/XI0/XI0_27/d_6_ XI11_6/XI0/XI0_27/d__6_ DECAP_INV_G11
XG3549 XI11_6/XI0/XI0_27/d_5_ XI11_6/XI0/XI0_27/d__5_ DECAP_INV_G11
XG3550 XI11_6/XI0/XI0_27/d_4_ XI11_6/XI0/XI0_27/d__4_ DECAP_INV_G11
XG3551 XI11_6/XI0/XI0_27/d_3_ XI11_6/XI0/XI0_27/d__3_ DECAP_INV_G11
XG3552 XI11_6/XI0/XI0_27/d_2_ XI11_6/XI0/XI0_27/d__2_ DECAP_INV_G11
XG3553 XI11_6/XI0/XI0_27/d_1_ XI11_6/XI0/XI0_27/d__1_ DECAP_INV_G11
XG3554 XI11_6/XI0/XI0_27/d_0_ XI11_6/XI0/XI0_27/d__0_ DECAP_INV_G11
XG3555 XI11_6/XI0/XI0_26/d__15_ XI11_6/XI0/XI0_26/d_15_ DECAP_INV_G11
XG3556 XI11_6/XI0/XI0_26/d__14_ XI11_6/XI0/XI0_26/d_14_ DECAP_INV_G11
XG3557 XI11_6/XI0/XI0_26/d__13_ XI11_6/XI0/XI0_26/d_13_ DECAP_INV_G11
XG3558 XI11_6/XI0/XI0_26/d__12_ XI11_6/XI0/XI0_26/d_12_ DECAP_INV_G11
XG3559 XI11_6/XI0/XI0_26/d__11_ XI11_6/XI0/XI0_26/d_11_ DECAP_INV_G11
XG3560 XI11_6/XI0/XI0_26/d__10_ XI11_6/XI0/XI0_26/d_10_ DECAP_INV_G11
XG3561 XI11_6/XI0/XI0_26/d__9_ XI11_6/XI0/XI0_26/d_9_ DECAP_INV_G11
XG3562 XI11_6/XI0/XI0_26/d__8_ XI11_6/XI0/XI0_26/d_8_ DECAP_INV_G11
XG3563 XI11_6/XI0/XI0_26/d__7_ XI11_6/XI0/XI0_26/d_7_ DECAP_INV_G11
XG3564 XI11_6/XI0/XI0_26/d__6_ XI11_6/XI0/XI0_26/d_6_ DECAP_INV_G11
XG3565 XI11_6/XI0/XI0_26/d__5_ XI11_6/XI0/XI0_26/d_5_ DECAP_INV_G11
XG3566 XI11_6/XI0/XI0_26/d__4_ XI11_6/XI0/XI0_26/d_4_ DECAP_INV_G11
XG3567 XI11_6/XI0/XI0_26/d__3_ XI11_6/XI0/XI0_26/d_3_ DECAP_INV_G11
XG3568 XI11_6/XI0/XI0_26/d__2_ XI11_6/XI0/XI0_26/d_2_ DECAP_INV_G11
XG3569 XI11_6/XI0/XI0_26/d__1_ XI11_6/XI0/XI0_26/d_1_ DECAP_INV_G11
XG3570 XI11_6/XI0/XI0_26/d__0_ XI11_6/XI0/XI0_26/d_0_ DECAP_INV_G11
XG3571 XI11_6/XI0/XI0_26/d_15_ XI11_6/XI0/XI0_26/d__15_ DECAP_INV_G11
XG3572 XI11_6/XI0/XI0_26/d_14_ XI11_6/XI0/XI0_26/d__14_ DECAP_INV_G11
XG3573 XI11_6/XI0/XI0_26/d_13_ XI11_6/XI0/XI0_26/d__13_ DECAP_INV_G11
XG3574 XI11_6/XI0/XI0_26/d_12_ XI11_6/XI0/XI0_26/d__12_ DECAP_INV_G11
XG3575 XI11_6/XI0/XI0_26/d_11_ XI11_6/XI0/XI0_26/d__11_ DECAP_INV_G11
XG3576 XI11_6/XI0/XI0_26/d_10_ XI11_6/XI0/XI0_26/d__10_ DECAP_INV_G11
XG3577 XI11_6/XI0/XI0_26/d_9_ XI11_6/XI0/XI0_26/d__9_ DECAP_INV_G11
XG3578 XI11_6/XI0/XI0_26/d_8_ XI11_6/XI0/XI0_26/d__8_ DECAP_INV_G11
XG3579 XI11_6/XI0/XI0_26/d_7_ XI11_6/XI0/XI0_26/d__7_ DECAP_INV_G11
XG3580 XI11_6/XI0/XI0_26/d_6_ XI11_6/XI0/XI0_26/d__6_ DECAP_INV_G11
XG3581 XI11_6/XI0/XI0_26/d_5_ XI11_6/XI0/XI0_26/d__5_ DECAP_INV_G11
XG3582 XI11_6/XI0/XI0_26/d_4_ XI11_6/XI0/XI0_26/d__4_ DECAP_INV_G11
XG3583 XI11_6/XI0/XI0_26/d_3_ XI11_6/XI0/XI0_26/d__3_ DECAP_INV_G11
XG3584 XI11_6/XI0/XI0_26/d_2_ XI11_6/XI0/XI0_26/d__2_ DECAP_INV_G11
XG3585 XI11_6/XI0/XI0_26/d_1_ XI11_6/XI0/XI0_26/d__1_ DECAP_INV_G11
XG3586 XI11_6/XI0/XI0_26/d_0_ XI11_6/XI0/XI0_26/d__0_ DECAP_INV_G11
XG3587 XI11_6/XI0/XI0_25/d__15_ XI11_6/XI0/XI0_25/d_15_ DECAP_INV_G11
XG3588 XI11_6/XI0/XI0_25/d__14_ XI11_6/XI0/XI0_25/d_14_ DECAP_INV_G11
XG3589 XI11_6/XI0/XI0_25/d__13_ XI11_6/XI0/XI0_25/d_13_ DECAP_INV_G11
XG3590 XI11_6/XI0/XI0_25/d__12_ XI11_6/XI0/XI0_25/d_12_ DECAP_INV_G11
XG3591 XI11_6/XI0/XI0_25/d__11_ XI11_6/XI0/XI0_25/d_11_ DECAP_INV_G11
XG3592 XI11_6/XI0/XI0_25/d__10_ XI11_6/XI0/XI0_25/d_10_ DECAP_INV_G11
XG3593 XI11_6/XI0/XI0_25/d__9_ XI11_6/XI0/XI0_25/d_9_ DECAP_INV_G11
XG3594 XI11_6/XI0/XI0_25/d__8_ XI11_6/XI0/XI0_25/d_8_ DECAP_INV_G11
XG3595 XI11_6/XI0/XI0_25/d__7_ XI11_6/XI0/XI0_25/d_7_ DECAP_INV_G11
XG3596 XI11_6/XI0/XI0_25/d__6_ XI11_6/XI0/XI0_25/d_6_ DECAP_INV_G11
XG3597 XI11_6/XI0/XI0_25/d__5_ XI11_6/XI0/XI0_25/d_5_ DECAP_INV_G11
XG3598 XI11_6/XI0/XI0_25/d__4_ XI11_6/XI0/XI0_25/d_4_ DECAP_INV_G11
XG3599 XI11_6/XI0/XI0_25/d__3_ XI11_6/XI0/XI0_25/d_3_ DECAP_INV_G11
XG3600 XI11_6/XI0/XI0_25/d__2_ XI11_6/XI0/XI0_25/d_2_ DECAP_INV_G11
XG3601 XI11_6/XI0/XI0_25/d__1_ XI11_6/XI0/XI0_25/d_1_ DECAP_INV_G11
XG3602 XI11_6/XI0/XI0_25/d__0_ XI11_6/XI0/XI0_25/d_0_ DECAP_INV_G11
XG3603 XI11_6/XI0/XI0_25/d_15_ XI11_6/XI0/XI0_25/d__15_ DECAP_INV_G11
XG3604 XI11_6/XI0/XI0_25/d_14_ XI11_6/XI0/XI0_25/d__14_ DECAP_INV_G11
XG3605 XI11_6/XI0/XI0_25/d_13_ XI11_6/XI0/XI0_25/d__13_ DECAP_INV_G11
XG3606 XI11_6/XI0/XI0_25/d_12_ XI11_6/XI0/XI0_25/d__12_ DECAP_INV_G11
XG3607 XI11_6/XI0/XI0_25/d_11_ XI11_6/XI0/XI0_25/d__11_ DECAP_INV_G11
XG3608 XI11_6/XI0/XI0_25/d_10_ XI11_6/XI0/XI0_25/d__10_ DECAP_INV_G11
XG3609 XI11_6/XI0/XI0_25/d_9_ XI11_6/XI0/XI0_25/d__9_ DECAP_INV_G11
XG3610 XI11_6/XI0/XI0_25/d_8_ XI11_6/XI0/XI0_25/d__8_ DECAP_INV_G11
XG3611 XI11_6/XI0/XI0_25/d_7_ XI11_6/XI0/XI0_25/d__7_ DECAP_INV_G11
XG3612 XI11_6/XI0/XI0_25/d_6_ XI11_6/XI0/XI0_25/d__6_ DECAP_INV_G11
XG3613 XI11_6/XI0/XI0_25/d_5_ XI11_6/XI0/XI0_25/d__5_ DECAP_INV_G11
XG3614 XI11_6/XI0/XI0_25/d_4_ XI11_6/XI0/XI0_25/d__4_ DECAP_INV_G11
XG3615 XI11_6/XI0/XI0_25/d_3_ XI11_6/XI0/XI0_25/d__3_ DECAP_INV_G11
XG3616 XI11_6/XI0/XI0_25/d_2_ XI11_6/XI0/XI0_25/d__2_ DECAP_INV_G11
XG3617 XI11_6/XI0/XI0_25/d_1_ XI11_6/XI0/XI0_25/d__1_ DECAP_INV_G11
XG3618 XI11_6/XI0/XI0_25/d_0_ XI11_6/XI0/XI0_25/d__0_ DECAP_INV_G11
XG3619 XI11_6/XI0/XI0_24/d__15_ XI11_6/XI0/XI0_24/d_15_ DECAP_INV_G11
XG3620 XI11_6/XI0/XI0_24/d__14_ XI11_6/XI0/XI0_24/d_14_ DECAP_INV_G11
XG3621 XI11_6/XI0/XI0_24/d__13_ XI11_6/XI0/XI0_24/d_13_ DECAP_INV_G11
XG3622 XI11_6/XI0/XI0_24/d__12_ XI11_6/XI0/XI0_24/d_12_ DECAP_INV_G11
XG3623 XI11_6/XI0/XI0_24/d__11_ XI11_6/XI0/XI0_24/d_11_ DECAP_INV_G11
XG3624 XI11_6/XI0/XI0_24/d__10_ XI11_6/XI0/XI0_24/d_10_ DECAP_INV_G11
XG3625 XI11_6/XI0/XI0_24/d__9_ XI11_6/XI0/XI0_24/d_9_ DECAP_INV_G11
XG3626 XI11_6/XI0/XI0_24/d__8_ XI11_6/XI0/XI0_24/d_8_ DECAP_INV_G11
XG3627 XI11_6/XI0/XI0_24/d__7_ XI11_6/XI0/XI0_24/d_7_ DECAP_INV_G11
XG3628 XI11_6/XI0/XI0_24/d__6_ XI11_6/XI0/XI0_24/d_6_ DECAP_INV_G11
XG3629 XI11_6/XI0/XI0_24/d__5_ XI11_6/XI0/XI0_24/d_5_ DECAP_INV_G11
XG3630 XI11_6/XI0/XI0_24/d__4_ XI11_6/XI0/XI0_24/d_4_ DECAP_INV_G11
XG3631 XI11_6/XI0/XI0_24/d__3_ XI11_6/XI0/XI0_24/d_3_ DECAP_INV_G11
XG3632 XI11_6/XI0/XI0_24/d__2_ XI11_6/XI0/XI0_24/d_2_ DECAP_INV_G11
XG3633 XI11_6/XI0/XI0_24/d__1_ XI11_6/XI0/XI0_24/d_1_ DECAP_INV_G11
XG3634 XI11_6/XI0/XI0_24/d__0_ XI11_6/XI0/XI0_24/d_0_ DECAP_INV_G11
XG3635 XI11_6/XI0/XI0_24/d_15_ XI11_6/XI0/XI0_24/d__15_ DECAP_INV_G11
XG3636 XI11_6/XI0/XI0_24/d_14_ XI11_6/XI0/XI0_24/d__14_ DECAP_INV_G11
XG3637 XI11_6/XI0/XI0_24/d_13_ XI11_6/XI0/XI0_24/d__13_ DECAP_INV_G11
XG3638 XI11_6/XI0/XI0_24/d_12_ XI11_6/XI0/XI0_24/d__12_ DECAP_INV_G11
XG3639 XI11_6/XI0/XI0_24/d_11_ XI11_6/XI0/XI0_24/d__11_ DECAP_INV_G11
XG3640 XI11_6/XI0/XI0_24/d_10_ XI11_6/XI0/XI0_24/d__10_ DECAP_INV_G11
XG3641 XI11_6/XI0/XI0_24/d_9_ XI11_6/XI0/XI0_24/d__9_ DECAP_INV_G11
XG3642 XI11_6/XI0/XI0_24/d_8_ XI11_6/XI0/XI0_24/d__8_ DECAP_INV_G11
XG3643 XI11_6/XI0/XI0_24/d_7_ XI11_6/XI0/XI0_24/d__7_ DECAP_INV_G11
XG3644 XI11_6/XI0/XI0_24/d_6_ XI11_6/XI0/XI0_24/d__6_ DECAP_INV_G11
XG3645 XI11_6/XI0/XI0_24/d_5_ XI11_6/XI0/XI0_24/d__5_ DECAP_INV_G11
XG3646 XI11_6/XI0/XI0_24/d_4_ XI11_6/XI0/XI0_24/d__4_ DECAP_INV_G11
XG3647 XI11_6/XI0/XI0_24/d_3_ XI11_6/XI0/XI0_24/d__3_ DECAP_INV_G11
XG3648 XI11_6/XI0/XI0_24/d_2_ XI11_6/XI0/XI0_24/d__2_ DECAP_INV_G11
XG3649 XI11_6/XI0/XI0_24/d_1_ XI11_6/XI0/XI0_24/d__1_ DECAP_INV_G11
XG3650 XI11_6/XI0/XI0_24/d_0_ XI11_6/XI0/XI0_24/d__0_ DECAP_INV_G11
XG3651 XI11_6/XI0/XI0_23/d__15_ XI11_6/XI0/XI0_23/d_15_ DECAP_INV_G11
XG3652 XI11_6/XI0/XI0_23/d__14_ XI11_6/XI0/XI0_23/d_14_ DECAP_INV_G11
XG3653 XI11_6/XI0/XI0_23/d__13_ XI11_6/XI0/XI0_23/d_13_ DECAP_INV_G11
XG3654 XI11_6/XI0/XI0_23/d__12_ XI11_6/XI0/XI0_23/d_12_ DECAP_INV_G11
XG3655 XI11_6/XI0/XI0_23/d__11_ XI11_6/XI0/XI0_23/d_11_ DECAP_INV_G11
XG3656 XI11_6/XI0/XI0_23/d__10_ XI11_6/XI0/XI0_23/d_10_ DECAP_INV_G11
XG3657 XI11_6/XI0/XI0_23/d__9_ XI11_6/XI0/XI0_23/d_9_ DECAP_INV_G11
XG3658 XI11_6/XI0/XI0_23/d__8_ XI11_6/XI0/XI0_23/d_8_ DECAP_INV_G11
XG3659 XI11_6/XI0/XI0_23/d__7_ XI11_6/XI0/XI0_23/d_7_ DECAP_INV_G11
XG3660 XI11_6/XI0/XI0_23/d__6_ XI11_6/XI0/XI0_23/d_6_ DECAP_INV_G11
XG3661 XI11_6/XI0/XI0_23/d__5_ XI11_6/XI0/XI0_23/d_5_ DECAP_INV_G11
XG3662 XI11_6/XI0/XI0_23/d__4_ XI11_6/XI0/XI0_23/d_4_ DECAP_INV_G11
XG3663 XI11_6/XI0/XI0_23/d__3_ XI11_6/XI0/XI0_23/d_3_ DECAP_INV_G11
XG3664 XI11_6/XI0/XI0_23/d__2_ XI11_6/XI0/XI0_23/d_2_ DECAP_INV_G11
XG3665 XI11_6/XI0/XI0_23/d__1_ XI11_6/XI0/XI0_23/d_1_ DECAP_INV_G11
XG3666 XI11_6/XI0/XI0_23/d__0_ XI11_6/XI0/XI0_23/d_0_ DECAP_INV_G11
XG3667 XI11_6/XI0/XI0_23/d_15_ XI11_6/XI0/XI0_23/d__15_ DECAP_INV_G11
XG3668 XI11_6/XI0/XI0_23/d_14_ XI11_6/XI0/XI0_23/d__14_ DECAP_INV_G11
XG3669 XI11_6/XI0/XI0_23/d_13_ XI11_6/XI0/XI0_23/d__13_ DECAP_INV_G11
XG3670 XI11_6/XI0/XI0_23/d_12_ XI11_6/XI0/XI0_23/d__12_ DECAP_INV_G11
XG3671 XI11_6/XI0/XI0_23/d_11_ XI11_6/XI0/XI0_23/d__11_ DECAP_INV_G11
XG3672 XI11_6/XI0/XI0_23/d_10_ XI11_6/XI0/XI0_23/d__10_ DECAP_INV_G11
XG3673 XI11_6/XI0/XI0_23/d_9_ XI11_6/XI0/XI0_23/d__9_ DECAP_INV_G11
XG3674 XI11_6/XI0/XI0_23/d_8_ XI11_6/XI0/XI0_23/d__8_ DECAP_INV_G11
XG3675 XI11_6/XI0/XI0_23/d_7_ XI11_6/XI0/XI0_23/d__7_ DECAP_INV_G11
XG3676 XI11_6/XI0/XI0_23/d_6_ XI11_6/XI0/XI0_23/d__6_ DECAP_INV_G11
XG3677 XI11_6/XI0/XI0_23/d_5_ XI11_6/XI0/XI0_23/d__5_ DECAP_INV_G11
XG3678 XI11_6/XI0/XI0_23/d_4_ XI11_6/XI0/XI0_23/d__4_ DECAP_INV_G11
XG3679 XI11_6/XI0/XI0_23/d_3_ XI11_6/XI0/XI0_23/d__3_ DECAP_INV_G11
XG3680 XI11_6/XI0/XI0_23/d_2_ XI11_6/XI0/XI0_23/d__2_ DECAP_INV_G11
XG3681 XI11_6/XI0/XI0_23/d_1_ XI11_6/XI0/XI0_23/d__1_ DECAP_INV_G11
XG3682 XI11_6/XI0/XI0_23/d_0_ XI11_6/XI0/XI0_23/d__0_ DECAP_INV_G11
XG3683 XI11_6/XI0/XI0_22/d__15_ XI11_6/XI0/XI0_22/d_15_ DECAP_INV_G11
XG3684 XI11_6/XI0/XI0_22/d__14_ XI11_6/XI0/XI0_22/d_14_ DECAP_INV_G11
XG3685 XI11_6/XI0/XI0_22/d__13_ XI11_6/XI0/XI0_22/d_13_ DECAP_INV_G11
XG3686 XI11_6/XI0/XI0_22/d__12_ XI11_6/XI0/XI0_22/d_12_ DECAP_INV_G11
XG3687 XI11_6/XI0/XI0_22/d__11_ XI11_6/XI0/XI0_22/d_11_ DECAP_INV_G11
XG3688 XI11_6/XI0/XI0_22/d__10_ XI11_6/XI0/XI0_22/d_10_ DECAP_INV_G11
XG3689 XI11_6/XI0/XI0_22/d__9_ XI11_6/XI0/XI0_22/d_9_ DECAP_INV_G11
XG3690 XI11_6/XI0/XI0_22/d__8_ XI11_6/XI0/XI0_22/d_8_ DECAP_INV_G11
XG3691 XI11_6/XI0/XI0_22/d__7_ XI11_6/XI0/XI0_22/d_7_ DECAP_INV_G11
XG3692 XI11_6/XI0/XI0_22/d__6_ XI11_6/XI0/XI0_22/d_6_ DECAP_INV_G11
XG3693 XI11_6/XI0/XI0_22/d__5_ XI11_6/XI0/XI0_22/d_5_ DECAP_INV_G11
XG3694 XI11_6/XI0/XI0_22/d__4_ XI11_6/XI0/XI0_22/d_4_ DECAP_INV_G11
XG3695 XI11_6/XI0/XI0_22/d__3_ XI11_6/XI0/XI0_22/d_3_ DECAP_INV_G11
XG3696 XI11_6/XI0/XI0_22/d__2_ XI11_6/XI0/XI0_22/d_2_ DECAP_INV_G11
XG3697 XI11_6/XI0/XI0_22/d__1_ XI11_6/XI0/XI0_22/d_1_ DECAP_INV_G11
XG3698 XI11_6/XI0/XI0_22/d__0_ XI11_6/XI0/XI0_22/d_0_ DECAP_INV_G11
XG3699 XI11_6/XI0/XI0_22/d_15_ XI11_6/XI0/XI0_22/d__15_ DECAP_INV_G11
XG3700 XI11_6/XI0/XI0_22/d_14_ XI11_6/XI0/XI0_22/d__14_ DECAP_INV_G11
XG3701 XI11_6/XI0/XI0_22/d_13_ XI11_6/XI0/XI0_22/d__13_ DECAP_INV_G11
XG3702 XI11_6/XI0/XI0_22/d_12_ XI11_6/XI0/XI0_22/d__12_ DECAP_INV_G11
XG3703 XI11_6/XI0/XI0_22/d_11_ XI11_6/XI0/XI0_22/d__11_ DECAP_INV_G11
XG3704 XI11_6/XI0/XI0_22/d_10_ XI11_6/XI0/XI0_22/d__10_ DECAP_INV_G11
XG3705 XI11_6/XI0/XI0_22/d_9_ XI11_6/XI0/XI0_22/d__9_ DECAP_INV_G11
XG3706 XI11_6/XI0/XI0_22/d_8_ XI11_6/XI0/XI0_22/d__8_ DECAP_INV_G11
XG3707 XI11_6/XI0/XI0_22/d_7_ XI11_6/XI0/XI0_22/d__7_ DECAP_INV_G11
XG3708 XI11_6/XI0/XI0_22/d_6_ XI11_6/XI0/XI0_22/d__6_ DECAP_INV_G11
XG3709 XI11_6/XI0/XI0_22/d_5_ XI11_6/XI0/XI0_22/d__5_ DECAP_INV_G11
XG3710 XI11_6/XI0/XI0_22/d_4_ XI11_6/XI0/XI0_22/d__4_ DECAP_INV_G11
XG3711 XI11_6/XI0/XI0_22/d_3_ XI11_6/XI0/XI0_22/d__3_ DECAP_INV_G11
XG3712 XI11_6/XI0/XI0_22/d_2_ XI11_6/XI0/XI0_22/d__2_ DECAP_INV_G11
XG3713 XI11_6/XI0/XI0_22/d_1_ XI11_6/XI0/XI0_22/d__1_ DECAP_INV_G11
XG3714 XI11_6/XI0/XI0_22/d_0_ XI11_6/XI0/XI0_22/d__0_ DECAP_INV_G11
XG3715 XI11_6/XI0/XI0_21/d__15_ XI11_6/XI0/XI0_21/d_15_ DECAP_INV_G11
XG3716 XI11_6/XI0/XI0_21/d__14_ XI11_6/XI0/XI0_21/d_14_ DECAP_INV_G11
XG3717 XI11_6/XI0/XI0_21/d__13_ XI11_6/XI0/XI0_21/d_13_ DECAP_INV_G11
XG3718 XI11_6/XI0/XI0_21/d__12_ XI11_6/XI0/XI0_21/d_12_ DECAP_INV_G11
XG3719 XI11_6/XI0/XI0_21/d__11_ XI11_6/XI0/XI0_21/d_11_ DECAP_INV_G11
XG3720 XI11_6/XI0/XI0_21/d__10_ XI11_6/XI0/XI0_21/d_10_ DECAP_INV_G11
XG3721 XI11_6/XI0/XI0_21/d__9_ XI11_6/XI0/XI0_21/d_9_ DECAP_INV_G11
XG3722 XI11_6/XI0/XI0_21/d__8_ XI11_6/XI0/XI0_21/d_8_ DECAP_INV_G11
XG3723 XI11_6/XI0/XI0_21/d__7_ XI11_6/XI0/XI0_21/d_7_ DECAP_INV_G11
XG3724 XI11_6/XI0/XI0_21/d__6_ XI11_6/XI0/XI0_21/d_6_ DECAP_INV_G11
XG3725 XI11_6/XI0/XI0_21/d__5_ XI11_6/XI0/XI0_21/d_5_ DECAP_INV_G11
XG3726 XI11_6/XI0/XI0_21/d__4_ XI11_6/XI0/XI0_21/d_4_ DECAP_INV_G11
XG3727 XI11_6/XI0/XI0_21/d__3_ XI11_6/XI0/XI0_21/d_3_ DECAP_INV_G11
XG3728 XI11_6/XI0/XI0_21/d__2_ XI11_6/XI0/XI0_21/d_2_ DECAP_INV_G11
XG3729 XI11_6/XI0/XI0_21/d__1_ XI11_6/XI0/XI0_21/d_1_ DECAP_INV_G11
XG3730 XI11_6/XI0/XI0_21/d__0_ XI11_6/XI0/XI0_21/d_0_ DECAP_INV_G11
XG3731 XI11_6/XI0/XI0_21/d_15_ XI11_6/XI0/XI0_21/d__15_ DECAP_INV_G11
XG3732 XI11_6/XI0/XI0_21/d_14_ XI11_6/XI0/XI0_21/d__14_ DECAP_INV_G11
XG3733 XI11_6/XI0/XI0_21/d_13_ XI11_6/XI0/XI0_21/d__13_ DECAP_INV_G11
XG3734 XI11_6/XI0/XI0_21/d_12_ XI11_6/XI0/XI0_21/d__12_ DECAP_INV_G11
XG3735 XI11_6/XI0/XI0_21/d_11_ XI11_6/XI0/XI0_21/d__11_ DECAP_INV_G11
XG3736 XI11_6/XI0/XI0_21/d_10_ XI11_6/XI0/XI0_21/d__10_ DECAP_INV_G11
XG3737 XI11_6/XI0/XI0_21/d_9_ XI11_6/XI0/XI0_21/d__9_ DECAP_INV_G11
XG3738 XI11_6/XI0/XI0_21/d_8_ XI11_6/XI0/XI0_21/d__8_ DECAP_INV_G11
XG3739 XI11_6/XI0/XI0_21/d_7_ XI11_6/XI0/XI0_21/d__7_ DECAP_INV_G11
XG3740 XI11_6/XI0/XI0_21/d_6_ XI11_6/XI0/XI0_21/d__6_ DECAP_INV_G11
XG3741 XI11_6/XI0/XI0_21/d_5_ XI11_6/XI0/XI0_21/d__5_ DECAP_INV_G11
XG3742 XI11_6/XI0/XI0_21/d_4_ XI11_6/XI0/XI0_21/d__4_ DECAP_INV_G11
XG3743 XI11_6/XI0/XI0_21/d_3_ XI11_6/XI0/XI0_21/d__3_ DECAP_INV_G11
XG3744 XI11_6/XI0/XI0_21/d_2_ XI11_6/XI0/XI0_21/d__2_ DECAP_INV_G11
XG3745 XI11_6/XI0/XI0_21/d_1_ XI11_6/XI0/XI0_21/d__1_ DECAP_INV_G11
XG3746 XI11_6/XI0/XI0_21/d_0_ XI11_6/XI0/XI0_21/d__0_ DECAP_INV_G11
XG3747 XI11_6/XI0/XI0_20/d__15_ XI11_6/XI0/XI0_20/d_15_ DECAP_INV_G11
XG3748 XI11_6/XI0/XI0_20/d__14_ XI11_6/XI0/XI0_20/d_14_ DECAP_INV_G11
XG3749 XI11_6/XI0/XI0_20/d__13_ XI11_6/XI0/XI0_20/d_13_ DECAP_INV_G11
XG3750 XI11_6/XI0/XI0_20/d__12_ XI11_6/XI0/XI0_20/d_12_ DECAP_INV_G11
XG3751 XI11_6/XI0/XI0_20/d__11_ XI11_6/XI0/XI0_20/d_11_ DECAP_INV_G11
XG3752 XI11_6/XI0/XI0_20/d__10_ XI11_6/XI0/XI0_20/d_10_ DECAP_INV_G11
XG3753 XI11_6/XI0/XI0_20/d__9_ XI11_6/XI0/XI0_20/d_9_ DECAP_INV_G11
XG3754 XI11_6/XI0/XI0_20/d__8_ XI11_6/XI0/XI0_20/d_8_ DECAP_INV_G11
XG3755 XI11_6/XI0/XI0_20/d__7_ XI11_6/XI0/XI0_20/d_7_ DECAP_INV_G11
XG3756 XI11_6/XI0/XI0_20/d__6_ XI11_6/XI0/XI0_20/d_6_ DECAP_INV_G11
XG3757 XI11_6/XI0/XI0_20/d__5_ XI11_6/XI0/XI0_20/d_5_ DECAP_INV_G11
XG3758 XI11_6/XI0/XI0_20/d__4_ XI11_6/XI0/XI0_20/d_4_ DECAP_INV_G11
XG3759 XI11_6/XI0/XI0_20/d__3_ XI11_6/XI0/XI0_20/d_3_ DECAP_INV_G11
XG3760 XI11_6/XI0/XI0_20/d__2_ XI11_6/XI0/XI0_20/d_2_ DECAP_INV_G11
XG3761 XI11_6/XI0/XI0_20/d__1_ XI11_6/XI0/XI0_20/d_1_ DECAP_INV_G11
XG3762 XI11_6/XI0/XI0_20/d__0_ XI11_6/XI0/XI0_20/d_0_ DECAP_INV_G11
XG3763 XI11_6/XI0/XI0_20/d_15_ XI11_6/XI0/XI0_20/d__15_ DECAP_INV_G11
XG3764 XI11_6/XI0/XI0_20/d_14_ XI11_6/XI0/XI0_20/d__14_ DECAP_INV_G11
XG3765 XI11_6/XI0/XI0_20/d_13_ XI11_6/XI0/XI0_20/d__13_ DECAP_INV_G11
XG3766 XI11_6/XI0/XI0_20/d_12_ XI11_6/XI0/XI0_20/d__12_ DECAP_INV_G11
XG3767 XI11_6/XI0/XI0_20/d_11_ XI11_6/XI0/XI0_20/d__11_ DECAP_INV_G11
XG3768 XI11_6/XI0/XI0_20/d_10_ XI11_6/XI0/XI0_20/d__10_ DECAP_INV_G11
XG3769 XI11_6/XI0/XI0_20/d_9_ XI11_6/XI0/XI0_20/d__9_ DECAP_INV_G11
XG3770 XI11_6/XI0/XI0_20/d_8_ XI11_6/XI0/XI0_20/d__8_ DECAP_INV_G11
XG3771 XI11_6/XI0/XI0_20/d_7_ XI11_6/XI0/XI0_20/d__7_ DECAP_INV_G11
XG3772 XI11_6/XI0/XI0_20/d_6_ XI11_6/XI0/XI0_20/d__6_ DECAP_INV_G11
XG3773 XI11_6/XI0/XI0_20/d_5_ XI11_6/XI0/XI0_20/d__5_ DECAP_INV_G11
XG3774 XI11_6/XI0/XI0_20/d_4_ XI11_6/XI0/XI0_20/d__4_ DECAP_INV_G11
XG3775 XI11_6/XI0/XI0_20/d_3_ XI11_6/XI0/XI0_20/d__3_ DECAP_INV_G11
XG3776 XI11_6/XI0/XI0_20/d_2_ XI11_6/XI0/XI0_20/d__2_ DECAP_INV_G11
XG3777 XI11_6/XI0/XI0_20/d_1_ XI11_6/XI0/XI0_20/d__1_ DECAP_INV_G11
XG3778 XI11_6/XI0/XI0_20/d_0_ XI11_6/XI0/XI0_20/d__0_ DECAP_INV_G11
XG3779 XI11_6/XI0/XI0_19/d__15_ XI11_6/XI0/XI0_19/d_15_ DECAP_INV_G11
XG3780 XI11_6/XI0/XI0_19/d__14_ XI11_6/XI0/XI0_19/d_14_ DECAP_INV_G11
XG3781 XI11_6/XI0/XI0_19/d__13_ XI11_6/XI0/XI0_19/d_13_ DECAP_INV_G11
XG3782 XI11_6/XI0/XI0_19/d__12_ XI11_6/XI0/XI0_19/d_12_ DECAP_INV_G11
XG3783 XI11_6/XI0/XI0_19/d__11_ XI11_6/XI0/XI0_19/d_11_ DECAP_INV_G11
XG3784 XI11_6/XI0/XI0_19/d__10_ XI11_6/XI0/XI0_19/d_10_ DECAP_INV_G11
XG3785 XI11_6/XI0/XI0_19/d__9_ XI11_6/XI0/XI0_19/d_9_ DECAP_INV_G11
XG3786 XI11_6/XI0/XI0_19/d__8_ XI11_6/XI0/XI0_19/d_8_ DECAP_INV_G11
XG3787 XI11_6/XI0/XI0_19/d__7_ XI11_6/XI0/XI0_19/d_7_ DECAP_INV_G11
XG3788 XI11_6/XI0/XI0_19/d__6_ XI11_6/XI0/XI0_19/d_6_ DECAP_INV_G11
XG3789 XI11_6/XI0/XI0_19/d__5_ XI11_6/XI0/XI0_19/d_5_ DECAP_INV_G11
XG3790 XI11_6/XI0/XI0_19/d__4_ XI11_6/XI0/XI0_19/d_4_ DECAP_INV_G11
XG3791 XI11_6/XI0/XI0_19/d__3_ XI11_6/XI0/XI0_19/d_3_ DECAP_INV_G11
XG3792 XI11_6/XI0/XI0_19/d__2_ XI11_6/XI0/XI0_19/d_2_ DECAP_INV_G11
XG3793 XI11_6/XI0/XI0_19/d__1_ XI11_6/XI0/XI0_19/d_1_ DECAP_INV_G11
XG3794 XI11_6/XI0/XI0_19/d__0_ XI11_6/XI0/XI0_19/d_0_ DECAP_INV_G11
XG3795 XI11_6/XI0/XI0_19/d_15_ XI11_6/XI0/XI0_19/d__15_ DECAP_INV_G11
XG3796 XI11_6/XI0/XI0_19/d_14_ XI11_6/XI0/XI0_19/d__14_ DECAP_INV_G11
XG3797 XI11_6/XI0/XI0_19/d_13_ XI11_6/XI0/XI0_19/d__13_ DECAP_INV_G11
XG3798 XI11_6/XI0/XI0_19/d_12_ XI11_6/XI0/XI0_19/d__12_ DECAP_INV_G11
XG3799 XI11_6/XI0/XI0_19/d_11_ XI11_6/XI0/XI0_19/d__11_ DECAP_INV_G11
XG3800 XI11_6/XI0/XI0_19/d_10_ XI11_6/XI0/XI0_19/d__10_ DECAP_INV_G11
XG3801 XI11_6/XI0/XI0_19/d_9_ XI11_6/XI0/XI0_19/d__9_ DECAP_INV_G11
XG3802 XI11_6/XI0/XI0_19/d_8_ XI11_6/XI0/XI0_19/d__8_ DECAP_INV_G11
XG3803 XI11_6/XI0/XI0_19/d_7_ XI11_6/XI0/XI0_19/d__7_ DECAP_INV_G11
XG3804 XI11_6/XI0/XI0_19/d_6_ XI11_6/XI0/XI0_19/d__6_ DECAP_INV_G11
XG3805 XI11_6/XI0/XI0_19/d_5_ XI11_6/XI0/XI0_19/d__5_ DECAP_INV_G11
XG3806 XI11_6/XI0/XI0_19/d_4_ XI11_6/XI0/XI0_19/d__4_ DECAP_INV_G11
XG3807 XI11_6/XI0/XI0_19/d_3_ XI11_6/XI0/XI0_19/d__3_ DECAP_INV_G11
XG3808 XI11_6/XI0/XI0_19/d_2_ XI11_6/XI0/XI0_19/d__2_ DECAP_INV_G11
XG3809 XI11_6/XI0/XI0_19/d_1_ XI11_6/XI0/XI0_19/d__1_ DECAP_INV_G11
XG3810 XI11_6/XI0/XI0_19/d_0_ XI11_6/XI0/XI0_19/d__0_ DECAP_INV_G11
XG3811 XI11_6/XI0/XI0_18/d__15_ XI11_6/XI0/XI0_18/d_15_ DECAP_INV_G11
XG3812 XI11_6/XI0/XI0_18/d__14_ XI11_6/XI0/XI0_18/d_14_ DECAP_INV_G11
XG3813 XI11_6/XI0/XI0_18/d__13_ XI11_6/XI0/XI0_18/d_13_ DECAP_INV_G11
XG3814 XI11_6/XI0/XI0_18/d__12_ XI11_6/XI0/XI0_18/d_12_ DECAP_INV_G11
XG3815 XI11_6/XI0/XI0_18/d__11_ XI11_6/XI0/XI0_18/d_11_ DECAP_INV_G11
XG3816 XI11_6/XI0/XI0_18/d__10_ XI11_6/XI0/XI0_18/d_10_ DECAP_INV_G11
XG3817 XI11_6/XI0/XI0_18/d__9_ XI11_6/XI0/XI0_18/d_9_ DECAP_INV_G11
XG3818 XI11_6/XI0/XI0_18/d__8_ XI11_6/XI0/XI0_18/d_8_ DECAP_INV_G11
XG3819 XI11_6/XI0/XI0_18/d__7_ XI11_6/XI0/XI0_18/d_7_ DECAP_INV_G11
XG3820 XI11_6/XI0/XI0_18/d__6_ XI11_6/XI0/XI0_18/d_6_ DECAP_INV_G11
XG3821 XI11_6/XI0/XI0_18/d__5_ XI11_6/XI0/XI0_18/d_5_ DECAP_INV_G11
XG3822 XI11_6/XI0/XI0_18/d__4_ XI11_6/XI0/XI0_18/d_4_ DECAP_INV_G11
XG3823 XI11_6/XI0/XI0_18/d__3_ XI11_6/XI0/XI0_18/d_3_ DECAP_INV_G11
XG3824 XI11_6/XI0/XI0_18/d__2_ XI11_6/XI0/XI0_18/d_2_ DECAP_INV_G11
XG3825 XI11_6/XI0/XI0_18/d__1_ XI11_6/XI0/XI0_18/d_1_ DECAP_INV_G11
XG3826 XI11_6/XI0/XI0_18/d__0_ XI11_6/XI0/XI0_18/d_0_ DECAP_INV_G11
XG3827 XI11_6/XI0/XI0_18/d_15_ XI11_6/XI0/XI0_18/d__15_ DECAP_INV_G11
XG3828 XI11_6/XI0/XI0_18/d_14_ XI11_6/XI0/XI0_18/d__14_ DECAP_INV_G11
XG3829 XI11_6/XI0/XI0_18/d_13_ XI11_6/XI0/XI0_18/d__13_ DECAP_INV_G11
XG3830 XI11_6/XI0/XI0_18/d_12_ XI11_6/XI0/XI0_18/d__12_ DECAP_INV_G11
XG3831 XI11_6/XI0/XI0_18/d_11_ XI11_6/XI0/XI0_18/d__11_ DECAP_INV_G11
XG3832 XI11_6/XI0/XI0_18/d_10_ XI11_6/XI0/XI0_18/d__10_ DECAP_INV_G11
XG3833 XI11_6/XI0/XI0_18/d_9_ XI11_6/XI0/XI0_18/d__9_ DECAP_INV_G11
XG3834 XI11_6/XI0/XI0_18/d_8_ XI11_6/XI0/XI0_18/d__8_ DECAP_INV_G11
XG3835 XI11_6/XI0/XI0_18/d_7_ XI11_6/XI0/XI0_18/d__7_ DECAP_INV_G11
XG3836 XI11_6/XI0/XI0_18/d_6_ XI11_6/XI0/XI0_18/d__6_ DECAP_INV_G11
XG3837 XI11_6/XI0/XI0_18/d_5_ XI11_6/XI0/XI0_18/d__5_ DECAP_INV_G11
XG3838 XI11_6/XI0/XI0_18/d_4_ XI11_6/XI0/XI0_18/d__4_ DECAP_INV_G11
XG3839 XI11_6/XI0/XI0_18/d_3_ XI11_6/XI0/XI0_18/d__3_ DECAP_INV_G11
XG3840 XI11_6/XI0/XI0_18/d_2_ XI11_6/XI0/XI0_18/d__2_ DECAP_INV_G11
XG3841 XI11_6/XI0/XI0_18/d_1_ XI11_6/XI0/XI0_18/d__1_ DECAP_INV_G11
XG3842 XI11_6/XI0/XI0_18/d_0_ XI11_6/XI0/XI0_18/d__0_ DECAP_INV_G11
XG3843 XI11_6/XI0/XI0_17/d__15_ XI11_6/XI0/XI0_17/d_15_ DECAP_INV_G11
XG3844 XI11_6/XI0/XI0_17/d__14_ XI11_6/XI0/XI0_17/d_14_ DECAP_INV_G11
XG3845 XI11_6/XI0/XI0_17/d__13_ XI11_6/XI0/XI0_17/d_13_ DECAP_INV_G11
XG3846 XI11_6/XI0/XI0_17/d__12_ XI11_6/XI0/XI0_17/d_12_ DECAP_INV_G11
XG3847 XI11_6/XI0/XI0_17/d__11_ XI11_6/XI0/XI0_17/d_11_ DECAP_INV_G11
XG3848 XI11_6/XI0/XI0_17/d__10_ XI11_6/XI0/XI0_17/d_10_ DECAP_INV_G11
XG3849 XI11_6/XI0/XI0_17/d__9_ XI11_6/XI0/XI0_17/d_9_ DECAP_INV_G11
XG3850 XI11_6/XI0/XI0_17/d__8_ XI11_6/XI0/XI0_17/d_8_ DECAP_INV_G11
XG3851 XI11_6/XI0/XI0_17/d__7_ XI11_6/XI0/XI0_17/d_7_ DECAP_INV_G11
XG3852 XI11_6/XI0/XI0_17/d__6_ XI11_6/XI0/XI0_17/d_6_ DECAP_INV_G11
XG3853 XI11_6/XI0/XI0_17/d__5_ XI11_6/XI0/XI0_17/d_5_ DECAP_INV_G11
XG3854 XI11_6/XI0/XI0_17/d__4_ XI11_6/XI0/XI0_17/d_4_ DECAP_INV_G11
XG3855 XI11_6/XI0/XI0_17/d__3_ XI11_6/XI0/XI0_17/d_3_ DECAP_INV_G11
XG3856 XI11_6/XI0/XI0_17/d__2_ XI11_6/XI0/XI0_17/d_2_ DECAP_INV_G11
XG3857 XI11_6/XI0/XI0_17/d__1_ XI11_6/XI0/XI0_17/d_1_ DECAP_INV_G11
XG3858 XI11_6/XI0/XI0_17/d__0_ XI11_6/XI0/XI0_17/d_0_ DECAP_INV_G11
XG3859 XI11_6/XI0/XI0_17/d_15_ XI11_6/XI0/XI0_17/d__15_ DECAP_INV_G11
XG3860 XI11_6/XI0/XI0_17/d_14_ XI11_6/XI0/XI0_17/d__14_ DECAP_INV_G11
XG3861 XI11_6/XI0/XI0_17/d_13_ XI11_6/XI0/XI0_17/d__13_ DECAP_INV_G11
XG3862 XI11_6/XI0/XI0_17/d_12_ XI11_6/XI0/XI0_17/d__12_ DECAP_INV_G11
XG3863 XI11_6/XI0/XI0_17/d_11_ XI11_6/XI0/XI0_17/d__11_ DECAP_INV_G11
XG3864 XI11_6/XI0/XI0_17/d_10_ XI11_6/XI0/XI0_17/d__10_ DECAP_INV_G11
XG3865 XI11_6/XI0/XI0_17/d_9_ XI11_6/XI0/XI0_17/d__9_ DECAP_INV_G11
XG3866 XI11_6/XI0/XI0_17/d_8_ XI11_6/XI0/XI0_17/d__8_ DECAP_INV_G11
XG3867 XI11_6/XI0/XI0_17/d_7_ XI11_6/XI0/XI0_17/d__7_ DECAP_INV_G11
XG3868 XI11_6/XI0/XI0_17/d_6_ XI11_6/XI0/XI0_17/d__6_ DECAP_INV_G11
XG3869 XI11_6/XI0/XI0_17/d_5_ XI11_6/XI0/XI0_17/d__5_ DECAP_INV_G11
XG3870 XI11_6/XI0/XI0_17/d_4_ XI11_6/XI0/XI0_17/d__4_ DECAP_INV_G11
XG3871 XI11_6/XI0/XI0_17/d_3_ XI11_6/XI0/XI0_17/d__3_ DECAP_INV_G11
XG3872 XI11_6/XI0/XI0_17/d_2_ XI11_6/XI0/XI0_17/d__2_ DECAP_INV_G11
XG3873 XI11_6/XI0/XI0_17/d_1_ XI11_6/XI0/XI0_17/d__1_ DECAP_INV_G11
XG3874 XI11_6/XI0/XI0_17/d_0_ XI11_6/XI0/XI0_17/d__0_ DECAP_INV_G11
XG3875 XI11_6/XI0/XI0_16/d__15_ XI11_6/XI0/XI0_16/d_15_ DECAP_INV_G11
XG3876 XI11_6/XI0/XI0_16/d__14_ XI11_6/XI0/XI0_16/d_14_ DECAP_INV_G11
XG3877 XI11_6/XI0/XI0_16/d__13_ XI11_6/XI0/XI0_16/d_13_ DECAP_INV_G11
XG3878 XI11_6/XI0/XI0_16/d__12_ XI11_6/XI0/XI0_16/d_12_ DECAP_INV_G11
XG3879 XI11_6/XI0/XI0_16/d__11_ XI11_6/XI0/XI0_16/d_11_ DECAP_INV_G11
XG3880 XI11_6/XI0/XI0_16/d__10_ XI11_6/XI0/XI0_16/d_10_ DECAP_INV_G11
XG3881 XI11_6/XI0/XI0_16/d__9_ XI11_6/XI0/XI0_16/d_9_ DECAP_INV_G11
XG3882 XI11_6/XI0/XI0_16/d__8_ XI11_6/XI0/XI0_16/d_8_ DECAP_INV_G11
XG3883 XI11_6/XI0/XI0_16/d__7_ XI11_6/XI0/XI0_16/d_7_ DECAP_INV_G11
XG3884 XI11_6/XI0/XI0_16/d__6_ XI11_6/XI0/XI0_16/d_6_ DECAP_INV_G11
XG3885 XI11_6/XI0/XI0_16/d__5_ XI11_6/XI0/XI0_16/d_5_ DECAP_INV_G11
XG3886 XI11_6/XI0/XI0_16/d__4_ XI11_6/XI0/XI0_16/d_4_ DECAP_INV_G11
XG3887 XI11_6/XI0/XI0_16/d__3_ XI11_6/XI0/XI0_16/d_3_ DECAP_INV_G11
XG3888 XI11_6/XI0/XI0_16/d__2_ XI11_6/XI0/XI0_16/d_2_ DECAP_INV_G11
XG3889 XI11_6/XI0/XI0_16/d__1_ XI11_6/XI0/XI0_16/d_1_ DECAP_INV_G11
XG3890 XI11_6/XI0/XI0_16/d__0_ XI11_6/XI0/XI0_16/d_0_ DECAP_INV_G11
XG3891 XI11_6/XI0/XI0_16/d_15_ XI11_6/XI0/XI0_16/d__15_ DECAP_INV_G11
XG3892 XI11_6/XI0/XI0_16/d_14_ XI11_6/XI0/XI0_16/d__14_ DECAP_INV_G11
XG3893 XI11_6/XI0/XI0_16/d_13_ XI11_6/XI0/XI0_16/d__13_ DECAP_INV_G11
XG3894 XI11_6/XI0/XI0_16/d_12_ XI11_6/XI0/XI0_16/d__12_ DECAP_INV_G11
XG3895 XI11_6/XI0/XI0_16/d_11_ XI11_6/XI0/XI0_16/d__11_ DECAP_INV_G11
XG3896 XI11_6/XI0/XI0_16/d_10_ XI11_6/XI0/XI0_16/d__10_ DECAP_INV_G11
XG3897 XI11_6/XI0/XI0_16/d_9_ XI11_6/XI0/XI0_16/d__9_ DECAP_INV_G11
XG3898 XI11_6/XI0/XI0_16/d_8_ XI11_6/XI0/XI0_16/d__8_ DECAP_INV_G11
XG3899 XI11_6/XI0/XI0_16/d_7_ XI11_6/XI0/XI0_16/d__7_ DECAP_INV_G11
XG3900 XI11_6/XI0/XI0_16/d_6_ XI11_6/XI0/XI0_16/d__6_ DECAP_INV_G11
XG3901 XI11_6/XI0/XI0_16/d_5_ XI11_6/XI0/XI0_16/d__5_ DECAP_INV_G11
XG3902 XI11_6/XI0/XI0_16/d_4_ XI11_6/XI0/XI0_16/d__4_ DECAP_INV_G11
XG3903 XI11_6/XI0/XI0_16/d_3_ XI11_6/XI0/XI0_16/d__3_ DECAP_INV_G11
XG3904 XI11_6/XI0/XI0_16/d_2_ XI11_6/XI0/XI0_16/d__2_ DECAP_INV_G11
XG3905 XI11_6/XI0/XI0_16/d_1_ XI11_6/XI0/XI0_16/d__1_ DECAP_INV_G11
XG3906 XI11_6/XI0/XI0_16/d_0_ XI11_6/XI0/XI0_16/d__0_ DECAP_INV_G11
XG3907 XI11_6/XI0/XI0_15/d__15_ XI11_6/XI0/XI0_15/d_15_ DECAP_INV_G11
XG3908 XI11_6/XI0/XI0_15/d__14_ XI11_6/XI0/XI0_15/d_14_ DECAP_INV_G11
XG3909 XI11_6/XI0/XI0_15/d__13_ XI11_6/XI0/XI0_15/d_13_ DECAP_INV_G11
XG3910 XI11_6/XI0/XI0_15/d__12_ XI11_6/XI0/XI0_15/d_12_ DECAP_INV_G11
XG3911 XI11_6/XI0/XI0_15/d__11_ XI11_6/XI0/XI0_15/d_11_ DECAP_INV_G11
XG3912 XI11_6/XI0/XI0_15/d__10_ XI11_6/XI0/XI0_15/d_10_ DECAP_INV_G11
XG3913 XI11_6/XI0/XI0_15/d__9_ XI11_6/XI0/XI0_15/d_9_ DECAP_INV_G11
XG3914 XI11_6/XI0/XI0_15/d__8_ XI11_6/XI0/XI0_15/d_8_ DECAP_INV_G11
XG3915 XI11_6/XI0/XI0_15/d__7_ XI11_6/XI0/XI0_15/d_7_ DECAP_INV_G11
XG3916 XI11_6/XI0/XI0_15/d__6_ XI11_6/XI0/XI0_15/d_6_ DECAP_INV_G11
XG3917 XI11_6/XI0/XI0_15/d__5_ XI11_6/XI0/XI0_15/d_5_ DECAP_INV_G11
XG3918 XI11_6/XI0/XI0_15/d__4_ XI11_6/XI0/XI0_15/d_4_ DECAP_INV_G11
XG3919 XI11_6/XI0/XI0_15/d__3_ XI11_6/XI0/XI0_15/d_3_ DECAP_INV_G11
XG3920 XI11_6/XI0/XI0_15/d__2_ XI11_6/XI0/XI0_15/d_2_ DECAP_INV_G11
XG3921 XI11_6/XI0/XI0_15/d__1_ XI11_6/XI0/XI0_15/d_1_ DECAP_INV_G11
XG3922 XI11_6/XI0/XI0_15/d__0_ XI11_6/XI0/XI0_15/d_0_ DECAP_INV_G11
XG3923 XI11_6/XI0/XI0_15/d_15_ XI11_6/XI0/XI0_15/d__15_ DECAP_INV_G11
XG3924 XI11_6/XI0/XI0_15/d_14_ XI11_6/XI0/XI0_15/d__14_ DECAP_INV_G11
XG3925 XI11_6/XI0/XI0_15/d_13_ XI11_6/XI0/XI0_15/d__13_ DECAP_INV_G11
XG3926 XI11_6/XI0/XI0_15/d_12_ XI11_6/XI0/XI0_15/d__12_ DECAP_INV_G11
XG3927 XI11_6/XI0/XI0_15/d_11_ XI11_6/XI0/XI0_15/d__11_ DECAP_INV_G11
XG3928 XI11_6/XI0/XI0_15/d_10_ XI11_6/XI0/XI0_15/d__10_ DECAP_INV_G11
XG3929 XI11_6/XI0/XI0_15/d_9_ XI11_6/XI0/XI0_15/d__9_ DECAP_INV_G11
XG3930 XI11_6/XI0/XI0_15/d_8_ XI11_6/XI0/XI0_15/d__8_ DECAP_INV_G11
XG3931 XI11_6/XI0/XI0_15/d_7_ XI11_6/XI0/XI0_15/d__7_ DECAP_INV_G11
XG3932 XI11_6/XI0/XI0_15/d_6_ XI11_6/XI0/XI0_15/d__6_ DECAP_INV_G11
XG3933 XI11_6/XI0/XI0_15/d_5_ XI11_6/XI0/XI0_15/d__5_ DECAP_INV_G11
XG3934 XI11_6/XI0/XI0_15/d_4_ XI11_6/XI0/XI0_15/d__4_ DECAP_INV_G11
XG3935 XI11_6/XI0/XI0_15/d_3_ XI11_6/XI0/XI0_15/d__3_ DECAP_INV_G11
XG3936 XI11_6/XI0/XI0_15/d_2_ XI11_6/XI0/XI0_15/d__2_ DECAP_INV_G11
XG3937 XI11_6/XI0/XI0_15/d_1_ XI11_6/XI0/XI0_15/d__1_ DECAP_INV_G11
XG3938 XI11_6/XI0/XI0_15/d_0_ XI11_6/XI0/XI0_15/d__0_ DECAP_INV_G11
XG3939 XI11_6/XI0/XI0_14/d__15_ XI11_6/XI0/XI0_14/d_15_ DECAP_INV_G11
XG3940 XI11_6/XI0/XI0_14/d__14_ XI11_6/XI0/XI0_14/d_14_ DECAP_INV_G11
XG3941 XI11_6/XI0/XI0_14/d__13_ XI11_6/XI0/XI0_14/d_13_ DECAP_INV_G11
XG3942 XI11_6/XI0/XI0_14/d__12_ XI11_6/XI0/XI0_14/d_12_ DECAP_INV_G11
XG3943 XI11_6/XI0/XI0_14/d__11_ XI11_6/XI0/XI0_14/d_11_ DECAP_INV_G11
XG3944 XI11_6/XI0/XI0_14/d__10_ XI11_6/XI0/XI0_14/d_10_ DECAP_INV_G11
XG3945 XI11_6/XI0/XI0_14/d__9_ XI11_6/XI0/XI0_14/d_9_ DECAP_INV_G11
XG3946 XI11_6/XI0/XI0_14/d__8_ XI11_6/XI0/XI0_14/d_8_ DECAP_INV_G11
XG3947 XI11_6/XI0/XI0_14/d__7_ XI11_6/XI0/XI0_14/d_7_ DECAP_INV_G11
XG3948 XI11_6/XI0/XI0_14/d__6_ XI11_6/XI0/XI0_14/d_6_ DECAP_INV_G11
XG3949 XI11_6/XI0/XI0_14/d__5_ XI11_6/XI0/XI0_14/d_5_ DECAP_INV_G11
XG3950 XI11_6/XI0/XI0_14/d__4_ XI11_6/XI0/XI0_14/d_4_ DECAP_INV_G11
XG3951 XI11_6/XI0/XI0_14/d__3_ XI11_6/XI0/XI0_14/d_3_ DECAP_INV_G11
XG3952 XI11_6/XI0/XI0_14/d__2_ XI11_6/XI0/XI0_14/d_2_ DECAP_INV_G11
XG3953 XI11_6/XI0/XI0_14/d__1_ XI11_6/XI0/XI0_14/d_1_ DECAP_INV_G11
XG3954 XI11_6/XI0/XI0_14/d__0_ XI11_6/XI0/XI0_14/d_0_ DECAP_INV_G11
XG3955 XI11_6/XI0/XI0_14/d_15_ XI11_6/XI0/XI0_14/d__15_ DECAP_INV_G11
XG3956 XI11_6/XI0/XI0_14/d_14_ XI11_6/XI0/XI0_14/d__14_ DECAP_INV_G11
XG3957 XI11_6/XI0/XI0_14/d_13_ XI11_6/XI0/XI0_14/d__13_ DECAP_INV_G11
XG3958 XI11_6/XI0/XI0_14/d_12_ XI11_6/XI0/XI0_14/d__12_ DECAP_INV_G11
XG3959 XI11_6/XI0/XI0_14/d_11_ XI11_6/XI0/XI0_14/d__11_ DECAP_INV_G11
XG3960 XI11_6/XI0/XI0_14/d_10_ XI11_6/XI0/XI0_14/d__10_ DECAP_INV_G11
XG3961 XI11_6/XI0/XI0_14/d_9_ XI11_6/XI0/XI0_14/d__9_ DECAP_INV_G11
XG3962 XI11_6/XI0/XI0_14/d_8_ XI11_6/XI0/XI0_14/d__8_ DECAP_INV_G11
XG3963 XI11_6/XI0/XI0_14/d_7_ XI11_6/XI0/XI0_14/d__7_ DECAP_INV_G11
XG3964 XI11_6/XI0/XI0_14/d_6_ XI11_6/XI0/XI0_14/d__6_ DECAP_INV_G11
XG3965 XI11_6/XI0/XI0_14/d_5_ XI11_6/XI0/XI0_14/d__5_ DECAP_INV_G11
XG3966 XI11_6/XI0/XI0_14/d_4_ XI11_6/XI0/XI0_14/d__4_ DECAP_INV_G11
XG3967 XI11_6/XI0/XI0_14/d_3_ XI11_6/XI0/XI0_14/d__3_ DECAP_INV_G11
XG3968 XI11_6/XI0/XI0_14/d_2_ XI11_6/XI0/XI0_14/d__2_ DECAP_INV_G11
XG3969 XI11_6/XI0/XI0_14/d_1_ XI11_6/XI0/XI0_14/d__1_ DECAP_INV_G11
XG3970 XI11_6/XI0/XI0_14/d_0_ XI11_6/XI0/XI0_14/d__0_ DECAP_INV_G11
XG3971 XI11_6/XI0/XI0_13/d__15_ XI11_6/XI0/XI0_13/d_15_ DECAP_INV_G11
XG3972 XI11_6/XI0/XI0_13/d__14_ XI11_6/XI0/XI0_13/d_14_ DECAP_INV_G11
XG3973 XI11_6/XI0/XI0_13/d__13_ XI11_6/XI0/XI0_13/d_13_ DECAP_INV_G11
XG3974 XI11_6/XI0/XI0_13/d__12_ XI11_6/XI0/XI0_13/d_12_ DECAP_INV_G11
XG3975 XI11_6/XI0/XI0_13/d__11_ XI11_6/XI0/XI0_13/d_11_ DECAP_INV_G11
XG3976 XI11_6/XI0/XI0_13/d__10_ XI11_6/XI0/XI0_13/d_10_ DECAP_INV_G11
XG3977 XI11_6/XI0/XI0_13/d__9_ XI11_6/XI0/XI0_13/d_9_ DECAP_INV_G11
XG3978 XI11_6/XI0/XI0_13/d__8_ XI11_6/XI0/XI0_13/d_8_ DECAP_INV_G11
XG3979 XI11_6/XI0/XI0_13/d__7_ XI11_6/XI0/XI0_13/d_7_ DECAP_INV_G11
XG3980 XI11_6/XI0/XI0_13/d__6_ XI11_6/XI0/XI0_13/d_6_ DECAP_INV_G11
XG3981 XI11_6/XI0/XI0_13/d__5_ XI11_6/XI0/XI0_13/d_5_ DECAP_INV_G11
XG3982 XI11_6/XI0/XI0_13/d__4_ XI11_6/XI0/XI0_13/d_4_ DECAP_INV_G11
XG3983 XI11_6/XI0/XI0_13/d__3_ XI11_6/XI0/XI0_13/d_3_ DECAP_INV_G11
XG3984 XI11_6/XI0/XI0_13/d__2_ XI11_6/XI0/XI0_13/d_2_ DECAP_INV_G11
XG3985 XI11_6/XI0/XI0_13/d__1_ XI11_6/XI0/XI0_13/d_1_ DECAP_INV_G11
XG3986 XI11_6/XI0/XI0_13/d__0_ XI11_6/XI0/XI0_13/d_0_ DECAP_INV_G11
XG3987 XI11_6/XI0/XI0_13/d_15_ XI11_6/XI0/XI0_13/d__15_ DECAP_INV_G11
XG3988 XI11_6/XI0/XI0_13/d_14_ XI11_6/XI0/XI0_13/d__14_ DECAP_INV_G11
XG3989 XI11_6/XI0/XI0_13/d_13_ XI11_6/XI0/XI0_13/d__13_ DECAP_INV_G11
XG3990 XI11_6/XI0/XI0_13/d_12_ XI11_6/XI0/XI0_13/d__12_ DECAP_INV_G11
XG3991 XI11_6/XI0/XI0_13/d_11_ XI11_6/XI0/XI0_13/d__11_ DECAP_INV_G11
XG3992 XI11_6/XI0/XI0_13/d_10_ XI11_6/XI0/XI0_13/d__10_ DECAP_INV_G11
XG3993 XI11_6/XI0/XI0_13/d_9_ XI11_6/XI0/XI0_13/d__9_ DECAP_INV_G11
XG3994 XI11_6/XI0/XI0_13/d_8_ XI11_6/XI0/XI0_13/d__8_ DECAP_INV_G11
XG3995 XI11_6/XI0/XI0_13/d_7_ XI11_6/XI0/XI0_13/d__7_ DECAP_INV_G11
XG3996 XI11_6/XI0/XI0_13/d_6_ XI11_6/XI0/XI0_13/d__6_ DECAP_INV_G11
XG3997 XI11_6/XI0/XI0_13/d_5_ XI11_6/XI0/XI0_13/d__5_ DECAP_INV_G11
XG3998 XI11_6/XI0/XI0_13/d_4_ XI11_6/XI0/XI0_13/d__4_ DECAP_INV_G11
XG3999 XI11_6/XI0/XI0_13/d_3_ XI11_6/XI0/XI0_13/d__3_ DECAP_INV_G11
XG4000 XI11_6/XI0/XI0_13/d_2_ XI11_6/XI0/XI0_13/d__2_ DECAP_INV_G11
XG4001 XI11_6/XI0/XI0_13/d_1_ XI11_6/XI0/XI0_13/d__1_ DECAP_INV_G11
XG4002 XI11_6/XI0/XI0_13/d_0_ XI11_6/XI0/XI0_13/d__0_ DECAP_INV_G11
XG4003 XI11_6/XI0/XI0_12/d__15_ XI11_6/XI0/XI0_12/d_15_ DECAP_INV_G11
XG4004 XI11_6/XI0/XI0_12/d__14_ XI11_6/XI0/XI0_12/d_14_ DECAP_INV_G11
XG4005 XI11_6/XI0/XI0_12/d__13_ XI11_6/XI0/XI0_12/d_13_ DECAP_INV_G11
XG4006 XI11_6/XI0/XI0_12/d__12_ XI11_6/XI0/XI0_12/d_12_ DECAP_INV_G11
XG4007 XI11_6/XI0/XI0_12/d__11_ XI11_6/XI0/XI0_12/d_11_ DECAP_INV_G11
XG4008 XI11_6/XI0/XI0_12/d__10_ XI11_6/XI0/XI0_12/d_10_ DECAP_INV_G11
XG4009 XI11_6/XI0/XI0_12/d__9_ XI11_6/XI0/XI0_12/d_9_ DECAP_INV_G11
XG4010 XI11_6/XI0/XI0_12/d__8_ XI11_6/XI0/XI0_12/d_8_ DECAP_INV_G11
XG4011 XI11_6/XI0/XI0_12/d__7_ XI11_6/XI0/XI0_12/d_7_ DECAP_INV_G11
XG4012 XI11_6/XI0/XI0_12/d__6_ XI11_6/XI0/XI0_12/d_6_ DECAP_INV_G11
XG4013 XI11_6/XI0/XI0_12/d__5_ XI11_6/XI0/XI0_12/d_5_ DECAP_INV_G11
XG4014 XI11_6/XI0/XI0_12/d__4_ XI11_6/XI0/XI0_12/d_4_ DECAP_INV_G11
XG4015 XI11_6/XI0/XI0_12/d__3_ XI11_6/XI0/XI0_12/d_3_ DECAP_INV_G11
XG4016 XI11_6/XI0/XI0_12/d__2_ XI11_6/XI0/XI0_12/d_2_ DECAP_INV_G11
XG4017 XI11_6/XI0/XI0_12/d__1_ XI11_6/XI0/XI0_12/d_1_ DECAP_INV_G11
XG4018 XI11_6/XI0/XI0_12/d__0_ XI11_6/XI0/XI0_12/d_0_ DECAP_INV_G11
XG4019 XI11_6/XI0/XI0_12/d_15_ XI11_6/XI0/XI0_12/d__15_ DECAP_INV_G11
XG4020 XI11_6/XI0/XI0_12/d_14_ XI11_6/XI0/XI0_12/d__14_ DECAP_INV_G11
XG4021 XI11_6/XI0/XI0_12/d_13_ XI11_6/XI0/XI0_12/d__13_ DECAP_INV_G11
XG4022 XI11_6/XI0/XI0_12/d_12_ XI11_6/XI0/XI0_12/d__12_ DECAP_INV_G11
XG4023 XI11_6/XI0/XI0_12/d_11_ XI11_6/XI0/XI0_12/d__11_ DECAP_INV_G11
XG4024 XI11_6/XI0/XI0_12/d_10_ XI11_6/XI0/XI0_12/d__10_ DECAP_INV_G11
XG4025 XI11_6/XI0/XI0_12/d_9_ XI11_6/XI0/XI0_12/d__9_ DECAP_INV_G11
XG4026 XI11_6/XI0/XI0_12/d_8_ XI11_6/XI0/XI0_12/d__8_ DECAP_INV_G11
XG4027 XI11_6/XI0/XI0_12/d_7_ XI11_6/XI0/XI0_12/d__7_ DECAP_INV_G11
XG4028 XI11_6/XI0/XI0_12/d_6_ XI11_6/XI0/XI0_12/d__6_ DECAP_INV_G11
XG4029 XI11_6/XI0/XI0_12/d_5_ XI11_6/XI0/XI0_12/d__5_ DECAP_INV_G11
XG4030 XI11_6/XI0/XI0_12/d_4_ XI11_6/XI0/XI0_12/d__4_ DECAP_INV_G11
XG4031 XI11_6/XI0/XI0_12/d_3_ XI11_6/XI0/XI0_12/d__3_ DECAP_INV_G11
XG4032 XI11_6/XI0/XI0_12/d_2_ XI11_6/XI0/XI0_12/d__2_ DECAP_INV_G11
XG4033 XI11_6/XI0/XI0_12/d_1_ XI11_6/XI0/XI0_12/d__1_ DECAP_INV_G11
XG4034 XI11_6/XI0/XI0_12/d_0_ XI11_6/XI0/XI0_12/d__0_ DECAP_INV_G11
XG4035 XI11_6/XI0/XI0_11/d__15_ XI11_6/XI0/XI0_11/d_15_ DECAP_INV_G11
XG4036 XI11_6/XI0/XI0_11/d__14_ XI11_6/XI0/XI0_11/d_14_ DECAP_INV_G11
XG4037 XI11_6/XI0/XI0_11/d__13_ XI11_6/XI0/XI0_11/d_13_ DECAP_INV_G11
XG4038 XI11_6/XI0/XI0_11/d__12_ XI11_6/XI0/XI0_11/d_12_ DECAP_INV_G11
XG4039 XI11_6/XI0/XI0_11/d__11_ XI11_6/XI0/XI0_11/d_11_ DECAP_INV_G11
XG4040 XI11_6/XI0/XI0_11/d__10_ XI11_6/XI0/XI0_11/d_10_ DECAP_INV_G11
XG4041 XI11_6/XI0/XI0_11/d__9_ XI11_6/XI0/XI0_11/d_9_ DECAP_INV_G11
XG4042 XI11_6/XI0/XI0_11/d__8_ XI11_6/XI0/XI0_11/d_8_ DECAP_INV_G11
XG4043 XI11_6/XI0/XI0_11/d__7_ XI11_6/XI0/XI0_11/d_7_ DECAP_INV_G11
XG4044 XI11_6/XI0/XI0_11/d__6_ XI11_6/XI0/XI0_11/d_6_ DECAP_INV_G11
XG4045 XI11_6/XI0/XI0_11/d__5_ XI11_6/XI0/XI0_11/d_5_ DECAP_INV_G11
XG4046 XI11_6/XI0/XI0_11/d__4_ XI11_6/XI0/XI0_11/d_4_ DECAP_INV_G11
XG4047 XI11_6/XI0/XI0_11/d__3_ XI11_6/XI0/XI0_11/d_3_ DECAP_INV_G11
XG4048 XI11_6/XI0/XI0_11/d__2_ XI11_6/XI0/XI0_11/d_2_ DECAP_INV_G11
XG4049 XI11_6/XI0/XI0_11/d__1_ XI11_6/XI0/XI0_11/d_1_ DECAP_INV_G11
XG4050 XI11_6/XI0/XI0_11/d__0_ XI11_6/XI0/XI0_11/d_0_ DECAP_INV_G11
XG4051 XI11_6/XI0/XI0_11/d_15_ XI11_6/XI0/XI0_11/d__15_ DECAP_INV_G11
XG4052 XI11_6/XI0/XI0_11/d_14_ XI11_6/XI0/XI0_11/d__14_ DECAP_INV_G11
XG4053 XI11_6/XI0/XI0_11/d_13_ XI11_6/XI0/XI0_11/d__13_ DECAP_INV_G11
XG4054 XI11_6/XI0/XI0_11/d_12_ XI11_6/XI0/XI0_11/d__12_ DECAP_INV_G11
XG4055 XI11_6/XI0/XI0_11/d_11_ XI11_6/XI0/XI0_11/d__11_ DECAP_INV_G11
XG4056 XI11_6/XI0/XI0_11/d_10_ XI11_6/XI0/XI0_11/d__10_ DECAP_INV_G11
XG4057 XI11_6/XI0/XI0_11/d_9_ XI11_6/XI0/XI0_11/d__9_ DECAP_INV_G11
XG4058 XI11_6/XI0/XI0_11/d_8_ XI11_6/XI0/XI0_11/d__8_ DECAP_INV_G11
XG4059 XI11_6/XI0/XI0_11/d_7_ XI11_6/XI0/XI0_11/d__7_ DECAP_INV_G11
XG4060 XI11_6/XI0/XI0_11/d_6_ XI11_6/XI0/XI0_11/d__6_ DECAP_INV_G11
XG4061 XI11_6/XI0/XI0_11/d_5_ XI11_6/XI0/XI0_11/d__5_ DECAP_INV_G11
XG4062 XI11_6/XI0/XI0_11/d_4_ XI11_6/XI0/XI0_11/d__4_ DECAP_INV_G11
XG4063 XI11_6/XI0/XI0_11/d_3_ XI11_6/XI0/XI0_11/d__3_ DECAP_INV_G11
XG4064 XI11_6/XI0/XI0_11/d_2_ XI11_6/XI0/XI0_11/d__2_ DECAP_INV_G11
XG4065 XI11_6/XI0/XI0_11/d_1_ XI11_6/XI0/XI0_11/d__1_ DECAP_INV_G11
XG4066 XI11_6/XI0/XI0_11/d_0_ XI11_6/XI0/XI0_11/d__0_ DECAP_INV_G11
XG4067 XI11_6/XI0/XI0_10/d__15_ XI11_6/XI0/XI0_10/d_15_ DECAP_INV_G11
XG4068 XI11_6/XI0/XI0_10/d__14_ XI11_6/XI0/XI0_10/d_14_ DECAP_INV_G11
XG4069 XI11_6/XI0/XI0_10/d__13_ XI11_6/XI0/XI0_10/d_13_ DECAP_INV_G11
XG4070 XI11_6/XI0/XI0_10/d__12_ XI11_6/XI0/XI0_10/d_12_ DECAP_INV_G11
XG4071 XI11_6/XI0/XI0_10/d__11_ XI11_6/XI0/XI0_10/d_11_ DECAP_INV_G11
XG4072 XI11_6/XI0/XI0_10/d__10_ XI11_6/XI0/XI0_10/d_10_ DECAP_INV_G11
XG4073 XI11_6/XI0/XI0_10/d__9_ XI11_6/XI0/XI0_10/d_9_ DECAP_INV_G11
XG4074 XI11_6/XI0/XI0_10/d__8_ XI11_6/XI0/XI0_10/d_8_ DECAP_INV_G11
XG4075 XI11_6/XI0/XI0_10/d__7_ XI11_6/XI0/XI0_10/d_7_ DECAP_INV_G11
XG4076 XI11_6/XI0/XI0_10/d__6_ XI11_6/XI0/XI0_10/d_6_ DECAP_INV_G11
XG4077 XI11_6/XI0/XI0_10/d__5_ XI11_6/XI0/XI0_10/d_5_ DECAP_INV_G11
XG4078 XI11_6/XI0/XI0_10/d__4_ XI11_6/XI0/XI0_10/d_4_ DECAP_INV_G11
XG4079 XI11_6/XI0/XI0_10/d__3_ XI11_6/XI0/XI0_10/d_3_ DECAP_INV_G11
XG4080 XI11_6/XI0/XI0_10/d__2_ XI11_6/XI0/XI0_10/d_2_ DECAP_INV_G11
XG4081 XI11_6/XI0/XI0_10/d__1_ XI11_6/XI0/XI0_10/d_1_ DECAP_INV_G11
XG4082 XI11_6/XI0/XI0_10/d__0_ XI11_6/XI0/XI0_10/d_0_ DECAP_INV_G11
XG4083 XI11_6/XI0/XI0_10/d_15_ XI11_6/XI0/XI0_10/d__15_ DECAP_INV_G11
XG4084 XI11_6/XI0/XI0_10/d_14_ XI11_6/XI0/XI0_10/d__14_ DECAP_INV_G11
XG4085 XI11_6/XI0/XI0_10/d_13_ XI11_6/XI0/XI0_10/d__13_ DECAP_INV_G11
XG4086 XI11_6/XI0/XI0_10/d_12_ XI11_6/XI0/XI0_10/d__12_ DECAP_INV_G11
XG4087 XI11_6/XI0/XI0_10/d_11_ XI11_6/XI0/XI0_10/d__11_ DECAP_INV_G11
XG4088 XI11_6/XI0/XI0_10/d_10_ XI11_6/XI0/XI0_10/d__10_ DECAP_INV_G11
XG4089 XI11_6/XI0/XI0_10/d_9_ XI11_6/XI0/XI0_10/d__9_ DECAP_INV_G11
XG4090 XI11_6/XI0/XI0_10/d_8_ XI11_6/XI0/XI0_10/d__8_ DECAP_INV_G11
XG4091 XI11_6/XI0/XI0_10/d_7_ XI11_6/XI0/XI0_10/d__7_ DECAP_INV_G11
XG4092 XI11_6/XI0/XI0_10/d_6_ XI11_6/XI0/XI0_10/d__6_ DECAP_INV_G11
XG4093 XI11_6/XI0/XI0_10/d_5_ XI11_6/XI0/XI0_10/d__5_ DECAP_INV_G11
XG4094 XI11_6/XI0/XI0_10/d_4_ XI11_6/XI0/XI0_10/d__4_ DECAP_INV_G11
XG4095 XI11_6/XI0/XI0_10/d_3_ XI11_6/XI0/XI0_10/d__3_ DECAP_INV_G11
XG4096 XI11_6/XI0/XI0_10/d_2_ XI11_6/XI0/XI0_10/d__2_ DECAP_INV_G11
XG4097 XI11_6/XI0/XI0_10/d_1_ XI11_6/XI0/XI0_10/d__1_ DECAP_INV_G11
XG4098 XI11_6/XI0/XI0_10/d_0_ XI11_6/XI0/XI0_10/d__0_ DECAP_INV_G11
XG4099 XI11_6/XI0/XI0_9/d__15_ XI11_6/XI0/XI0_9/d_15_ DECAP_INV_G11
XG4100 XI11_6/XI0/XI0_9/d__14_ XI11_6/XI0/XI0_9/d_14_ DECAP_INV_G11
XG4101 XI11_6/XI0/XI0_9/d__13_ XI11_6/XI0/XI0_9/d_13_ DECAP_INV_G11
XG4102 XI11_6/XI0/XI0_9/d__12_ XI11_6/XI0/XI0_9/d_12_ DECAP_INV_G11
XG4103 XI11_6/XI0/XI0_9/d__11_ XI11_6/XI0/XI0_9/d_11_ DECAP_INV_G11
XG4104 XI11_6/XI0/XI0_9/d__10_ XI11_6/XI0/XI0_9/d_10_ DECAP_INV_G11
XG4105 XI11_6/XI0/XI0_9/d__9_ XI11_6/XI0/XI0_9/d_9_ DECAP_INV_G11
XG4106 XI11_6/XI0/XI0_9/d__8_ XI11_6/XI0/XI0_9/d_8_ DECAP_INV_G11
XG4107 XI11_6/XI0/XI0_9/d__7_ XI11_6/XI0/XI0_9/d_7_ DECAP_INV_G11
XG4108 XI11_6/XI0/XI0_9/d__6_ XI11_6/XI0/XI0_9/d_6_ DECAP_INV_G11
XG4109 XI11_6/XI0/XI0_9/d__5_ XI11_6/XI0/XI0_9/d_5_ DECAP_INV_G11
XG4110 XI11_6/XI0/XI0_9/d__4_ XI11_6/XI0/XI0_9/d_4_ DECAP_INV_G11
XG4111 XI11_6/XI0/XI0_9/d__3_ XI11_6/XI0/XI0_9/d_3_ DECAP_INV_G11
XG4112 XI11_6/XI0/XI0_9/d__2_ XI11_6/XI0/XI0_9/d_2_ DECAP_INV_G11
XG4113 XI11_6/XI0/XI0_9/d__1_ XI11_6/XI0/XI0_9/d_1_ DECAP_INV_G11
XG4114 XI11_6/XI0/XI0_9/d__0_ XI11_6/XI0/XI0_9/d_0_ DECAP_INV_G11
XG4115 XI11_6/XI0/XI0_9/d_15_ XI11_6/XI0/XI0_9/d__15_ DECAP_INV_G11
XG4116 XI11_6/XI0/XI0_9/d_14_ XI11_6/XI0/XI0_9/d__14_ DECAP_INV_G11
XG4117 XI11_6/XI0/XI0_9/d_13_ XI11_6/XI0/XI0_9/d__13_ DECAP_INV_G11
XG4118 XI11_6/XI0/XI0_9/d_12_ XI11_6/XI0/XI0_9/d__12_ DECAP_INV_G11
XG4119 XI11_6/XI0/XI0_9/d_11_ XI11_6/XI0/XI0_9/d__11_ DECAP_INV_G11
XG4120 XI11_6/XI0/XI0_9/d_10_ XI11_6/XI0/XI0_9/d__10_ DECAP_INV_G11
XG4121 XI11_6/XI0/XI0_9/d_9_ XI11_6/XI0/XI0_9/d__9_ DECAP_INV_G11
XG4122 XI11_6/XI0/XI0_9/d_8_ XI11_6/XI0/XI0_9/d__8_ DECAP_INV_G11
XG4123 XI11_6/XI0/XI0_9/d_7_ XI11_6/XI0/XI0_9/d__7_ DECAP_INV_G11
XG4124 XI11_6/XI0/XI0_9/d_6_ XI11_6/XI0/XI0_9/d__6_ DECAP_INV_G11
XG4125 XI11_6/XI0/XI0_9/d_5_ XI11_6/XI0/XI0_9/d__5_ DECAP_INV_G11
XG4126 XI11_6/XI0/XI0_9/d_4_ XI11_6/XI0/XI0_9/d__4_ DECAP_INV_G11
XG4127 XI11_6/XI0/XI0_9/d_3_ XI11_6/XI0/XI0_9/d__3_ DECAP_INV_G11
XG4128 XI11_6/XI0/XI0_9/d_2_ XI11_6/XI0/XI0_9/d__2_ DECAP_INV_G11
XG4129 XI11_6/XI0/XI0_9/d_1_ XI11_6/XI0/XI0_9/d__1_ DECAP_INV_G11
XG4130 XI11_6/XI0/XI0_9/d_0_ XI11_6/XI0/XI0_9/d__0_ DECAP_INV_G11
XG4131 XI11_6/XI0/XI0_8/d__15_ XI11_6/XI0/XI0_8/d_15_ DECAP_INV_G11
XG4132 XI11_6/XI0/XI0_8/d__14_ XI11_6/XI0/XI0_8/d_14_ DECAP_INV_G11
XG4133 XI11_6/XI0/XI0_8/d__13_ XI11_6/XI0/XI0_8/d_13_ DECAP_INV_G11
XG4134 XI11_6/XI0/XI0_8/d__12_ XI11_6/XI0/XI0_8/d_12_ DECAP_INV_G11
XG4135 XI11_6/XI0/XI0_8/d__11_ XI11_6/XI0/XI0_8/d_11_ DECAP_INV_G11
XG4136 XI11_6/XI0/XI0_8/d__10_ XI11_6/XI0/XI0_8/d_10_ DECAP_INV_G11
XG4137 XI11_6/XI0/XI0_8/d__9_ XI11_6/XI0/XI0_8/d_9_ DECAP_INV_G11
XG4138 XI11_6/XI0/XI0_8/d__8_ XI11_6/XI0/XI0_8/d_8_ DECAP_INV_G11
XG4139 XI11_6/XI0/XI0_8/d__7_ XI11_6/XI0/XI0_8/d_7_ DECAP_INV_G11
XG4140 XI11_6/XI0/XI0_8/d__6_ XI11_6/XI0/XI0_8/d_6_ DECAP_INV_G11
XG4141 XI11_6/XI0/XI0_8/d__5_ XI11_6/XI0/XI0_8/d_5_ DECAP_INV_G11
XG4142 XI11_6/XI0/XI0_8/d__4_ XI11_6/XI0/XI0_8/d_4_ DECAP_INV_G11
XG4143 XI11_6/XI0/XI0_8/d__3_ XI11_6/XI0/XI0_8/d_3_ DECAP_INV_G11
XG4144 XI11_6/XI0/XI0_8/d__2_ XI11_6/XI0/XI0_8/d_2_ DECAP_INV_G11
XG4145 XI11_6/XI0/XI0_8/d__1_ XI11_6/XI0/XI0_8/d_1_ DECAP_INV_G11
XG4146 XI11_6/XI0/XI0_8/d__0_ XI11_6/XI0/XI0_8/d_0_ DECAP_INV_G11
XG4147 XI11_6/XI0/XI0_8/d_15_ XI11_6/XI0/XI0_8/d__15_ DECAP_INV_G11
XG4148 XI11_6/XI0/XI0_8/d_14_ XI11_6/XI0/XI0_8/d__14_ DECAP_INV_G11
XG4149 XI11_6/XI0/XI0_8/d_13_ XI11_6/XI0/XI0_8/d__13_ DECAP_INV_G11
XG4150 XI11_6/XI0/XI0_8/d_12_ XI11_6/XI0/XI0_8/d__12_ DECAP_INV_G11
XG4151 XI11_6/XI0/XI0_8/d_11_ XI11_6/XI0/XI0_8/d__11_ DECAP_INV_G11
XG4152 XI11_6/XI0/XI0_8/d_10_ XI11_6/XI0/XI0_8/d__10_ DECAP_INV_G11
XG4153 XI11_6/XI0/XI0_8/d_9_ XI11_6/XI0/XI0_8/d__9_ DECAP_INV_G11
XG4154 XI11_6/XI0/XI0_8/d_8_ XI11_6/XI0/XI0_8/d__8_ DECAP_INV_G11
XG4155 XI11_6/XI0/XI0_8/d_7_ XI11_6/XI0/XI0_8/d__7_ DECAP_INV_G11
XG4156 XI11_6/XI0/XI0_8/d_6_ XI11_6/XI0/XI0_8/d__6_ DECAP_INV_G11
XG4157 XI11_6/XI0/XI0_8/d_5_ XI11_6/XI0/XI0_8/d__5_ DECAP_INV_G11
XG4158 XI11_6/XI0/XI0_8/d_4_ XI11_6/XI0/XI0_8/d__4_ DECAP_INV_G11
XG4159 XI11_6/XI0/XI0_8/d_3_ XI11_6/XI0/XI0_8/d__3_ DECAP_INV_G11
XG4160 XI11_6/XI0/XI0_8/d_2_ XI11_6/XI0/XI0_8/d__2_ DECAP_INV_G11
XG4161 XI11_6/XI0/XI0_8/d_1_ XI11_6/XI0/XI0_8/d__1_ DECAP_INV_G11
XG4162 XI11_6/XI0/XI0_8/d_0_ XI11_6/XI0/XI0_8/d__0_ DECAP_INV_G11
XG4163 XI11_6/XI0/XI0_7/d__15_ XI11_6/XI0/XI0_7/d_15_ DECAP_INV_G11
XG4164 XI11_6/XI0/XI0_7/d__14_ XI11_6/XI0/XI0_7/d_14_ DECAP_INV_G11
XG4165 XI11_6/XI0/XI0_7/d__13_ XI11_6/XI0/XI0_7/d_13_ DECAP_INV_G11
XG4166 XI11_6/XI0/XI0_7/d__12_ XI11_6/XI0/XI0_7/d_12_ DECAP_INV_G11
XG4167 XI11_6/XI0/XI0_7/d__11_ XI11_6/XI0/XI0_7/d_11_ DECAP_INV_G11
XG4168 XI11_6/XI0/XI0_7/d__10_ XI11_6/XI0/XI0_7/d_10_ DECAP_INV_G11
XG4169 XI11_6/XI0/XI0_7/d__9_ XI11_6/XI0/XI0_7/d_9_ DECAP_INV_G11
XG4170 XI11_6/XI0/XI0_7/d__8_ XI11_6/XI0/XI0_7/d_8_ DECAP_INV_G11
XG4171 XI11_6/XI0/XI0_7/d__7_ XI11_6/XI0/XI0_7/d_7_ DECAP_INV_G11
XG4172 XI11_6/XI0/XI0_7/d__6_ XI11_6/XI0/XI0_7/d_6_ DECAP_INV_G11
XG4173 XI11_6/XI0/XI0_7/d__5_ XI11_6/XI0/XI0_7/d_5_ DECAP_INV_G11
XG4174 XI11_6/XI0/XI0_7/d__4_ XI11_6/XI0/XI0_7/d_4_ DECAP_INV_G11
XG4175 XI11_6/XI0/XI0_7/d__3_ XI11_6/XI0/XI0_7/d_3_ DECAP_INV_G11
XG4176 XI11_6/XI0/XI0_7/d__2_ XI11_6/XI0/XI0_7/d_2_ DECAP_INV_G11
XG4177 XI11_6/XI0/XI0_7/d__1_ XI11_6/XI0/XI0_7/d_1_ DECAP_INV_G11
XG4178 XI11_6/XI0/XI0_7/d__0_ XI11_6/XI0/XI0_7/d_0_ DECAP_INV_G11
XG4179 XI11_6/XI0/XI0_7/d_15_ XI11_6/XI0/XI0_7/d__15_ DECAP_INV_G11
XG4180 XI11_6/XI0/XI0_7/d_14_ XI11_6/XI0/XI0_7/d__14_ DECAP_INV_G11
XG4181 XI11_6/XI0/XI0_7/d_13_ XI11_6/XI0/XI0_7/d__13_ DECAP_INV_G11
XG4182 XI11_6/XI0/XI0_7/d_12_ XI11_6/XI0/XI0_7/d__12_ DECAP_INV_G11
XG4183 XI11_6/XI0/XI0_7/d_11_ XI11_6/XI0/XI0_7/d__11_ DECAP_INV_G11
XG4184 XI11_6/XI0/XI0_7/d_10_ XI11_6/XI0/XI0_7/d__10_ DECAP_INV_G11
XG4185 XI11_6/XI0/XI0_7/d_9_ XI11_6/XI0/XI0_7/d__9_ DECAP_INV_G11
XG4186 XI11_6/XI0/XI0_7/d_8_ XI11_6/XI0/XI0_7/d__8_ DECAP_INV_G11
XG4187 XI11_6/XI0/XI0_7/d_7_ XI11_6/XI0/XI0_7/d__7_ DECAP_INV_G11
XG4188 XI11_6/XI0/XI0_7/d_6_ XI11_6/XI0/XI0_7/d__6_ DECAP_INV_G11
XG4189 XI11_6/XI0/XI0_7/d_5_ XI11_6/XI0/XI0_7/d__5_ DECAP_INV_G11
XG4190 XI11_6/XI0/XI0_7/d_4_ XI11_6/XI0/XI0_7/d__4_ DECAP_INV_G11
XG4191 XI11_6/XI0/XI0_7/d_3_ XI11_6/XI0/XI0_7/d__3_ DECAP_INV_G11
XG4192 XI11_6/XI0/XI0_7/d_2_ XI11_6/XI0/XI0_7/d__2_ DECAP_INV_G11
XG4193 XI11_6/XI0/XI0_7/d_1_ XI11_6/XI0/XI0_7/d__1_ DECAP_INV_G11
XG4194 XI11_6/XI0/XI0_7/d_0_ XI11_6/XI0/XI0_7/d__0_ DECAP_INV_G11
XG4195 XI11_6/XI0/XI0_6/d__15_ XI11_6/XI0/XI0_6/d_15_ DECAP_INV_G11
XG4196 XI11_6/XI0/XI0_6/d__14_ XI11_6/XI0/XI0_6/d_14_ DECAP_INV_G11
XG4197 XI11_6/XI0/XI0_6/d__13_ XI11_6/XI0/XI0_6/d_13_ DECAP_INV_G11
XG4198 XI11_6/XI0/XI0_6/d__12_ XI11_6/XI0/XI0_6/d_12_ DECAP_INV_G11
XG4199 XI11_6/XI0/XI0_6/d__11_ XI11_6/XI0/XI0_6/d_11_ DECAP_INV_G11
XG4200 XI11_6/XI0/XI0_6/d__10_ XI11_6/XI0/XI0_6/d_10_ DECAP_INV_G11
XG4201 XI11_6/XI0/XI0_6/d__9_ XI11_6/XI0/XI0_6/d_9_ DECAP_INV_G11
XG4202 XI11_6/XI0/XI0_6/d__8_ XI11_6/XI0/XI0_6/d_8_ DECAP_INV_G11
XG4203 XI11_6/XI0/XI0_6/d__7_ XI11_6/XI0/XI0_6/d_7_ DECAP_INV_G11
XG4204 XI11_6/XI0/XI0_6/d__6_ XI11_6/XI0/XI0_6/d_6_ DECAP_INV_G11
XG4205 XI11_6/XI0/XI0_6/d__5_ XI11_6/XI0/XI0_6/d_5_ DECAP_INV_G11
XG4206 XI11_6/XI0/XI0_6/d__4_ XI11_6/XI0/XI0_6/d_4_ DECAP_INV_G11
XG4207 XI11_6/XI0/XI0_6/d__3_ XI11_6/XI0/XI0_6/d_3_ DECAP_INV_G11
XG4208 XI11_6/XI0/XI0_6/d__2_ XI11_6/XI0/XI0_6/d_2_ DECAP_INV_G11
XG4209 XI11_6/XI0/XI0_6/d__1_ XI11_6/XI0/XI0_6/d_1_ DECAP_INV_G11
XG4210 XI11_6/XI0/XI0_6/d__0_ XI11_6/XI0/XI0_6/d_0_ DECAP_INV_G11
XG4211 XI11_6/XI0/XI0_6/d_15_ XI11_6/XI0/XI0_6/d__15_ DECAP_INV_G11
XG4212 XI11_6/XI0/XI0_6/d_14_ XI11_6/XI0/XI0_6/d__14_ DECAP_INV_G11
XG4213 XI11_6/XI0/XI0_6/d_13_ XI11_6/XI0/XI0_6/d__13_ DECAP_INV_G11
XG4214 XI11_6/XI0/XI0_6/d_12_ XI11_6/XI0/XI0_6/d__12_ DECAP_INV_G11
XG4215 XI11_6/XI0/XI0_6/d_11_ XI11_6/XI0/XI0_6/d__11_ DECAP_INV_G11
XG4216 XI11_6/XI0/XI0_6/d_10_ XI11_6/XI0/XI0_6/d__10_ DECAP_INV_G11
XG4217 XI11_6/XI0/XI0_6/d_9_ XI11_6/XI0/XI0_6/d__9_ DECAP_INV_G11
XG4218 XI11_6/XI0/XI0_6/d_8_ XI11_6/XI0/XI0_6/d__8_ DECAP_INV_G11
XG4219 XI11_6/XI0/XI0_6/d_7_ XI11_6/XI0/XI0_6/d__7_ DECAP_INV_G11
XG4220 XI11_6/XI0/XI0_6/d_6_ XI11_6/XI0/XI0_6/d__6_ DECAP_INV_G11
XG4221 XI11_6/XI0/XI0_6/d_5_ XI11_6/XI0/XI0_6/d__5_ DECAP_INV_G11
XG4222 XI11_6/XI0/XI0_6/d_4_ XI11_6/XI0/XI0_6/d__4_ DECAP_INV_G11
XG4223 XI11_6/XI0/XI0_6/d_3_ XI11_6/XI0/XI0_6/d__3_ DECAP_INV_G11
XG4224 XI11_6/XI0/XI0_6/d_2_ XI11_6/XI0/XI0_6/d__2_ DECAP_INV_G11
XG4225 XI11_6/XI0/XI0_6/d_1_ XI11_6/XI0/XI0_6/d__1_ DECAP_INV_G11
XG4226 XI11_6/XI0/XI0_6/d_0_ XI11_6/XI0/XI0_6/d__0_ DECAP_INV_G11
XG4227 XI11_6/XI0/XI0_5/d__15_ XI11_6/XI0/XI0_5/d_15_ DECAP_INV_G11
XG4228 XI11_6/XI0/XI0_5/d__14_ XI11_6/XI0/XI0_5/d_14_ DECAP_INV_G11
XG4229 XI11_6/XI0/XI0_5/d__13_ XI11_6/XI0/XI0_5/d_13_ DECAP_INV_G11
XG4230 XI11_6/XI0/XI0_5/d__12_ XI11_6/XI0/XI0_5/d_12_ DECAP_INV_G11
XG4231 XI11_6/XI0/XI0_5/d__11_ XI11_6/XI0/XI0_5/d_11_ DECAP_INV_G11
XG4232 XI11_6/XI0/XI0_5/d__10_ XI11_6/XI0/XI0_5/d_10_ DECAP_INV_G11
XG4233 XI11_6/XI0/XI0_5/d__9_ XI11_6/XI0/XI0_5/d_9_ DECAP_INV_G11
XG4234 XI11_6/XI0/XI0_5/d__8_ XI11_6/XI0/XI0_5/d_8_ DECAP_INV_G11
XG4235 XI11_6/XI0/XI0_5/d__7_ XI11_6/XI0/XI0_5/d_7_ DECAP_INV_G11
XG4236 XI11_6/XI0/XI0_5/d__6_ XI11_6/XI0/XI0_5/d_6_ DECAP_INV_G11
XG4237 XI11_6/XI0/XI0_5/d__5_ XI11_6/XI0/XI0_5/d_5_ DECAP_INV_G11
XG4238 XI11_6/XI0/XI0_5/d__4_ XI11_6/XI0/XI0_5/d_4_ DECAP_INV_G11
XG4239 XI11_6/XI0/XI0_5/d__3_ XI11_6/XI0/XI0_5/d_3_ DECAP_INV_G11
XG4240 XI11_6/XI0/XI0_5/d__2_ XI11_6/XI0/XI0_5/d_2_ DECAP_INV_G11
XG4241 XI11_6/XI0/XI0_5/d__1_ XI11_6/XI0/XI0_5/d_1_ DECAP_INV_G11
XG4242 XI11_6/XI0/XI0_5/d__0_ XI11_6/XI0/XI0_5/d_0_ DECAP_INV_G11
XG4243 XI11_6/XI0/XI0_5/d_15_ XI11_6/XI0/XI0_5/d__15_ DECAP_INV_G11
XG4244 XI11_6/XI0/XI0_5/d_14_ XI11_6/XI0/XI0_5/d__14_ DECAP_INV_G11
XG4245 XI11_6/XI0/XI0_5/d_13_ XI11_6/XI0/XI0_5/d__13_ DECAP_INV_G11
XG4246 XI11_6/XI0/XI0_5/d_12_ XI11_6/XI0/XI0_5/d__12_ DECAP_INV_G11
XG4247 XI11_6/XI0/XI0_5/d_11_ XI11_6/XI0/XI0_5/d__11_ DECAP_INV_G11
XG4248 XI11_6/XI0/XI0_5/d_10_ XI11_6/XI0/XI0_5/d__10_ DECAP_INV_G11
XG4249 XI11_6/XI0/XI0_5/d_9_ XI11_6/XI0/XI0_5/d__9_ DECAP_INV_G11
XG4250 XI11_6/XI0/XI0_5/d_8_ XI11_6/XI0/XI0_5/d__8_ DECAP_INV_G11
XG4251 XI11_6/XI0/XI0_5/d_7_ XI11_6/XI0/XI0_5/d__7_ DECAP_INV_G11
XG4252 XI11_6/XI0/XI0_5/d_6_ XI11_6/XI0/XI0_5/d__6_ DECAP_INV_G11
XG4253 XI11_6/XI0/XI0_5/d_5_ XI11_6/XI0/XI0_5/d__5_ DECAP_INV_G11
XG4254 XI11_6/XI0/XI0_5/d_4_ XI11_6/XI0/XI0_5/d__4_ DECAP_INV_G11
XG4255 XI11_6/XI0/XI0_5/d_3_ XI11_6/XI0/XI0_5/d__3_ DECAP_INV_G11
XG4256 XI11_6/XI0/XI0_5/d_2_ XI11_6/XI0/XI0_5/d__2_ DECAP_INV_G11
XG4257 XI11_6/XI0/XI0_5/d_1_ XI11_6/XI0/XI0_5/d__1_ DECAP_INV_G11
XG4258 XI11_6/XI0/XI0_5/d_0_ XI11_6/XI0/XI0_5/d__0_ DECAP_INV_G11
XG4259 XI11_6/XI0/XI0_4/d__15_ XI11_6/XI0/XI0_4/d_15_ DECAP_INV_G11
XG4260 XI11_6/XI0/XI0_4/d__14_ XI11_6/XI0/XI0_4/d_14_ DECAP_INV_G11
XG4261 XI11_6/XI0/XI0_4/d__13_ XI11_6/XI0/XI0_4/d_13_ DECAP_INV_G11
XG4262 XI11_6/XI0/XI0_4/d__12_ XI11_6/XI0/XI0_4/d_12_ DECAP_INV_G11
XG4263 XI11_6/XI0/XI0_4/d__11_ XI11_6/XI0/XI0_4/d_11_ DECAP_INV_G11
XG4264 XI11_6/XI0/XI0_4/d__10_ XI11_6/XI0/XI0_4/d_10_ DECAP_INV_G11
XG4265 XI11_6/XI0/XI0_4/d__9_ XI11_6/XI0/XI0_4/d_9_ DECAP_INV_G11
XG4266 XI11_6/XI0/XI0_4/d__8_ XI11_6/XI0/XI0_4/d_8_ DECAP_INV_G11
XG4267 XI11_6/XI0/XI0_4/d__7_ XI11_6/XI0/XI0_4/d_7_ DECAP_INV_G11
XG4268 XI11_6/XI0/XI0_4/d__6_ XI11_6/XI0/XI0_4/d_6_ DECAP_INV_G11
XG4269 XI11_6/XI0/XI0_4/d__5_ XI11_6/XI0/XI0_4/d_5_ DECAP_INV_G11
XG4270 XI11_6/XI0/XI0_4/d__4_ XI11_6/XI0/XI0_4/d_4_ DECAP_INV_G11
XG4271 XI11_6/XI0/XI0_4/d__3_ XI11_6/XI0/XI0_4/d_3_ DECAP_INV_G11
XG4272 XI11_6/XI0/XI0_4/d__2_ XI11_6/XI0/XI0_4/d_2_ DECAP_INV_G11
XG4273 XI11_6/XI0/XI0_4/d__1_ XI11_6/XI0/XI0_4/d_1_ DECAP_INV_G11
XG4274 XI11_6/XI0/XI0_4/d__0_ XI11_6/XI0/XI0_4/d_0_ DECAP_INV_G11
XG4275 XI11_6/XI0/XI0_4/d_15_ XI11_6/XI0/XI0_4/d__15_ DECAP_INV_G11
XG4276 XI11_6/XI0/XI0_4/d_14_ XI11_6/XI0/XI0_4/d__14_ DECAP_INV_G11
XG4277 XI11_6/XI0/XI0_4/d_13_ XI11_6/XI0/XI0_4/d__13_ DECAP_INV_G11
XG4278 XI11_6/XI0/XI0_4/d_12_ XI11_6/XI0/XI0_4/d__12_ DECAP_INV_G11
XG4279 XI11_6/XI0/XI0_4/d_11_ XI11_6/XI0/XI0_4/d__11_ DECAP_INV_G11
XG4280 XI11_6/XI0/XI0_4/d_10_ XI11_6/XI0/XI0_4/d__10_ DECAP_INV_G11
XG4281 XI11_6/XI0/XI0_4/d_9_ XI11_6/XI0/XI0_4/d__9_ DECAP_INV_G11
XG4282 XI11_6/XI0/XI0_4/d_8_ XI11_6/XI0/XI0_4/d__8_ DECAP_INV_G11
XG4283 XI11_6/XI0/XI0_4/d_7_ XI11_6/XI0/XI0_4/d__7_ DECAP_INV_G11
XG4284 XI11_6/XI0/XI0_4/d_6_ XI11_6/XI0/XI0_4/d__6_ DECAP_INV_G11
XG4285 XI11_6/XI0/XI0_4/d_5_ XI11_6/XI0/XI0_4/d__5_ DECAP_INV_G11
XG4286 XI11_6/XI0/XI0_4/d_4_ XI11_6/XI0/XI0_4/d__4_ DECAP_INV_G11
XG4287 XI11_6/XI0/XI0_4/d_3_ XI11_6/XI0/XI0_4/d__3_ DECAP_INV_G11
XG4288 XI11_6/XI0/XI0_4/d_2_ XI11_6/XI0/XI0_4/d__2_ DECAP_INV_G11
XG4289 XI11_6/XI0/XI0_4/d_1_ XI11_6/XI0/XI0_4/d__1_ DECAP_INV_G11
XG4290 XI11_6/XI0/XI0_4/d_0_ XI11_6/XI0/XI0_4/d__0_ DECAP_INV_G11
XG4291 XI11_6/XI0/XI0_3/d__15_ XI11_6/XI0/XI0_3/d_15_ DECAP_INV_G11
XG4292 XI11_6/XI0/XI0_3/d__14_ XI11_6/XI0/XI0_3/d_14_ DECAP_INV_G11
XG4293 XI11_6/XI0/XI0_3/d__13_ XI11_6/XI0/XI0_3/d_13_ DECAP_INV_G11
XG4294 XI11_6/XI0/XI0_3/d__12_ XI11_6/XI0/XI0_3/d_12_ DECAP_INV_G11
XG4295 XI11_6/XI0/XI0_3/d__11_ XI11_6/XI0/XI0_3/d_11_ DECAP_INV_G11
XG4296 XI11_6/XI0/XI0_3/d__10_ XI11_6/XI0/XI0_3/d_10_ DECAP_INV_G11
XG4297 XI11_6/XI0/XI0_3/d__9_ XI11_6/XI0/XI0_3/d_9_ DECAP_INV_G11
XG4298 XI11_6/XI0/XI0_3/d__8_ XI11_6/XI0/XI0_3/d_8_ DECAP_INV_G11
XG4299 XI11_6/XI0/XI0_3/d__7_ XI11_6/XI0/XI0_3/d_7_ DECAP_INV_G11
XG4300 XI11_6/XI0/XI0_3/d__6_ XI11_6/XI0/XI0_3/d_6_ DECAP_INV_G11
XG4301 XI11_6/XI0/XI0_3/d__5_ XI11_6/XI0/XI0_3/d_5_ DECAP_INV_G11
XG4302 XI11_6/XI0/XI0_3/d__4_ XI11_6/XI0/XI0_3/d_4_ DECAP_INV_G11
XG4303 XI11_6/XI0/XI0_3/d__3_ XI11_6/XI0/XI0_3/d_3_ DECAP_INV_G11
XG4304 XI11_6/XI0/XI0_3/d__2_ XI11_6/XI0/XI0_3/d_2_ DECAP_INV_G11
XG4305 XI11_6/XI0/XI0_3/d__1_ XI11_6/XI0/XI0_3/d_1_ DECAP_INV_G11
XG4306 XI11_6/XI0/XI0_3/d__0_ XI11_6/XI0/XI0_3/d_0_ DECAP_INV_G11
XG4307 XI11_6/XI0/XI0_3/d_15_ XI11_6/XI0/XI0_3/d__15_ DECAP_INV_G11
XG4308 XI11_6/XI0/XI0_3/d_14_ XI11_6/XI0/XI0_3/d__14_ DECAP_INV_G11
XG4309 XI11_6/XI0/XI0_3/d_13_ XI11_6/XI0/XI0_3/d__13_ DECAP_INV_G11
XG4310 XI11_6/XI0/XI0_3/d_12_ XI11_6/XI0/XI0_3/d__12_ DECAP_INV_G11
XG4311 XI11_6/XI0/XI0_3/d_11_ XI11_6/XI0/XI0_3/d__11_ DECAP_INV_G11
XG4312 XI11_6/XI0/XI0_3/d_10_ XI11_6/XI0/XI0_3/d__10_ DECAP_INV_G11
XG4313 XI11_6/XI0/XI0_3/d_9_ XI11_6/XI0/XI0_3/d__9_ DECAP_INV_G11
XG4314 XI11_6/XI0/XI0_3/d_8_ XI11_6/XI0/XI0_3/d__8_ DECAP_INV_G11
XG4315 XI11_6/XI0/XI0_3/d_7_ XI11_6/XI0/XI0_3/d__7_ DECAP_INV_G11
XG4316 XI11_6/XI0/XI0_3/d_6_ XI11_6/XI0/XI0_3/d__6_ DECAP_INV_G11
XG4317 XI11_6/XI0/XI0_3/d_5_ XI11_6/XI0/XI0_3/d__5_ DECAP_INV_G11
XG4318 XI11_6/XI0/XI0_3/d_4_ XI11_6/XI0/XI0_3/d__4_ DECAP_INV_G11
XG4319 XI11_6/XI0/XI0_3/d_3_ XI11_6/XI0/XI0_3/d__3_ DECAP_INV_G11
XG4320 XI11_6/XI0/XI0_3/d_2_ XI11_6/XI0/XI0_3/d__2_ DECAP_INV_G11
XG4321 XI11_6/XI0/XI0_3/d_1_ XI11_6/XI0/XI0_3/d__1_ DECAP_INV_G11
XG4322 XI11_6/XI0/XI0_3/d_0_ XI11_6/XI0/XI0_3/d__0_ DECAP_INV_G11
XG4323 XI11_6/XI0/XI0_2/d__15_ XI11_6/XI0/XI0_2/d_15_ DECAP_INV_G11
XG4324 XI11_6/XI0/XI0_2/d__14_ XI11_6/XI0/XI0_2/d_14_ DECAP_INV_G11
XG4325 XI11_6/XI0/XI0_2/d__13_ XI11_6/XI0/XI0_2/d_13_ DECAP_INV_G11
XG4326 XI11_6/XI0/XI0_2/d__12_ XI11_6/XI0/XI0_2/d_12_ DECAP_INV_G11
XG4327 XI11_6/XI0/XI0_2/d__11_ XI11_6/XI0/XI0_2/d_11_ DECAP_INV_G11
XG4328 XI11_6/XI0/XI0_2/d__10_ XI11_6/XI0/XI0_2/d_10_ DECAP_INV_G11
XG4329 XI11_6/XI0/XI0_2/d__9_ XI11_6/XI0/XI0_2/d_9_ DECAP_INV_G11
XG4330 XI11_6/XI0/XI0_2/d__8_ XI11_6/XI0/XI0_2/d_8_ DECAP_INV_G11
XG4331 XI11_6/XI0/XI0_2/d__7_ XI11_6/XI0/XI0_2/d_7_ DECAP_INV_G11
XG4332 XI11_6/XI0/XI0_2/d__6_ XI11_6/XI0/XI0_2/d_6_ DECAP_INV_G11
XG4333 XI11_6/XI0/XI0_2/d__5_ XI11_6/XI0/XI0_2/d_5_ DECAP_INV_G11
XG4334 XI11_6/XI0/XI0_2/d__4_ XI11_6/XI0/XI0_2/d_4_ DECAP_INV_G11
XG4335 XI11_6/XI0/XI0_2/d__3_ XI11_6/XI0/XI0_2/d_3_ DECAP_INV_G11
XG4336 XI11_6/XI0/XI0_2/d__2_ XI11_6/XI0/XI0_2/d_2_ DECAP_INV_G11
XG4337 XI11_6/XI0/XI0_2/d__1_ XI11_6/XI0/XI0_2/d_1_ DECAP_INV_G11
XG4338 XI11_6/XI0/XI0_2/d__0_ XI11_6/XI0/XI0_2/d_0_ DECAP_INV_G11
XG4339 XI11_6/XI0/XI0_2/d_15_ XI11_6/XI0/XI0_2/d__15_ DECAP_INV_G11
XG4340 XI11_6/XI0/XI0_2/d_14_ XI11_6/XI0/XI0_2/d__14_ DECAP_INV_G11
XG4341 XI11_6/XI0/XI0_2/d_13_ XI11_6/XI0/XI0_2/d__13_ DECAP_INV_G11
XG4342 XI11_6/XI0/XI0_2/d_12_ XI11_6/XI0/XI0_2/d__12_ DECAP_INV_G11
XG4343 XI11_6/XI0/XI0_2/d_11_ XI11_6/XI0/XI0_2/d__11_ DECAP_INV_G11
XG4344 XI11_6/XI0/XI0_2/d_10_ XI11_6/XI0/XI0_2/d__10_ DECAP_INV_G11
XG4345 XI11_6/XI0/XI0_2/d_9_ XI11_6/XI0/XI0_2/d__9_ DECAP_INV_G11
XG4346 XI11_6/XI0/XI0_2/d_8_ XI11_6/XI0/XI0_2/d__8_ DECAP_INV_G11
XG4347 XI11_6/XI0/XI0_2/d_7_ XI11_6/XI0/XI0_2/d__7_ DECAP_INV_G11
XG4348 XI11_6/XI0/XI0_2/d_6_ XI11_6/XI0/XI0_2/d__6_ DECAP_INV_G11
XG4349 XI11_6/XI0/XI0_2/d_5_ XI11_6/XI0/XI0_2/d__5_ DECAP_INV_G11
XG4350 XI11_6/XI0/XI0_2/d_4_ XI11_6/XI0/XI0_2/d__4_ DECAP_INV_G11
XG4351 XI11_6/XI0/XI0_2/d_3_ XI11_6/XI0/XI0_2/d__3_ DECAP_INV_G11
XG4352 XI11_6/XI0/XI0_2/d_2_ XI11_6/XI0/XI0_2/d__2_ DECAP_INV_G11
XG4353 XI11_6/XI0/XI0_2/d_1_ XI11_6/XI0/XI0_2/d__1_ DECAP_INV_G11
XG4354 XI11_6/XI0/XI0_2/d_0_ XI11_6/XI0/XI0_2/d__0_ DECAP_INV_G11
XG4355 XI11_6/XI0/XI0_1/d__15_ XI11_6/XI0/XI0_1/d_15_ DECAP_INV_G11
XG4356 XI11_6/XI0/XI0_1/d__14_ XI11_6/XI0/XI0_1/d_14_ DECAP_INV_G11
XG4357 XI11_6/XI0/XI0_1/d__13_ XI11_6/XI0/XI0_1/d_13_ DECAP_INV_G11
XG4358 XI11_6/XI0/XI0_1/d__12_ XI11_6/XI0/XI0_1/d_12_ DECAP_INV_G11
XG4359 XI11_6/XI0/XI0_1/d__11_ XI11_6/XI0/XI0_1/d_11_ DECAP_INV_G11
XG4360 XI11_6/XI0/XI0_1/d__10_ XI11_6/XI0/XI0_1/d_10_ DECAP_INV_G11
XG4361 XI11_6/XI0/XI0_1/d__9_ XI11_6/XI0/XI0_1/d_9_ DECAP_INV_G11
XG4362 XI11_6/XI0/XI0_1/d__8_ XI11_6/XI0/XI0_1/d_8_ DECAP_INV_G11
XG4363 XI11_6/XI0/XI0_1/d__7_ XI11_6/XI0/XI0_1/d_7_ DECAP_INV_G11
XG4364 XI11_6/XI0/XI0_1/d__6_ XI11_6/XI0/XI0_1/d_6_ DECAP_INV_G11
XG4365 XI11_6/XI0/XI0_1/d__5_ XI11_6/XI0/XI0_1/d_5_ DECAP_INV_G11
XG4366 XI11_6/XI0/XI0_1/d__4_ XI11_6/XI0/XI0_1/d_4_ DECAP_INV_G11
XG4367 XI11_6/XI0/XI0_1/d__3_ XI11_6/XI0/XI0_1/d_3_ DECAP_INV_G11
XG4368 XI11_6/XI0/XI0_1/d__2_ XI11_6/XI0/XI0_1/d_2_ DECAP_INV_G11
XG4369 XI11_6/XI0/XI0_1/d__1_ XI11_6/XI0/XI0_1/d_1_ DECAP_INV_G11
XG4370 XI11_6/XI0/XI0_1/d__0_ XI11_6/XI0/XI0_1/d_0_ DECAP_INV_G11
XG4371 XI11_6/XI0/XI0_1/d_15_ XI11_6/XI0/XI0_1/d__15_ DECAP_INV_G11
XG4372 XI11_6/XI0/XI0_1/d_14_ XI11_6/XI0/XI0_1/d__14_ DECAP_INV_G11
XG4373 XI11_6/XI0/XI0_1/d_13_ XI11_6/XI0/XI0_1/d__13_ DECAP_INV_G11
XG4374 XI11_6/XI0/XI0_1/d_12_ XI11_6/XI0/XI0_1/d__12_ DECAP_INV_G11
XG4375 XI11_6/XI0/XI0_1/d_11_ XI11_6/XI0/XI0_1/d__11_ DECAP_INV_G11
XG4376 XI11_6/XI0/XI0_1/d_10_ XI11_6/XI0/XI0_1/d__10_ DECAP_INV_G11
XG4377 XI11_6/XI0/XI0_1/d_9_ XI11_6/XI0/XI0_1/d__9_ DECAP_INV_G11
XG4378 XI11_6/XI0/XI0_1/d_8_ XI11_6/XI0/XI0_1/d__8_ DECAP_INV_G11
XG4379 XI11_6/XI0/XI0_1/d_7_ XI11_6/XI0/XI0_1/d__7_ DECAP_INV_G11
XG4380 XI11_6/XI0/XI0_1/d_6_ XI11_6/XI0/XI0_1/d__6_ DECAP_INV_G11
XG4381 XI11_6/XI0/XI0_1/d_5_ XI11_6/XI0/XI0_1/d__5_ DECAP_INV_G11
XG4382 XI11_6/XI0/XI0_1/d_4_ XI11_6/XI0/XI0_1/d__4_ DECAP_INV_G11
XG4383 XI11_6/XI0/XI0_1/d_3_ XI11_6/XI0/XI0_1/d__3_ DECAP_INV_G11
XG4384 XI11_6/XI0/XI0_1/d_2_ XI11_6/XI0/XI0_1/d__2_ DECAP_INV_G11
XG4385 XI11_6/XI0/XI0_1/d_1_ XI11_6/XI0/XI0_1/d__1_ DECAP_INV_G11
XG4386 XI11_6/XI0/XI0_1/d_0_ XI11_6/XI0/XI0_1/d__0_ DECAP_INV_G11
XG4387 XI11_6/XI0/XI0_0/d__15_ XI11_6/XI0/XI0_0/d_15_ DECAP_INV_G11
XG4388 XI11_6/XI0/XI0_0/d__14_ XI11_6/XI0/XI0_0/d_14_ DECAP_INV_G11
XG4389 XI11_6/XI0/XI0_0/d__13_ XI11_6/XI0/XI0_0/d_13_ DECAP_INV_G11
XG4390 XI11_6/XI0/XI0_0/d__12_ XI11_6/XI0/XI0_0/d_12_ DECAP_INV_G11
XG4391 XI11_6/XI0/XI0_0/d__11_ XI11_6/XI0/XI0_0/d_11_ DECAP_INV_G11
XG4392 XI11_6/XI0/XI0_0/d__10_ XI11_6/XI0/XI0_0/d_10_ DECAP_INV_G11
XG4393 XI11_6/XI0/XI0_0/d__9_ XI11_6/XI0/XI0_0/d_9_ DECAP_INV_G11
XG4394 XI11_6/XI0/XI0_0/d__8_ XI11_6/XI0/XI0_0/d_8_ DECAP_INV_G11
XG4395 XI11_6/XI0/XI0_0/d__7_ XI11_6/XI0/XI0_0/d_7_ DECAP_INV_G11
XG4396 XI11_6/XI0/XI0_0/d__6_ XI11_6/XI0/XI0_0/d_6_ DECAP_INV_G11
XG4397 XI11_6/XI0/XI0_0/d__5_ XI11_6/XI0/XI0_0/d_5_ DECAP_INV_G11
XG4398 XI11_6/XI0/XI0_0/d__4_ XI11_6/XI0/XI0_0/d_4_ DECAP_INV_G11
XG4399 XI11_6/XI0/XI0_0/d__3_ XI11_6/XI0/XI0_0/d_3_ DECAP_INV_G11
XG4400 XI11_6/XI0/XI0_0/d__2_ XI11_6/XI0/XI0_0/d_2_ DECAP_INV_G11
XG4401 XI11_6/XI0/XI0_0/d__1_ XI11_6/XI0/XI0_0/d_1_ DECAP_INV_G11
XG4402 XI11_6/XI0/XI0_0/d__0_ XI11_6/XI0/XI0_0/d_0_ DECAP_INV_G11
XG4403 XI11_6/XI0/XI0_0/d_15_ XI11_6/XI0/XI0_0/d__15_ DECAP_INV_G11
XG4404 XI11_6/XI0/XI0_0/d_14_ XI11_6/XI0/XI0_0/d__14_ DECAP_INV_G11
XG4405 XI11_6/XI0/XI0_0/d_13_ XI11_6/XI0/XI0_0/d__13_ DECAP_INV_G11
XG4406 XI11_6/XI0/XI0_0/d_12_ XI11_6/XI0/XI0_0/d__12_ DECAP_INV_G11
XG4407 XI11_6/XI0/XI0_0/d_11_ XI11_6/XI0/XI0_0/d__11_ DECAP_INV_G11
XG4408 XI11_6/XI0/XI0_0/d_10_ XI11_6/XI0/XI0_0/d__10_ DECAP_INV_G11
XG4409 XI11_6/XI0/XI0_0/d_9_ XI11_6/XI0/XI0_0/d__9_ DECAP_INV_G11
XG4410 XI11_6/XI0/XI0_0/d_8_ XI11_6/XI0/XI0_0/d__8_ DECAP_INV_G11
XG4411 XI11_6/XI0/XI0_0/d_7_ XI11_6/XI0/XI0_0/d__7_ DECAP_INV_G11
XG4412 XI11_6/XI0/XI0_0/d_6_ XI11_6/XI0/XI0_0/d__6_ DECAP_INV_G11
XG4413 XI11_6/XI0/XI0_0/d_5_ XI11_6/XI0/XI0_0/d__5_ DECAP_INV_G11
XG4414 XI11_6/XI0/XI0_0/d_4_ XI11_6/XI0/XI0_0/d__4_ DECAP_INV_G11
XG4415 XI11_6/XI0/XI0_0/d_3_ XI11_6/XI0/XI0_0/d__3_ DECAP_INV_G11
XG4416 XI11_6/XI0/XI0_0/d_2_ XI11_6/XI0/XI0_0/d__2_ DECAP_INV_G11
XG4417 XI11_6/XI0/XI0_0/d_1_ XI11_6/XI0/XI0_0/d__1_ DECAP_INV_G11
XG4418 XI11_6/XI0/XI0_0/d_0_ XI11_6/XI0/XI0_0/d__0_ DECAP_INV_G11
XG4419 XI11_5/XI3/net17 XI11_5/XI3/net5 DECAP_INV_G7
XG4420 XI11_5/XI3/net5 XI11_5/preck DECAP_INV_G8
XG4421 sck_bar XI11_5/XI3/net018 DECAP_INV_G9
XG4422 XI11_5/XI3/net018 XI11_5/XI3/net012 DECAP_INV_G9
XG4423 XI11_5/XI3/net014 XI11_5/XI3/net7 DECAP_INV_G9
XG4424 XI11_5/XI3/net012 XI11_5/XI3/net014 DECAP_INV_G9
XG4425 XI11_5/XI4/net063 XI11_5/XI4/net0112 DECAP_INV_G10
XG4426 XI11_5/XI4/net26 XI11_5/XI4/net089 DECAP_INV_G10
XG4427 XI11_5/XI4/data_out XI11_5/XI4/data_out_ DECAP_INV_G10
XG4428 XI11_5/XI4/net20 XI11_5/XI4/net0103 DECAP_INV_G10
XG4429 XI11_5/net12 XI11_5/XI4/net32 DECAP_INV_G7
XG4430 XI11_5/net9 XI11_5/XI4/net52 DECAP_INV_G7
XG4431 XI11_5/XI4/data_out_ XI11_5/XI4/data_out DECAP_INV_G10
XG4432 XI11_5/XI0/XI0_63/d__15_ XI11_5/XI0/XI0_63/d_15_ DECAP_INV_G11
XG4433 XI11_5/XI0/XI0_63/d__14_ XI11_5/XI0/XI0_63/d_14_ DECAP_INV_G11
XG4434 XI11_5/XI0/XI0_63/d__13_ XI11_5/XI0/XI0_63/d_13_ DECAP_INV_G11
XG4435 XI11_5/XI0/XI0_63/d__12_ XI11_5/XI0/XI0_63/d_12_ DECAP_INV_G11
XG4436 XI11_5/XI0/XI0_63/d__11_ XI11_5/XI0/XI0_63/d_11_ DECAP_INV_G11
XG4437 XI11_5/XI0/XI0_63/d__10_ XI11_5/XI0/XI0_63/d_10_ DECAP_INV_G11
XG4438 XI11_5/XI0/XI0_63/d__9_ XI11_5/XI0/XI0_63/d_9_ DECAP_INV_G11
XG4439 XI11_5/XI0/XI0_63/d__8_ XI11_5/XI0/XI0_63/d_8_ DECAP_INV_G11
XG4440 XI11_5/XI0/XI0_63/d__7_ XI11_5/XI0/XI0_63/d_7_ DECAP_INV_G11
XG4441 XI11_5/XI0/XI0_63/d__6_ XI11_5/XI0/XI0_63/d_6_ DECAP_INV_G11
XG4442 XI11_5/XI0/XI0_63/d__5_ XI11_5/XI0/XI0_63/d_5_ DECAP_INV_G11
XG4443 XI11_5/XI0/XI0_63/d__4_ XI11_5/XI0/XI0_63/d_4_ DECAP_INV_G11
XG4444 XI11_5/XI0/XI0_63/d__3_ XI11_5/XI0/XI0_63/d_3_ DECAP_INV_G11
XG4445 XI11_5/XI0/XI0_63/d__2_ XI11_5/XI0/XI0_63/d_2_ DECAP_INV_G11
XG4446 XI11_5/XI0/XI0_63/d__1_ XI11_5/XI0/XI0_63/d_1_ DECAP_INV_G11
XG4447 XI11_5/XI0/XI0_63/d__0_ XI11_5/XI0/XI0_63/d_0_ DECAP_INV_G11
XG4448 XI11_5/XI0/XI0_63/d_15_ XI11_5/XI0/XI0_63/d__15_ DECAP_INV_G11
XG4449 XI11_5/XI0/XI0_63/d_14_ XI11_5/XI0/XI0_63/d__14_ DECAP_INV_G11
XG4450 XI11_5/XI0/XI0_63/d_13_ XI11_5/XI0/XI0_63/d__13_ DECAP_INV_G11
XG4451 XI11_5/XI0/XI0_63/d_12_ XI11_5/XI0/XI0_63/d__12_ DECAP_INV_G11
XG4452 XI11_5/XI0/XI0_63/d_11_ XI11_5/XI0/XI0_63/d__11_ DECAP_INV_G11
XG4453 XI11_5/XI0/XI0_63/d_10_ XI11_5/XI0/XI0_63/d__10_ DECAP_INV_G11
XG4454 XI11_5/XI0/XI0_63/d_9_ XI11_5/XI0/XI0_63/d__9_ DECAP_INV_G11
XG4455 XI11_5/XI0/XI0_63/d_8_ XI11_5/XI0/XI0_63/d__8_ DECAP_INV_G11
XG4456 XI11_5/XI0/XI0_63/d_7_ XI11_5/XI0/XI0_63/d__7_ DECAP_INV_G11
XG4457 XI11_5/XI0/XI0_63/d_6_ XI11_5/XI0/XI0_63/d__6_ DECAP_INV_G11
XG4458 XI11_5/XI0/XI0_63/d_5_ XI11_5/XI0/XI0_63/d__5_ DECAP_INV_G11
XG4459 XI11_5/XI0/XI0_63/d_4_ XI11_5/XI0/XI0_63/d__4_ DECAP_INV_G11
XG4460 XI11_5/XI0/XI0_63/d_3_ XI11_5/XI0/XI0_63/d__3_ DECAP_INV_G11
XG4461 XI11_5/XI0/XI0_63/d_2_ XI11_5/XI0/XI0_63/d__2_ DECAP_INV_G11
XG4462 XI11_5/XI0/XI0_63/d_1_ XI11_5/XI0/XI0_63/d__1_ DECAP_INV_G11
XG4463 XI11_5/XI0/XI0_63/d_0_ XI11_5/XI0/XI0_63/d__0_ DECAP_INV_G11
XG4464 XI11_5/XI0/XI0_62/d__15_ XI11_5/XI0/XI0_62/d_15_ DECAP_INV_G11
XG4465 XI11_5/XI0/XI0_62/d__14_ XI11_5/XI0/XI0_62/d_14_ DECAP_INV_G11
XG4466 XI11_5/XI0/XI0_62/d__13_ XI11_5/XI0/XI0_62/d_13_ DECAP_INV_G11
XG4467 XI11_5/XI0/XI0_62/d__12_ XI11_5/XI0/XI0_62/d_12_ DECAP_INV_G11
XG4468 XI11_5/XI0/XI0_62/d__11_ XI11_5/XI0/XI0_62/d_11_ DECAP_INV_G11
XG4469 XI11_5/XI0/XI0_62/d__10_ XI11_5/XI0/XI0_62/d_10_ DECAP_INV_G11
XG4470 XI11_5/XI0/XI0_62/d__9_ XI11_5/XI0/XI0_62/d_9_ DECAP_INV_G11
XG4471 XI11_5/XI0/XI0_62/d__8_ XI11_5/XI0/XI0_62/d_8_ DECAP_INV_G11
XG4472 XI11_5/XI0/XI0_62/d__7_ XI11_5/XI0/XI0_62/d_7_ DECAP_INV_G11
XG4473 XI11_5/XI0/XI0_62/d__6_ XI11_5/XI0/XI0_62/d_6_ DECAP_INV_G11
XG4474 XI11_5/XI0/XI0_62/d__5_ XI11_5/XI0/XI0_62/d_5_ DECAP_INV_G11
XG4475 XI11_5/XI0/XI0_62/d__4_ XI11_5/XI0/XI0_62/d_4_ DECAP_INV_G11
XG4476 XI11_5/XI0/XI0_62/d__3_ XI11_5/XI0/XI0_62/d_3_ DECAP_INV_G11
XG4477 XI11_5/XI0/XI0_62/d__2_ XI11_5/XI0/XI0_62/d_2_ DECAP_INV_G11
XG4478 XI11_5/XI0/XI0_62/d__1_ XI11_5/XI0/XI0_62/d_1_ DECAP_INV_G11
XG4479 XI11_5/XI0/XI0_62/d__0_ XI11_5/XI0/XI0_62/d_0_ DECAP_INV_G11
XG4480 XI11_5/XI0/XI0_62/d_15_ XI11_5/XI0/XI0_62/d__15_ DECAP_INV_G11
XG4481 XI11_5/XI0/XI0_62/d_14_ XI11_5/XI0/XI0_62/d__14_ DECAP_INV_G11
XG4482 XI11_5/XI0/XI0_62/d_13_ XI11_5/XI0/XI0_62/d__13_ DECAP_INV_G11
XG4483 XI11_5/XI0/XI0_62/d_12_ XI11_5/XI0/XI0_62/d__12_ DECAP_INV_G11
XG4484 XI11_5/XI0/XI0_62/d_11_ XI11_5/XI0/XI0_62/d__11_ DECAP_INV_G11
XG4485 XI11_5/XI0/XI0_62/d_10_ XI11_5/XI0/XI0_62/d__10_ DECAP_INV_G11
XG4486 XI11_5/XI0/XI0_62/d_9_ XI11_5/XI0/XI0_62/d__9_ DECAP_INV_G11
XG4487 XI11_5/XI0/XI0_62/d_8_ XI11_5/XI0/XI0_62/d__8_ DECAP_INV_G11
XG4488 XI11_5/XI0/XI0_62/d_7_ XI11_5/XI0/XI0_62/d__7_ DECAP_INV_G11
XG4489 XI11_5/XI0/XI0_62/d_6_ XI11_5/XI0/XI0_62/d__6_ DECAP_INV_G11
XG4490 XI11_5/XI0/XI0_62/d_5_ XI11_5/XI0/XI0_62/d__5_ DECAP_INV_G11
XG4491 XI11_5/XI0/XI0_62/d_4_ XI11_5/XI0/XI0_62/d__4_ DECAP_INV_G11
XG4492 XI11_5/XI0/XI0_62/d_3_ XI11_5/XI0/XI0_62/d__3_ DECAP_INV_G11
XG4493 XI11_5/XI0/XI0_62/d_2_ XI11_5/XI0/XI0_62/d__2_ DECAP_INV_G11
XG4494 XI11_5/XI0/XI0_62/d_1_ XI11_5/XI0/XI0_62/d__1_ DECAP_INV_G11
XG4495 XI11_5/XI0/XI0_62/d_0_ XI11_5/XI0/XI0_62/d__0_ DECAP_INV_G11
XG4496 XI11_5/XI0/XI0_61/d__15_ XI11_5/XI0/XI0_61/d_15_ DECAP_INV_G11
XG4497 XI11_5/XI0/XI0_61/d__14_ XI11_5/XI0/XI0_61/d_14_ DECAP_INV_G11
XG4498 XI11_5/XI0/XI0_61/d__13_ XI11_5/XI0/XI0_61/d_13_ DECAP_INV_G11
XG4499 XI11_5/XI0/XI0_61/d__12_ XI11_5/XI0/XI0_61/d_12_ DECAP_INV_G11
XG4500 XI11_5/XI0/XI0_61/d__11_ XI11_5/XI0/XI0_61/d_11_ DECAP_INV_G11
XG4501 XI11_5/XI0/XI0_61/d__10_ XI11_5/XI0/XI0_61/d_10_ DECAP_INV_G11
XG4502 XI11_5/XI0/XI0_61/d__9_ XI11_5/XI0/XI0_61/d_9_ DECAP_INV_G11
XG4503 XI11_5/XI0/XI0_61/d__8_ XI11_5/XI0/XI0_61/d_8_ DECAP_INV_G11
XG4504 XI11_5/XI0/XI0_61/d__7_ XI11_5/XI0/XI0_61/d_7_ DECAP_INV_G11
XG4505 XI11_5/XI0/XI0_61/d__6_ XI11_5/XI0/XI0_61/d_6_ DECAP_INV_G11
XG4506 XI11_5/XI0/XI0_61/d__5_ XI11_5/XI0/XI0_61/d_5_ DECAP_INV_G11
XG4507 XI11_5/XI0/XI0_61/d__4_ XI11_5/XI0/XI0_61/d_4_ DECAP_INV_G11
XG4508 XI11_5/XI0/XI0_61/d__3_ XI11_5/XI0/XI0_61/d_3_ DECAP_INV_G11
XG4509 XI11_5/XI0/XI0_61/d__2_ XI11_5/XI0/XI0_61/d_2_ DECAP_INV_G11
XG4510 XI11_5/XI0/XI0_61/d__1_ XI11_5/XI0/XI0_61/d_1_ DECAP_INV_G11
XG4511 XI11_5/XI0/XI0_61/d__0_ XI11_5/XI0/XI0_61/d_0_ DECAP_INV_G11
XG4512 XI11_5/XI0/XI0_61/d_15_ XI11_5/XI0/XI0_61/d__15_ DECAP_INV_G11
XG4513 XI11_5/XI0/XI0_61/d_14_ XI11_5/XI0/XI0_61/d__14_ DECAP_INV_G11
XG4514 XI11_5/XI0/XI0_61/d_13_ XI11_5/XI0/XI0_61/d__13_ DECAP_INV_G11
XG4515 XI11_5/XI0/XI0_61/d_12_ XI11_5/XI0/XI0_61/d__12_ DECAP_INV_G11
XG4516 XI11_5/XI0/XI0_61/d_11_ XI11_5/XI0/XI0_61/d__11_ DECAP_INV_G11
XG4517 XI11_5/XI0/XI0_61/d_10_ XI11_5/XI0/XI0_61/d__10_ DECAP_INV_G11
XG4518 XI11_5/XI0/XI0_61/d_9_ XI11_5/XI0/XI0_61/d__9_ DECAP_INV_G11
XG4519 XI11_5/XI0/XI0_61/d_8_ XI11_5/XI0/XI0_61/d__8_ DECAP_INV_G11
XG4520 XI11_5/XI0/XI0_61/d_7_ XI11_5/XI0/XI0_61/d__7_ DECAP_INV_G11
XG4521 XI11_5/XI0/XI0_61/d_6_ XI11_5/XI0/XI0_61/d__6_ DECAP_INV_G11
XG4522 XI11_5/XI0/XI0_61/d_5_ XI11_5/XI0/XI0_61/d__5_ DECAP_INV_G11
XG4523 XI11_5/XI0/XI0_61/d_4_ XI11_5/XI0/XI0_61/d__4_ DECAP_INV_G11
XG4524 XI11_5/XI0/XI0_61/d_3_ XI11_5/XI0/XI0_61/d__3_ DECAP_INV_G11
XG4525 XI11_5/XI0/XI0_61/d_2_ XI11_5/XI0/XI0_61/d__2_ DECAP_INV_G11
XG4526 XI11_5/XI0/XI0_61/d_1_ XI11_5/XI0/XI0_61/d__1_ DECAP_INV_G11
XG4527 XI11_5/XI0/XI0_61/d_0_ XI11_5/XI0/XI0_61/d__0_ DECAP_INV_G11
XG4528 XI11_5/XI0/XI0_60/d__15_ XI11_5/XI0/XI0_60/d_15_ DECAP_INV_G11
XG4529 XI11_5/XI0/XI0_60/d__14_ XI11_5/XI0/XI0_60/d_14_ DECAP_INV_G11
XG4530 XI11_5/XI0/XI0_60/d__13_ XI11_5/XI0/XI0_60/d_13_ DECAP_INV_G11
XG4531 XI11_5/XI0/XI0_60/d__12_ XI11_5/XI0/XI0_60/d_12_ DECAP_INV_G11
XG4532 XI11_5/XI0/XI0_60/d__11_ XI11_5/XI0/XI0_60/d_11_ DECAP_INV_G11
XG4533 XI11_5/XI0/XI0_60/d__10_ XI11_5/XI0/XI0_60/d_10_ DECAP_INV_G11
XG4534 XI11_5/XI0/XI0_60/d__9_ XI11_5/XI0/XI0_60/d_9_ DECAP_INV_G11
XG4535 XI11_5/XI0/XI0_60/d__8_ XI11_5/XI0/XI0_60/d_8_ DECAP_INV_G11
XG4536 XI11_5/XI0/XI0_60/d__7_ XI11_5/XI0/XI0_60/d_7_ DECAP_INV_G11
XG4537 XI11_5/XI0/XI0_60/d__6_ XI11_5/XI0/XI0_60/d_6_ DECAP_INV_G11
XG4538 XI11_5/XI0/XI0_60/d__5_ XI11_5/XI0/XI0_60/d_5_ DECAP_INV_G11
XG4539 XI11_5/XI0/XI0_60/d__4_ XI11_5/XI0/XI0_60/d_4_ DECAP_INV_G11
XG4540 XI11_5/XI0/XI0_60/d__3_ XI11_5/XI0/XI0_60/d_3_ DECAP_INV_G11
XG4541 XI11_5/XI0/XI0_60/d__2_ XI11_5/XI0/XI0_60/d_2_ DECAP_INV_G11
XG4542 XI11_5/XI0/XI0_60/d__1_ XI11_5/XI0/XI0_60/d_1_ DECAP_INV_G11
XG4543 XI11_5/XI0/XI0_60/d__0_ XI11_5/XI0/XI0_60/d_0_ DECAP_INV_G11
XG4544 XI11_5/XI0/XI0_60/d_15_ XI11_5/XI0/XI0_60/d__15_ DECAP_INV_G11
XG4545 XI11_5/XI0/XI0_60/d_14_ XI11_5/XI0/XI0_60/d__14_ DECAP_INV_G11
XG4546 XI11_5/XI0/XI0_60/d_13_ XI11_5/XI0/XI0_60/d__13_ DECAP_INV_G11
XG4547 XI11_5/XI0/XI0_60/d_12_ XI11_5/XI0/XI0_60/d__12_ DECAP_INV_G11
XG4548 XI11_5/XI0/XI0_60/d_11_ XI11_5/XI0/XI0_60/d__11_ DECAP_INV_G11
XG4549 XI11_5/XI0/XI0_60/d_10_ XI11_5/XI0/XI0_60/d__10_ DECAP_INV_G11
XG4550 XI11_5/XI0/XI0_60/d_9_ XI11_5/XI0/XI0_60/d__9_ DECAP_INV_G11
XG4551 XI11_5/XI0/XI0_60/d_8_ XI11_5/XI0/XI0_60/d__8_ DECAP_INV_G11
XG4552 XI11_5/XI0/XI0_60/d_7_ XI11_5/XI0/XI0_60/d__7_ DECAP_INV_G11
XG4553 XI11_5/XI0/XI0_60/d_6_ XI11_5/XI0/XI0_60/d__6_ DECAP_INV_G11
XG4554 XI11_5/XI0/XI0_60/d_5_ XI11_5/XI0/XI0_60/d__5_ DECAP_INV_G11
XG4555 XI11_5/XI0/XI0_60/d_4_ XI11_5/XI0/XI0_60/d__4_ DECAP_INV_G11
XG4556 XI11_5/XI0/XI0_60/d_3_ XI11_5/XI0/XI0_60/d__3_ DECAP_INV_G11
XG4557 XI11_5/XI0/XI0_60/d_2_ XI11_5/XI0/XI0_60/d__2_ DECAP_INV_G11
XG4558 XI11_5/XI0/XI0_60/d_1_ XI11_5/XI0/XI0_60/d__1_ DECAP_INV_G11
XG4559 XI11_5/XI0/XI0_60/d_0_ XI11_5/XI0/XI0_60/d__0_ DECAP_INV_G11
XG4560 XI11_5/XI0/XI0_59/d__15_ XI11_5/XI0/XI0_59/d_15_ DECAP_INV_G11
XG4561 XI11_5/XI0/XI0_59/d__14_ XI11_5/XI0/XI0_59/d_14_ DECAP_INV_G11
XG4562 XI11_5/XI0/XI0_59/d__13_ XI11_5/XI0/XI0_59/d_13_ DECAP_INV_G11
XG4563 XI11_5/XI0/XI0_59/d__12_ XI11_5/XI0/XI0_59/d_12_ DECAP_INV_G11
XG4564 XI11_5/XI0/XI0_59/d__11_ XI11_5/XI0/XI0_59/d_11_ DECAP_INV_G11
XG4565 XI11_5/XI0/XI0_59/d__10_ XI11_5/XI0/XI0_59/d_10_ DECAP_INV_G11
XG4566 XI11_5/XI0/XI0_59/d__9_ XI11_5/XI0/XI0_59/d_9_ DECAP_INV_G11
XG4567 XI11_5/XI0/XI0_59/d__8_ XI11_5/XI0/XI0_59/d_8_ DECAP_INV_G11
XG4568 XI11_5/XI0/XI0_59/d__7_ XI11_5/XI0/XI0_59/d_7_ DECAP_INV_G11
XG4569 XI11_5/XI0/XI0_59/d__6_ XI11_5/XI0/XI0_59/d_6_ DECAP_INV_G11
XG4570 XI11_5/XI0/XI0_59/d__5_ XI11_5/XI0/XI0_59/d_5_ DECAP_INV_G11
XG4571 XI11_5/XI0/XI0_59/d__4_ XI11_5/XI0/XI0_59/d_4_ DECAP_INV_G11
XG4572 XI11_5/XI0/XI0_59/d__3_ XI11_5/XI0/XI0_59/d_3_ DECAP_INV_G11
XG4573 XI11_5/XI0/XI0_59/d__2_ XI11_5/XI0/XI0_59/d_2_ DECAP_INV_G11
XG4574 XI11_5/XI0/XI0_59/d__1_ XI11_5/XI0/XI0_59/d_1_ DECAP_INV_G11
XG4575 XI11_5/XI0/XI0_59/d__0_ XI11_5/XI0/XI0_59/d_0_ DECAP_INV_G11
XG4576 XI11_5/XI0/XI0_59/d_15_ XI11_5/XI0/XI0_59/d__15_ DECAP_INV_G11
XG4577 XI11_5/XI0/XI0_59/d_14_ XI11_5/XI0/XI0_59/d__14_ DECAP_INV_G11
XG4578 XI11_5/XI0/XI0_59/d_13_ XI11_5/XI0/XI0_59/d__13_ DECAP_INV_G11
XG4579 XI11_5/XI0/XI0_59/d_12_ XI11_5/XI0/XI0_59/d__12_ DECAP_INV_G11
XG4580 XI11_5/XI0/XI0_59/d_11_ XI11_5/XI0/XI0_59/d__11_ DECAP_INV_G11
XG4581 XI11_5/XI0/XI0_59/d_10_ XI11_5/XI0/XI0_59/d__10_ DECAP_INV_G11
XG4582 XI11_5/XI0/XI0_59/d_9_ XI11_5/XI0/XI0_59/d__9_ DECAP_INV_G11
XG4583 XI11_5/XI0/XI0_59/d_8_ XI11_5/XI0/XI0_59/d__8_ DECAP_INV_G11
XG4584 XI11_5/XI0/XI0_59/d_7_ XI11_5/XI0/XI0_59/d__7_ DECAP_INV_G11
XG4585 XI11_5/XI0/XI0_59/d_6_ XI11_5/XI0/XI0_59/d__6_ DECAP_INV_G11
XG4586 XI11_5/XI0/XI0_59/d_5_ XI11_5/XI0/XI0_59/d__5_ DECAP_INV_G11
XG4587 XI11_5/XI0/XI0_59/d_4_ XI11_5/XI0/XI0_59/d__4_ DECAP_INV_G11
XG4588 XI11_5/XI0/XI0_59/d_3_ XI11_5/XI0/XI0_59/d__3_ DECAP_INV_G11
XG4589 XI11_5/XI0/XI0_59/d_2_ XI11_5/XI0/XI0_59/d__2_ DECAP_INV_G11
XG4590 XI11_5/XI0/XI0_59/d_1_ XI11_5/XI0/XI0_59/d__1_ DECAP_INV_G11
XG4591 XI11_5/XI0/XI0_59/d_0_ XI11_5/XI0/XI0_59/d__0_ DECAP_INV_G11
XG4592 XI11_5/XI0/XI0_58/d__15_ XI11_5/XI0/XI0_58/d_15_ DECAP_INV_G11
XG4593 XI11_5/XI0/XI0_58/d__14_ XI11_5/XI0/XI0_58/d_14_ DECAP_INV_G11
XG4594 XI11_5/XI0/XI0_58/d__13_ XI11_5/XI0/XI0_58/d_13_ DECAP_INV_G11
XG4595 XI11_5/XI0/XI0_58/d__12_ XI11_5/XI0/XI0_58/d_12_ DECAP_INV_G11
XG4596 XI11_5/XI0/XI0_58/d__11_ XI11_5/XI0/XI0_58/d_11_ DECAP_INV_G11
XG4597 XI11_5/XI0/XI0_58/d__10_ XI11_5/XI0/XI0_58/d_10_ DECAP_INV_G11
XG4598 XI11_5/XI0/XI0_58/d__9_ XI11_5/XI0/XI0_58/d_9_ DECAP_INV_G11
XG4599 XI11_5/XI0/XI0_58/d__8_ XI11_5/XI0/XI0_58/d_8_ DECAP_INV_G11
XG4600 XI11_5/XI0/XI0_58/d__7_ XI11_5/XI0/XI0_58/d_7_ DECAP_INV_G11
XG4601 XI11_5/XI0/XI0_58/d__6_ XI11_5/XI0/XI0_58/d_6_ DECAP_INV_G11
XG4602 XI11_5/XI0/XI0_58/d__5_ XI11_5/XI0/XI0_58/d_5_ DECAP_INV_G11
XG4603 XI11_5/XI0/XI0_58/d__4_ XI11_5/XI0/XI0_58/d_4_ DECAP_INV_G11
XG4604 XI11_5/XI0/XI0_58/d__3_ XI11_5/XI0/XI0_58/d_3_ DECAP_INV_G11
XG4605 XI11_5/XI0/XI0_58/d__2_ XI11_5/XI0/XI0_58/d_2_ DECAP_INV_G11
XG4606 XI11_5/XI0/XI0_58/d__1_ XI11_5/XI0/XI0_58/d_1_ DECAP_INV_G11
XG4607 XI11_5/XI0/XI0_58/d__0_ XI11_5/XI0/XI0_58/d_0_ DECAP_INV_G11
XG4608 XI11_5/XI0/XI0_58/d_15_ XI11_5/XI0/XI0_58/d__15_ DECAP_INV_G11
XG4609 XI11_5/XI0/XI0_58/d_14_ XI11_5/XI0/XI0_58/d__14_ DECAP_INV_G11
XG4610 XI11_5/XI0/XI0_58/d_13_ XI11_5/XI0/XI0_58/d__13_ DECAP_INV_G11
XG4611 XI11_5/XI0/XI0_58/d_12_ XI11_5/XI0/XI0_58/d__12_ DECAP_INV_G11
XG4612 XI11_5/XI0/XI0_58/d_11_ XI11_5/XI0/XI0_58/d__11_ DECAP_INV_G11
XG4613 XI11_5/XI0/XI0_58/d_10_ XI11_5/XI0/XI0_58/d__10_ DECAP_INV_G11
XG4614 XI11_5/XI0/XI0_58/d_9_ XI11_5/XI0/XI0_58/d__9_ DECAP_INV_G11
XG4615 XI11_5/XI0/XI0_58/d_8_ XI11_5/XI0/XI0_58/d__8_ DECAP_INV_G11
XG4616 XI11_5/XI0/XI0_58/d_7_ XI11_5/XI0/XI0_58/d__7_ DECAP_INV_G11
XG4617 XI11_5/XI0/XI0_58/d_6_ XI11_5/XI0/XI0_58/d__6_ DECAP_INV_G11
XG4618 XI11_5/XI0/XI0_58/d_5_ XI11_5/XI0/XI0_58/d__5_ DECAP_INV_G11
XG4619 XI11_5/XI0/XI0_58/d_4_ XI11_5/XI0/XI0_58/d__4_ DECAP_INV_G11
XG4620 XI11_5/XI0/XI0_58/d_3_ XI11_5/XI0/XI0_58/d__3_ DECAP_INV_G11
XG4621 XI11_5/XI0/XI0_58/d_2_ XI11_5/XI0/XI0_58/d__2_ DECAP_INV_G11
XG4622 XI11_5/XI0/XI0_58/d_1_ XI11_5/XI0/XI0_58/d__1_ DECAP_INV_G11
XG4623 XI11_5/XI0/XI0_58/d_0_ XI11_5/XI0/XI0_58/d__0_ DECAP_INV_G11
XG4624 XI11_5/XI0/XI0_57/d__15_ XI11_5/XI0/XI0_57/d_15_ DECAP_INV_G11
XG4625 XI11_5/XI0/XI0_57/d__14_ XI11_5/XI0/XI0_57/d_14_ DECAP_INV_G11
XG4626 XI11_5/XI0/XI0_57/d__13_ XI11_5/XI0/XI0_57/d_13_ DECAP_INV_G11
XG4627 XI11_5/XI0/XI0_57/d__12_ XI11_5/XI0/XI0_57/d_12_ DECAP_INV_G11
XG4628 XI11_5/XI0/XI0_57/d__11_ XI11_5/XI0/XI0_57/d_11_ DECAP_INV_G11
XG4629 XI11_5/XI0/XI0_57/d__10_ XI11_5/XI0/XI0_57/d_10_ DECAP_INV_G11
XG4630 XI11_5/XI0/XI0_57/d__9_ XI11_5/XI0/XI0_57/d_9_ DECAP_INV_G11
XG4631 XI11_5/XI0/XI0_57/d__8_ XI11_5/XI0/XI0_57/d_8_ DECAP_INV_G11
XG4632 XI11_5/XI0/XI0_57/d__7_ XI11_5/XI0/XI0_57/d_7_ DECAP_INV_G11
XG4633 XI11_5/XI0/XI0_57/d__6_ XI11_5/XI0/XI0_57/d_6_ DECAP_INV_G11
XG4634 XI11_5/XI0/XI0_57/d__5_ XI11_5/XI0/XI0_57/d_5_ DECAP_INV_G11
XG4635 XI11_5/XI0/XI0_57/d__4_ XI11_5/XI0/XI0_57/d_4_ DECAP_INV_G11
XG4636 XI11_5/XI0/XI0_57/d__3_ XI11_5/XI0/XI0_57/d_3_ DECAP_INV_G11
XG4637 XI11_5/XI0/XI0_57/d__2_ XI11_5/XI0/XI0_57/d_2_ DECAP_INV_G11
XG4638 XI11_5/XI0/XI0_57/d__1_ XI11_5/XI0/XI0_57/d_1_ DECAP_INV_G11
XG4639 XI11_5/XI0/XI0_57/d__0_ XI11_5/XI0/XI0_57/d_0_ DECAP_INV_G11
XG4640 XI11_5/XI0/XI0_57/d_15_ XI11_5/XI0/XI0_57/d__15_ DECAP_INV_G11
XG4641 XI11_5/XI0/XI0_57/d_14_ XI11_5/XI0/XI0_57/d__14_ DECAP_INV_G11
XG4642 XI11_5/XI0/XI0_57/d_13_ XI11_5/XI0/XI0_57/d__13_ DECAP_INV_G11
XG4643 XI11_5/XI0/XI0_57/d_12_ XI11_5/XI0/XI0_57/d__12_ DECAP_INV_G11
XG4644 XI11_5/XI0/XI0_57/d_11_ XI11_5/XI0/XI0_57/d__11_ DECAP_INV_G11
XG4645 XI11_5/XI0/XI0_57/d_10_ XI11_5/XI0/XI0_57/d__10_ DECAP_INV_G11
XG4646 XI11_5/XI0/XI0_57/d_9_ XI11_5/XI0/XI0_57/d__9_ DECAP_INV_G11
XG4647 XI11_5/XI0/XI0_57/d_8_ XI11_5/XI0/XI0_57/d__8_ DECAP_INV_G11
XG4648 XI11_5/XI0/XI0_57/d_7_ XI11_5/XI0/XI0_57/d__7_ DECAP_INV_G11
XG4649 XI11_5/XI0/XI0_57/d_6_ XI11_5/XI0/XI0_57/d__6_ DECAP_INV_G11
XG4650 XI11_5/XI0/XI0_57/d_5_ XI11_5/XI0/XI0_57/d__5_ DECAP_INV_G11
XG4651 XI11_5/XI0/XI0_57/d_4_ XI11_5/XI0/XI0_57/d__4_ DECAP_INV_G11
XG4652 XI11_5/XI0/XI0_57/d_3_ XI11_5/XI0/XI0_57/d__3_ DECAP_INV_G11
XG4653 XI11_5/XI0/XI0_57/d_2_ XI11_5/XI0/XI0_57/d__2_ DECAP_INV_G11
XG4654 XI11_5/XI0/XI0_57/d_1_ XI11_5/XI0/XI0_57/d__1_ DECAP_INV_G11
XG4655 XI11_5/XI0/XI0_57/d_0_ XI11_5/XI0/XI0_57/d__0_ DECAP_INV_G11
XG4656 XI11_5/XI0/XI0_56/d__15_ XI11_5/XI0/XI0_56/d_15_ DECAP_INV_G11
XG4657 XI11_5/XI0/XI0_56/d__14_ XI11_5/XI0/XI0_56/d_14_ DECAP_INV_G11
XG4658 XI11_5/XI0/XI0_56/d__13_ XI11_5/XI0/XI0_56/d_13_ DECAP_INV_G11
XG4659 XI11_5/XI0/XI0_56/d__12_ XI11_5/XI0/XI0_56/d_12_ DECAP_INV_G11
XG4660 XI11_5/XI0/XI0_56/d__11_ XI11_5/XI0/XI0_56/d_11_ DECAP_INV_G11
XG4661 XI11_5/XI0/XI0_56/d__10_ XI11_5/XI0/XI0_56/d_10_ DECAP_INV_G11
XG4662 XI11_5/XI0/XI0_56/d__9_ XI11_5/XI0/XI0_56/d_9_ DECAP_INV_G11
XG4663 XI11_5/XI0/XI0_56/d__8_ XI11_5/XI0/XI0_56/d_8_ DECAP_INV_G11
XG4664 XI11_5/XI0/XI0_56/d__7_ XI11_5/XI0/XI0_56/d_7_ DECAP_INV_G11
XG4665 XI11_5/XI0/XI0_56/d__6_ XI11_5/XI0/XI0_56/d_6_ DECAP_INV_G11
XG4666 XI11_5/XI0/XI0_56/d__5_ XI11_5/XI0/XI0_56/d_5_ DECAP_INV_G11
XG4667 XI11_5/XI0/XI0_56/d__4_ XI11_5/XI0/XI0_56/d_4_ DECAP_INV_G11
XG4668 XI11_5/XI0/XI0_56/d__3_ XI11_5/XI0/XI0_56/d_3_ DECAP_INV_G11
XG4669 XI11_5/XI0/XI0_56/d__2_ XI11_5/XI0/XI0_56/d_2_ DECAP_INV_G11
XG4670 XI11_5/XI0/XI0_56/d__1_ XI11_5/XI0/XI0_56/d_1_ DECAP_INV_G11
XG4671 XI11_5/XI0/XI0_56/d__0_ XI11_5/XI0/XI0_56/d_0_ DECAP_INV_G11
XG4672 XI11_5/XI0/XI0_56/d_15_ XI11_5/XI0/XI0_56/d__15_ DECAP_INV_G11
XG4673 XI11_5/XI0/XI0_56/d_14_ XI11_5/XI0/XI0_56/d__14_ DECAP_INV_G11
XG4674 XI11_5/XI0/XI0_56/d_13_ XI11_5/XI0/XI0_56/d__13_ DECAP_INV_G11
XG4675 XI11_5/XI0/XI0_56/d_12_ XI11_5/XI0/XI0_56/d__12_ DECAP_INV_G11
XG4676 XI11_5/XI0/XI0_56/d_11_ XI11_5/XI0/XI0_56/d__11_ DECAP_INV_G11
XG4677 XI11_5/XI0/XI0_56/d_10_ XI11_5/XI0/XI0_56/d__10_ DECAP_INV_G11
XG4678 XI11_5/XI0/XI0_56/d_9_ XI11_5/XI0/XI0_56/d__9_ DECAP_INV_G11
XG4679 XI11_5/XI0/XI0_56/d_8_ XI11_5/XI0/XI0_56/d__8_ DECAP_INV_G11
XG4680 XI11_5/XI0/XI0_56/d_7_ XI11_5/XI0/XI0_56/d__7_ DECAP_INV_G11
XG4681 XI11_5/XI0/XI0_56/d_6_ XI11_5/XI0/XI0_56/d__6_ DECAP_INV_G11
XG4682 XI11_5/XI0/XI0_56/d_5_ XI11_5/XI0/XI0_56/d__5_ DECAP_INV_G11
XG4683 XI11_5/XI0/XI0_56/d_4_ XI11_5/XI0/XI0_56/d__4_ DECAP_INV_G11
XG4684 XI11_5/XI0/XI0_56/d_3_ XI11_5/XI0/XI0_56/d__3_ DECAP_INV_G11
XG4685 XI11_5/XI0/XI0_56/d_2_ XI11_5/XI0/XI0_56/d__2_ DECAP_INV_G11
XG4686 XI11_5/XI0/XI0_56/d_1_ XI11_5/XI0/XI0_56/d__1_ DECAP_INV_G11
XG4687 XI11_5/XI0/XI0_56/d_0_ XI11_5/XI0/XI0_56/d__0_ DECAP_INV_G11
XG4688 XI11_5/XI0/XI0_55/d__15_ XI11_5/XI0/XI0_55/d_15_ DECAP_INV_G11
XG4689 XI11_5/XI0/XI0_55/d__14_ XI11_5/XI0/XI0_55/d_14_ DECAP_INV_G11
XG4690 XI11_5/XI0/XI0_55/d__13_ XI11_5/XI0/XI0_55/d_13_ DECAP_INV_G11
XG4691 XI11_5/XI0/XI0_55/d__12_ XI11_5/XI0/XI0_55/d_12_ DECAP_INV_G11
XG4692 XI11_5/XI0/XI0_55/d__11_ XI11_5/XI0/XI0_55/d_11_ DECAP_INV_G11
XG4693 XI11_5/XI0/XI0_55/d__10_ XI11_5/XI0/XI0_55/d_10_ DECAP_INV_G11
XG4694 XI11_5/XI0/XI0_55/d__9_ XI11_5/XI0/XI0_55/d_9_ DECAP_INV_G11
XG4695 XI11_5/XI0/XI0_55/d__8_ XI11_5/XI0/XI0_55/d_8_ DECAP_INV_G11
XG4696 XI11_5/XI0/XI0_55/d__7_ XI11_5/XI0/XI0_55/d_7_ DECAP_INV_G11
XG4697 XI11_5/XI0/XI0_55/d__6_ XI11_5/XI0/XI0_55/d_6_ DECAP_INV_G11
XG4698 XI11_5/XI0/XI0_55/d__5_ XI11_5/XI0/XI0_55/d_5_ DECAP_INV_G11
XG4699 XI11_5/XI0/XI0_55/d__4_ XI11_5/XI0/XI0_55/d_4_ DECAP_INV_G11
XG4700 XI11_5/XI0/XI0_55/d__3_ XI11_5/XI0/XI0_55/d_3_ DECAP_INV_G11
XG4701 XI11_5/XI0/XI0_55/d__2_ XI11_5/XI0/XI0_55/d_2_ DECAP_INV_G11
XG4702 XI11_5/XI0/XI0_55/d__1_ XI11_5/XI0/XI0_55/d_1_ DECAP_INV_G11
XG4703 XI11_5/XI0/XI0_55/d__0_ XI11_5/XI0/XI0_55/d_0_ DECAP_INV_G11
XG4704 XI11_5/XI0/XI0_55/d_15_ XI11_5/XI0/XI0_55/d__15_ DECAP_INV_G11
XG4705 XI11_5/XI0/XI0_55/d_14_ XI11_5/XI0/XI0_55/d__14_ DECAP_INV_G11
XG4706 XI11_5/XI0/XI0_55/d_13_ XI11_5/XI0/XI0_55/d__13_ DECAP_INV_G11
XG4707 XI11_5/XI0/XI0_55/d_12_ XI11_5/XI0/XI0_55/d__12_ DECAP_INV_G11
XG4708 XI11_5/XI0/XI0_55/d_11_ XI11_5/XI0/XI0_55/d__11_ DECAP_INV_G11
XG4709 XI11_5/XI0/XI0_55/d_10_ XI11_5/XI0/XI0_55/d__10_ DECAP_INV_G11
XG4710 XI11_5/XI0/XI0_55/d_9_ XI11_5/XI0/XI0_55/d__9_ DECAP_INV_G11
XG4711 XI11_5/XI0/XI0_55/d_8_ XI11_5/XI0/XI0_55/d__8_ DECAP_INV_G11
XG4712 XI11_5/XI0/XI0_55/d_7_ XI11_5/XI0/XI0_55/d__7_ DECAP_INV_G11
XG4713 XI11_5/XI0/XI0_55/d_6_ XI11_5/XI0/XI0_55/d__6_ DECAP_INV_G11
XG4714 XI11_5/XI0/XI0_55/d_5_ XI11_5/XI0/XI0_55/d__5_ DECAP_INV_G11
XG4715 XI11_5/XI0/XI0_55/d_4_ XI11_5/XI0/XI0_55/d__4_ DECAP_INV_G11
XG4716 XI11_5/XI0/XI0_55/d_3_ XI11_5/XI0/XI0_55/d__3_ DECAP_INV_G11
XG4717 XI11_5/XI0/XI0_55/d_2_ XI11_5/XI0/XI0_55/d__2_ DECAP_INV_G11
XG4718 XI11_5/XI0/XI0_55/d_1_ XI11_5/XI0/XI0_55/d__1_ DECAP_INV_G11
XG4719 XI11_5/XI0/XI0_55/d_0_ XI11_5/XI0/XI0_55/d__0_ DECAP_INV_G11
XG4720 XI11_5/XI0/XI0_54/d__15_ XI11_5/XI0/XI0_54/d_15_ DECAP_INV_G11
XG4721 XI11_5/XI0/XI0_54/d__14_ XI11_5/XI0/XI0_54/d_14_ DECAP_INV_G11
XG4722 XI11_5/XI0/XI0_54/d__13_ XI11_5/XI0/XI0_54/d_13_ DECAP_INV_G11
XG4723 XI11_5/XI0/XI0_54/d__12_ XI11_5/XI0/XI0_54/d_12_ DECAP_INV_G11
XG4724 XI11_5/XI0/XI0_54/d__11_ XI11_5/XI0/XI0_54/d_11_ DECAP_INV_G11
XG4725 XI11_5/XI0/XI0_54/d__10_ XI11_5/XI0/XI0_54/d_10_ DECAP_INV_G11
XG4726 XI11_5/XI0/XI0_54/d__9_ XI11_5/XI0/XI0_54/d_9_ DECAP_INV_G11
XG4727 XI11_5/XI0/XI0_54/d__8_ XI11_5/XI0/XI0_54/d_8_ DECAP_INV_G11
XG4728 XI11_5/XI0/XI0_54/d__7_ XI11_5/XI0/XI0_54/d_7_ DECAP_INV_G11
XG4729 XI11_5/XI0/XI0_54/d__6_ XI11_5/XI0/XI0_54/d_6_ DECAP_INV_G11
XG4730 XI11_5/XI0/XI0_54/d__5_ XI11_5/XI0/XI0_54/d_5_ DECAP_INV_G11
XG4731 XI11_5/XI0/XI0_54/d__4_ XI11_5/XI0/XI0_54/d_4_ DECAP_INV_G11
XG4732 XI11_5/XI0/XI0_54/d__3_ XI11_5/XI0/XI0_54/d_3_ DECAP_INV_G11
XG4733 XI11_5/XI0/XI0_54/d__2_ XI11_5/XI0/XI0_54/d_2_ DECAP_INV_G11
XG4734 XI11_5/XI0/XI0_54/d__1_ XI11_5/XI0/XI0_54/d_1_ DECAP_INV_G11
XG4735 XI11_5/XI0/XI0_54/d__0_ XI11_5/XI0/XI0_54/d_0_ DECAP_INV_G11
XG4736 XI11_5/XI0/XI0_54/d_15_ XI11_5/XI0/XI0_54/d__15_ DECAP_INV_G11
XG4737 XI11_5/XI0/XI0_54/d_14_ XI11_5/XI0/XI0_54/d__14_ DECAP_INV_G11
XG4738 XI11_5/XI0/XI0_54/d_13_ XI11_5/XI0/XI0_54/d__13_ DECAP_INV_G11
XG4739 XI11_5/XI0/XI0_54/d_12_ XI11_5/XI0/XI0_54/d__12_ DECAP_INV_G11
XG4740 XI11_5/XI0/XI0_54/d_11_ XI11_5/XI0/XI0_54/d__11_ DECAP_INV_G11
XG4741 XI11_5/XI0/XI0_54/d_10_ XI11_5/XI0/XI0_54/d__10_ DECAP_INV_G11
XG4742 XI11_5/XI0/XI0_54/d_9_ XI11_5/XI0/XI0_54/d__9_ DECAP_INV_G11
XG4743 XI11_5/XI0/XI0_54/d_8_ XI11_5/XI0/XI0_54/d__8_ DECAP_INV_G11
XG4744 XI11_5/XI0/XI0_54/d_7_ XI11_5/XI0/XI0_54/d__7_ DECAP_INV_G11
XG4745 XI11_5/XI0/XI0_54/d_6_ XI11_5/XI0/XI0_54/d__6_ DECAP_INV_G11
XG4746 XI11_5/XI0/XI0_54/d_5_ XI11_5/XI0/XI0_54/d__5_ DECAP_INV_G11
XG4747 XI11_5/XI0/XI0_54/d_4_ XI11_5/XI0/XI0_54/d__4_ DECAP_INV_G11
XG4748 XI11_5/XI0/XI0_54/d_3_ XI11_5/XI0/XI0_54/d__3_ DECAP_INV_G11
XG4749 XI11_5/XI0/XI0_54/d_2_ XI11_5/XI0/XI0_54/d__2_ DECAP_INV_G11
XG4750 XI11_5/XI0/XI0_54/d_1_ XI11_5/XI0/XI0_54/d__1_ DECAP_INV_G11
XG4751 XI11_5/XI0/XI0_54/d_0_ XI11_5/XI0/XI0_54/d__0_ DECAP_INV_G11
XG4752 XI11_5/XI0/XI0_53/d__15_ XI11_5/XI0/XI0_53/d_15_ DECAP_INV_G11
XG4753 XI11_5/XI0/XI0_53/d__14_ XI11_5/XI0/XI0_53/d_14_ DECAP_INV_G11
XG4754 XI11_5/XI0/XI0_53/d__13_ XI11_5/XI0/XI0_53/d_13_ DECAP_INV_G11
XG4755 XI11_5/XI0/XI0_53/d__12_ XI11_5/XI0/XI0_53/d_12_ DECAP_INV_G11
XG4756 XI11_5/XI0/XI0_53/d__11_ XI11_5/XI0/XI0_53/d_11_ DECAP_INV_G11
XG4757 XI11_5/XI0/XI0_53/d__10_ XI11_5/XI0/XI0_53/d_10_ DECAP_INV_G11
XG4758 XI11_5/XI0/XI0_53/d__9_ XI11_5/XI0/XI0_53/d_9_ DECAP_INV_G11
XG4759 XI11_5/XI0/XI0_53/d__8_ XI11_5/XI0/XI0_53/d_8_ DECAP_INV_G11
XG4760 XI11_5/XI0/XI0_53/d__7_ XI11_5/XI0/XI0_53/d_7_ DECAP_INV_G11
XG4761 XI11_5/XI0/XI0_53/d__6_ XI11_5/XI0/XI0_53/d_6_ DECAP_INV_G11
XG4762 XI11_5/XI0/XI0_53/d__5_ XI11_5/XI0/XI0_53/d_5_ DECAP_INV_G11
XG4763 XI11_5/XI0/XI0_53/d__4_ XI11_5/XI0/XI0_53/d_4_ DECAP_INV_G11
XG4764 XI11_5/XI0/XI0_53/d__3_ XI11_5/XI0/XI0_53/d_3_ DECAP_INV_G11
XG4765 XI11_5/XI0/XI0_53/d__2_ XI11_5/XI0/XI0_53/d_2_ DECAP_INV_G11
XG4766 XI11_5/XI0/XI0_53/d__1_ XI11_5/XI0/XI0_53/d_1_ DECAP_INV_G11
XG4767 XI11_5/XI0/XI0_53/d__0_ XI11_5/XI0/XI0_53/d_0_ DECAP_INV_G11
XG4768 XI11_5/XI0/XI0_53/d_15_ XI11_5/XI0/XI0_53/d__15_ DECAP_INV_G11
XG4769 XI11_5/XI0/XI0_53/d_14_ XI11_5/XI0/XI0_53/d__14_ DECAP_INV_G11
XG4770 XI11_5/XI0/XI0_53/d_13_ XI11_5/XI0/XI0_53/d__13_ DECAP_INV_G11
XG4771 XI11_5/XI0/XI0_53/d_12_ XI11_5/XI0/XI0_53/d__12_ DECAP_INV_G11
XG4772 XI11_5/XI0/XI0_53/d_11_ XI11_5/XI0/XI0_53/d__11_ DECAP_INV_G11
XG4773 XI11_5/XI0/XI0_53/d_10_ XI11_5/XI0/XI0_53/d__10_ DECAP_INV_G11
XG4774 XI11_5/XI0/XI0_53/d_9_ XI11_5/XI0/XI0_53/d__9_ DECAP_INV_G11
XG4775 XI11_5/XI0/XI0_53/d_8_ XI11_5/XI0/XI0_53/d__8_ DECAP_INV_G11
XG4776 XI11_5/XI0/XI0_53/d_7_ XI11_5/XI0/XI0_53/d__7_ DECAP_INV_G11
XG4777 XI11_5/XI0/XI0_53/d_6_ XI11_5/XI0/XI0_53/d__6_ DECAP_INV_G11
XG4778 XI11_5/XI0/XI0_53/d_5_ XI11_5/XI0/XI0_53/d__5_ DECAP_INV_G11
XG4779 XI11_5/XI0/XI0_53/d_4_ XI11_5/XI0/XI0_53/d__4_ DECAP_INV_G11
XG4780 XI11_5/XI0/XI0_53/d_3_ XI11_5/XI0/XI0_53/d__3_ DECAP_INV_G11
XG4781 XI11_5/XI0/XI0_53/d_2_ XI11_5/XI0/XI0_53/d__2_ DECAP_INV_G11
XG4782 XI11_5/XI0/XI0_53/d_1_ XI11_5/XI0/XI0_53/d__1_ DECAP_INV_G11
XG4783 XI11_5/XI0/XI0_53/d_0_ XI11_5/XI0/XI0_53/d__0_ DECAP_INV_G11
XG4784 XI11_5/XI0/XI0_52/d__15_ XI11_5/XI0/XI0_52/d_15_ DECAP_INV_G11
XG4785 XI11_5/XI0/XI0_52/d__14_ XI11_5/XI0/XI0_52/d_14_ DECAP_INV_G11
XG4786 XI11_5/XI0/XI0_52/d__13_ XI11_5/XI0/XI0_52/d_13_ DECAP_INV_G11
XG4787 XI11_5/XI0/XI0_52/d__12_ XI11_5/XI0/XI0_52/d_12_ DECAP_INV_G11
XG4788 XI11_5/XI0/XI0_52/d__11_ XI11_5/XI0/XI0_52/d_11_ DECAP_INV_G11
XG4789 XI11_5/XI0/XI0_52/d__10_ XI11_5/XI0/XI0_52/d_10_ DECAP_INV_G11
XG4790 XI11_5/XI0/XI0_52/d__9_ XI11_5/XI0/XI0_52/d_9_ DECAP_INV_G11
XG4791 XI11_5/XI0/XI0_52/d__8_ XI11_5/XI0/XI0_52/d_8_ DECAP_INV_G11
XG4792 XI11_5/XI0/XI0_52/d__7_ XI11_5/XI0/XI0_52/d_7_ DECAP_INV_G11
XG4793 XI11_5/XI0/XI0_52/d__6_ XI11_5/XI0/XI0_52/d_6_ DECAP_INV_G11
XG4794 XI11_5/XI0/XI0_52/d__5_ XI11_5/XI0/XI0_52/d_5_ DECAP_INV_G11
XG4795 XI11_5/XI0/XI0_52/d__4_ XI11_5/XI0/XI0_52/d_4_ DECAP_INV_G11
XG4796 XI11_5/XI0/XI0_52/d__3_ XI11_5/XI0/XI0_52/d_3_ DECAP_INV_G11
XG4797 XI11_5/XI0/XI0_52/d__2_ XI11_5/XI0/XI0_52/d_2_ DECAP_INV_G11
XG4798 XI11_5/XI0/XI0_52/d__1_ XI11_5/XI0/XI0_52/d_1_ DECAP_INV_G11
XG4799 XI11_5/XI0/XI0_52/d__0_ XI11_5/XI0/XI0_52/d_0_ DECAP_INV_G11
XG4800 XI11_5/XI0/XI0_52/d_15_ XI11_5/XI0/XI0_52/d__15_ DECAP_INV_G11
XG4801 XI11_5/XI0/XI0_52/d_14_ XI11_5/XI0/XI0_52/d__14_ DECAP_INV_G11
XG4802 XI11_5/XI0/XI0_52/d_13_ XI11_5/XI0/XI0_52/d__13_ DECAP_INV_G11
XG4803 XI11_5/XI0/XI0_52/d_12_ XI11_5/XI0/XI0_52/d__12_ DECAP_INV_G11
XG4804 XI11_5/XI0/XI0_52/d_11_ XI11_5/XI0/XI0_52/d__11_ DECAP_INV_G11
XG4805 XI11_5/XI0/XI0_52/d_10_ XI11_5/XI0/XI0_52/d__10_ DECAP_INV_G11
XG4806 XI11_5/XI0/XI0_52/d_9_ XI11_5/XI0/XI0_52/d__9_ DECAP_INV_G11
XG4807 XI11_5/XI0/XI0_52/d_8_ XI11_5/XI0/XI0_52/d__8_ DECAP_INV_G11
XG4808 XI11_5/XI0/XI0_52/d_7_ XI11_5/XI0/XI0_52/d__7_ DECAP_INV_G11
XG4809 XI11_5/XI0/XI0_52/d_6_ XI11_5/XI0/XI0_52/d__6_ DECAP_INV_G11
XG4810 XI11_5/XI0/XI0_52/d_5_ XI11_5/XI0/XI0_52/d__5_ DECAP_INV_G11
XG4811 XI11_5/XI0/XI0_52/d_4_ XI11_5/XI0/XI0_52/d__4_ DECAP_INV_G11
XG4812 XI11_5/XI0/XI0_52/d_3_ XI11_5/XI0/XI0_52/d__3_ DECAP_INV_G11
XG4813 XI11_5/XI0/XI0_52/d_2_ XI11_5/XI0/XI0_52/d__2_ DECAP_INV_G11
XG4814 XI11_5/XI0/XI0_52/d_1_ XI11_5/XI0/XI0_52/d__1_ DECAP_INV_G11
XG4815 XI11_5/XI0/XI0_52/d_0_ XI11_5/XI0/XI0_52/d__0_ DECAP_INV_G11
XG4816 XI11_5/XI0/XI0_51/d__15_ XI11_5/XI0/XI0_51/d_15_ DECAP_INV_G11
XG4817 XI11_5/XI0/XI0_51/d__14_ XI11_5/XI0/XI0_51/d_14_ DECAP_INV_G11
XG4818 XI11_5/XI0/XI0_51/d__13_ XI11_5/XI0/XI0_51/d_13_ DECAP_INV_G11
XG4819 XI11_5/XI0/XI0_51/d__12_ XI11_5/XI0/XI0_51/d_12_ DECAP_INV_G11
XG4820 XI11_5/XI0/XI0_51/d__11_ XI11_5/XI0/XI0_51/d_11_ DECAP_INV_G11
XG4821 XI11_5/XI0/XI0_51/d__10_ XI11_5/XI0/XI0_51/d_10_ DECAP_INV_G11
XG4822 XI11_5/XI0/XI0_51/d__9_ XI11_5/XI0/XI0_51/d_9_ DECAP_INV_G11
XG4823 XI11_5/XI0/XI0_51/d__8_ XI11_5/XI0/XI0_51/d_8_ DECAP_INV_G11
XG4824 XI11_5/XI0/XI0_51/d__7_ XI11_5/XI0/XI0_51/d_7_ DECAP_INV_G11
XG4825 XI11_5/XI0/XI0_51/d__6_ XI11_5/XI0/XI0_51/d_6_ DECAP_INV_G11
XG4826 XI11_5/XI0/XI0_51/d__5_ XI11_5/XI0/XI0_51/d_5_ DECAP_INV_G11
XG4827 XI11_5/XI0/XI0_51/d__4_ XI11_5/XI0/XI0_51/d_4_ DECAP_INV_G11
XG4828 XI11_5/XI0/XI0_51/d__3_ XI11_5/XI0/XI0_51/d_3_ DECAP_INV_G11
XG4829 XI11_5/XI0/XI0_51/d__2_ XI11_5/XI0/XI0_51/d_2_ DECAP_INV_G11
XG4830 XI11_5/XI0/XI0_51/d__1_ XI11_5/XI0/XI0_51/d_1_ DECAP_INV_G11
XG4831 XI11_5/XI0/XI0_51/d__0_ XI11_5/XI0/XI0_51/d_0_ DECAP_INV_G11
XG4832 XI11_5/XI0/XI0_51/d_15_ XI11_5/XI0/XI0_51/d__15_ DECAP_INV_G11
XG4833 XI11_5/XI0/XI0_51/d_14_ XI11_5/XI0/XI0_51/d__14_ DECAP_INV_G11
XG4834 XI11_5/XI0/XI0_51/d_13_ XI11_5/XI0/XI0_51/d__13_ DECAP_INV_G11
XG4835 XI11_5/XI0/XI0_51/d_12_ XI11_5/XI0/XI0_51/d__12_ DECAP_INV_G11
XG4836 XI11_5/XI0/XI0_51/d_11_ XI11_5/XI0/XI0_51/d__11_ DECAP_INV_G11
XG4837 XI11_5/XI0/XI0_51/d_10_ XI11_5/XI0/XI0_51/d__10_ DECAP_INV_G11
XG4838 XI11_5/XI0/XI0_51/d_9_ XI11_5/XI0/XI0_51/d__9_ DECAP_INV_G11
XG4839 XI11_5/XI0/XI0_51/d_8_ XI11_5/XI0/XI0_51/d__8_ DECAP_INV_G11
XG4840 XI11_5/XI0/XI0_51/d_7_ XI11_5/XI0/XI0_51/d__7_ DECAP_INV_G11
XG4841 XI11_5/XI0/XI0_51/d_6_ XI11_5/XI0/XI0_51/d__6_ DECAP_INV_G11
XG4842 XI11_5/XI0/XI0_51/d_5_ XI11_5/XI0/XI0_51/d__5_ DECAP_INV_G11
XG4843 XI11_5/XI0/XI0_51/d_4_ XI11_5/XI0/XI0_51/d__4_ DECAP_INV_G11
XG4844 XI11_5/XI0/XI0_51/d_3_ XI11_5/XI0/XI0_51/d__3_ DECAP_INV_G11
XG4845 XI11_5/XI0/XI0_51/d_2_ XI11_5/XI0/XI0_51/d__2_ DECAP_INV_G11
XG4846 XI11_5/XI0/XI0_51/d_1_ XI11_5/XI0/XI0_51/d__1_ DECAP_INV_G11
XG4847 XI11_5/XI0/XI0_51/d_0_ XI11_5/XI0/XI0_51/d__0_ DECAP_INV_G11
XG4848 XI11_5/XI0/XI0_50/d__15_ XI11_5/XI0/XI0_50/d_15_ DECAP_INV_G11
XG4849 XI11_5/XI0/XI0_50/d__14_ XI11_5/XI0/XI0_50/d_14_ DECAP_INV_G11
XG4850 XI11_5/XI0/XI0_50/d__13_ XI11_5/XI0/XI0_50/d_13_ DECAP_INV_G11
XG4851 XI11_5/XI0/XI0_50/d__12_ XI11_5/XI0/XI0_50/d_12_ DECAP_INV_G11
XG4852 XI11_5/XI0/XI0_50/d__11_ XI11_5/XI0/XI0_50/d_11_ DECAP_INV_G11
XG4853 XI11_5/XI0/XI0_50/d__10_ XI11_5/XI0/XI0_50/d_10_ DECAP_INV_G11
XG4854 XI11_5/XI0/XI0_50/d__9_ XI11_5/XI0/XI0_50/d_9_ DECAP_INV_G11
XG4855 XI11_5/XI0/XI0_50/d__8_ XI11_5/XI0/XI0_50/d_8_ DECAP_INV_G11
XG4856 XI11_5/XI0/XI0_50/d__7_ XI11_5/XI0/XI0_50/d_7_ DECAP_INV_G11
XG4857 XI11_5/XI0/XI0_50/d__6_ XI11_5/XI0/XI0_50/d_6_ DECAP_INV_G11
XG4858 XI11_5/XI0/XI0_50/d__5_ XI11_5/XI0/XI0_50/d_5_ DECAP_INV_G11
XG4859 XI11_5/XI0/XI0_50/d__4_ XI11_5/XI0/XI0_50/d_4_ DECAP_INV_G11
XG4860 XI11_5/XI0/XI0_50/d__3_ XI11_5/XI0/XI0_50/d_3_ DECAP_INV_G11
XG4861 XI11_5/XI0/XI0_50/d__2_ XI11_5/XI0/XI0_50/d_2_ DECAP_INV_G11
XG4862 XI11_5/XI0/XI0_50/d__1_ XI11_5/XI0/XI0_50/d_1_ DECAP_INV_G11
XG4863 XI11_5/XI0/XI0_50/d__0_ XI11_5/XI0/XI0_50/d_0_ DECAP_INV_G11
XG4864 XI11_5/XI0/XI0_50/d_15_ XI11_5/XI0/XI0_50/d__15_ DECAP_INV_G11
XG4865 XI11_5/XI0/XI0_50/d_14_ XI11_5/XI0/XI0_50/d__14_ DECAP_INV_G11
XG4866 XI11_5/XI0/XI0_50/d_13_ XI11_5/XI0/XI0_50/d__13_ DECAP_INV_G11
XG4867 XI11_5/XI0/XI0_50/d_12_ XI11_5/XI0/XI0_50/d__12_ DECAP_INV_G11
XG4868 XI11_5/XI0/XI0_50/d_11_ XI11_5/XI0/XI0_50/d__11_ DECAP_INV_G11
XG4869 XI11_5/XI0/XI0_50/d_10_ XI11_5/XI0/XI0_50/d__10_ DECAP_INV_G11
XG4870 XI11_5/XI0/XI0_50/d_9_ XI11_5/XI0/XI0_50/d__9_ DECAP_INV_G11
XG4871 XI11_5/XI0/XI0_50/d_8_ XI11_5/XI0/XI0_50/d__8_ DECAP_INV_G11
XG4872 XI11_5/XI0/XI0_50/d_7_ XI11_5/XI0/XI0_50/d__7_ DECAP_INV_G11
XG4873 XI11_5/XI0/XI0_50/d_6_ XI11_5/XI0/XI0_50/d__6_ DECAP_INV_G11
XG4874 XI11_5/XI0/XI0_50/d_5_ XI11_5/XI0/XI0_50/d__5_ DECAP_INV_G11
XG4875 XI11_5/XI0/XI0_50/d_4_ XI11_5/XI0/XI0_50/d__4_ DECAP_INV_G11
XG4876 XI11_5/XI0/XI0_50/d_3_ XI11_5/XI0/XI0_50/d__3_ DECAP_INV_G11
XG4877 XI11_5/XI0/XI0_50/d_2_ XI11_5/XI0/XI0_50/d__2_ DECAP_INV_G11
XG4878 XI11_5/XI0/XI0_50/d_1_ XI11_5/XI0/XI0_50/d__1_ DECAP_INV_G11
XG4879 XI11_5/XI0/XI0_50/d_0_ XI11_5/XI0/XI0_50/d__0_ DECAP_INV_G11
XG4880 XI11_5/XI0/XI0_49/d__15_ XI11_5/XI0/XI0_49/d_15_ DECAP_INV_G11
XG4881 XI11_5/XI0/XI0_49/d__14_ XI11_5/XI0/XI0_49/d_14_ DECAP_INV_G11
XG4882 XI11_5/XI0/XI0_49/d__13_ XI11_5/XI0/XI0_49/d_13_ DECAP_INV_G11
XG4883 XI11_5/XI0/XI0_49/d__12_ XI11_5/XI0/XI0_49/d_12_ DECAP_INV_G11
XG4884 XI11_5/XI0/XI0_49/d__11_ XI11_5/XI0/XI0_49/d_11_ DECAP_INV_G11
XG4885 XI11_5/XI0/XI0_49/d__10_ XI11_5/XI0/XI0_49/d_10_ DECAP_INV_G11
XG4886 XI11_5/XI0/XI0_49/d__9_ XI11_5/XI0/XI0_49/d_9_ DECAP_INV_G11
XG4887 XI11_5/XI0/XI0_49/d__8_ XI11_5/XI0/XI0_49/d_8_ DECAP_INV_G11
XG4888 XI11_5/XI0/XI0_49/d__7_ XI11_5/XI0/XI0_49/d_7_ DECAP_INV_G11
XG4889 XI11_5/XI0/XI0_49/d__6_ XI11_5/XI0/XI0_49/d_6_ DECAP_INV_G11
XG4890 XI11_5/XI0/XI0_49/d__5_ XI11_5/XI0/XI0_49/d_5_ DECAP_INV_G11
XG4891 XI11_5/XI0/XI0_49/d__4_ XI11_5/XI0/XI0_49/d_4_ DECAP_INV_G11
XG4892 XI11_5/XI0/XI0_49/d__3_ XI11_5/XI0/XI0_49/d_3_ DECAP_INV_G11
XG4893 XI11_5/XI0/XI0_49/d__2_ XI11_5/XI0/XI0_49/d_2_ DECAP_INV_G11
XG4894 XI11_5/XI0/XI0_49/d__1_ XI11_5/XI0/XI0_49/d_1_ DECAP_INV_G11
XG4895 XI11_5/XI0/XI0_49/d__0_ XI11_5/XI0/XI0_49/d_0_ DECAP_INV_G11
XG4896 XI11_5/XI0/XI0_49/d_15_ XI11_5/XI0/XI0_49/d__15_ DECAP_INV_G11
XG4897 XI11_5/XI0/XI0_49/d_14_ XI11_5/XI0/XI0_49/d__14_ DECAP_INV_G11
XG4898 XI11_5/XI0/XI0_49/d_13_ XI11_5/XI0/XI0_49/d__13_ DECAP_INV_G11
XG4899 XI11_5/XI0/XI0_49/d_12_ XI11_5/XI0/XI0_49/d__12_ DECAP_INV_G11
XG4900 XI11_5/XI0/XI0_49/d_11_ XI11_5/XI0/XI0_49/d__11_ DECAP_INV_G11
XG4901 XI11_5/XI0/XI0_49/d_10_ XI11_5/XI0/XI0_49/d__10_ DECAP_INV_G11
XG4902 XI11_5/XI0/XI0_49/d_9_ XI11_5/XI0/XI0_49/d__9_ DECAP_INV_G11
XG4903 XI11_5/XI0/XI0_49/d_8_ XI11_5/XI0/XI0_49/d__8_ DECAP_INV_G11
XG4904 XI11_5/XI0/XI0_49/d_7_ XI11_5/XI0/XI0_49/d__7_ DECAP_INV_G11
XG4905 XI11_5/XI0/XI0_49/d_6_ XI11_5/XI0/XI0_49/d__6_ DECAP_INV_G11
XG4906 XI11_5/XI0/XI0_49/d_5_ XI11_5/XI0/XI0_49/d__5_ DECAP_INV_G11
XG4907 XI11_5/XI0/XI0_49/d_4_ XI11_5/XI0/XI0_49/d__4_ DECAP_INV_G11
XG4908 XI11_5/XI0/XI0_49/d_3_ XI11_5/XI0/XI0_49/d__3_ DECAP_INV_G11
XG4909 XI11_5/XI0/XI0_49/d_2_ XI11_5/XI0/XI0_49/d__2_ DECAP_INV_G11
XG4910 XI11_5/XI0/XI0_49/d_1_ XI11_5/XI0/XI0_49/d__1_ DECAP_INV_G11
XG4911 XI11_5/XI0/XI0_49/d_0_ XI11_5/XI0/XI0_49/d__0_ DECAP_INV_G11
XG4912 XI11_5/XI0/XI0_48/d__15_ XI11_5/XI0/XI0_48/d_15_ DECAP_INV_G11
XG4913 XI11_5/XI0/XI0_48/d__14_ XI11_5/XI0/XI0_48/d_14_ DECAP_INV_G11
XG4914 XI11_5/XI0/XI0_48/d__13_ XI11_5/XI0/XI0_48/d_13_ DECAP_INV_G11
XG4915 XI11_5/XI0/XI0_48/d__12_ XI11_5/XI0/XI0_48/d_12_ DECAP_INV_G11
XG4916 XI11_5/XI0/XI0_48/d__11_ XI11_5/XI0/XI0_48/d_11_ DECAP_INV_G11
XG4917 XI11_5/XI0/XI0_48/d__10_ XI11_5/XI0/XI0_48/d_10_ DECAP_INV_G11
XG4918 XI11_5/XI0/XI0_48/d__9_ XI11_5/XI0/XI0_48/d_9_ DECAP_INV_G11
XG4919 XI11_5/XI0/XI0_48/d__8_ XI11_5/XI0/XI0_48/d_8_ DECAP_INV_G11
XG4920 XI11_5/XI0/XI0_48/d__7_ XI11_5/XI0/XI0_48/d_7_ DECAP_INV_G11
XG4921 XI11_5/XI0/XI0_48/d__6_ XI11_5/XI0/XI0_48/d_6_ DECAP_INV_G11
XG4922 XI11_5/XI0/XI0_48/d__5_ XI11_5/XI0/XI0_48/d_5_ DECAP_INV_G11
XG4923 XI11_5/XI0/XI0_48/d__4_ XI11_5/XI0/XI0_48/d_4_ DECAP_INV_G11
XG4924 XI11_5/XI0/XI0_48/d__3_ XI11_5/XI0/XI0_48/d_3_ DECAP_INV_G11
XG4925 XI11_5/XI0/XI0_48/d__2_ XI11_5/XI0/XI0_48/d_2_ DECAP_INV_G11
XG4926 XI11_5/XI0/XI0_48/d__1_ XI11_5/XI0/XI0_48/d_1_ DECAP_INV_G11
XG4927 XI11_5/XI0/XI0_48/d__0_ XI11_5/XI0/XI0_48/d_0_ DECAP_INV_G11
XG4928 XI11_5/XI0/XI0_48/d_15_ XI11_5/XI0/XI0_48/d__15_ DECAP_INV_G11
XG4929 XI11_5/XI0/XI0_48/d_14_ XI11_5/XI0/XI0_48/d__14_ DECAP_INV_G11
XG4930 XI11_5/XI0/XI0_48/d_13_ XI11_5/XI0/XI0_48/d__13_ DECAP_INV_G11
XG4931 XI11_5/XI0/XI0_48/d_12_ XI11_5/XI0/XI0_48/d__12_ DECAP_INV_G11
XG4932 XI11_5/XI0/XI0_48/d_11_ XI11_5/XI0/XI0_48/d__11_ DECAP_INV_G11
XG4933 XI11_5/XI0/XI0_48/d_10_ XI11_5/XI0/XI0_48/d__10_ DECAP_INV_G11
XG4934 XI11_5/XI0/XI0_48/d_9_ XI11_5/XI0/XI0_48/d__9_ DECAP_INV_G11
XG4935 XI11_5/XI0/XI0_48/d_8_ XI11_5/XI0/XI0_48/d__8_ DECAP_INV_G11
XG4936 XI11_5/XI0/XI0_48/d_7_ XI11_5/XI0/XI0_48/d__7_ DECAP_INV_G11
XG4937 XI11_5/XI0/XI0_48/d_6_ XI11_5/XI0/XI0_48/d__6_ DECAP_INV_G11
XG4938 XI11_5/XI0/XI0_48/d_5_ XI11_5/XI0/XI0_48/d__5_ DECAP_INV_G11
XG4939 XI11_5/XI0/XI0_48/d_4_ XI11_5/XI0/XI0_48/d__4_ DECAP_INV_G11
XG4940 XI11_5/XI0/XI0_48/d_3_ XI11_5/XI0/XI0_48/d__3_ DECAP_INV_G11
XG4941 XI11_5/XI0/XI0_48/d_2_ XI11_5/XI0/XI0_48/d__2_ DECAP_INV_G11
XG4942 XI11_5/XI0/XI0_48/d_1_ XI11_5/XI0/XI0_48/d__1_ DECAP_INV_G11
XG4943 XI11_5/XI0/XI0_48/d_0_ XI11_5/XI0/XI0_48/d__0_ DECAP_INV_G11
XG4944 XI11_5/XI0/XI0_47/d__15_ XI11_5/XI0/XI0_47/d_15_ DECAP_INV_G11
XG4945 XI11_5/XI0/XI0_47/d__14_ XI11_5/XI0/XI0_47/d_14_ DECAP_INV_G11
XG4946 XI11_5/XI0/XI0_47/d__13_ XI11_5/XI0/XI0_47/d_13_ DECAP_INV_G11
XG4947 XI11_5/XI0/XI0_47/d__12_ XI11_5/XI0/XI0_47/d_12_ DECAP_INV_G11
XG4948 XI11_5/XI0/XI0_47/d__11_ XI11_5/XI0/XI0_47/d_11_ DECAP_INV_G11
XG4949 XI11_5/XI0/XI0_47/d__10_ XI11_5/XI0/XI0_47/d_10_ DECAP_INV_G11
XG4950 XI11_5/XI0/XI0_47/d__9_ XI11_5/XI0/XI0_47/d_9_ DECAP_INV_G11
XG4951 XI11_5/XI0/XI0_47/d__8_ XI11_5/XI0/XI0_47/d_8_ DECAP_INV_G11
XG4952 XI11_5/XI0/XI0_47/d__7_ XI11_5/XI0/XI0_47/d_7_ DECAP_INV_G11
XG4953 XI11_5/XI0/XI0_47/d__6_ XI11_5/XI0/XI0_47/d_6_ DECAP_INV_G11
XG4954 XI11_5/XI0/XI0_47/d__5_ XI11_5/XI0/XI0_47/d_5_ DECAP_INV_G11
XG4955 XI11_5/XI0/XI0_47/d__4_ XI11_5/XI0/XI0_47/d_4_ DECAP_INV_G11
XG4956 XI11_5/XI0/XI0_47/d__3_ XI11_5/XI0/XI0_47/d_3_ DECAP_INV_G11
XG4957 XI11_5/XI0/XI0_47/d__2_ XI11_5/XI0/XI0_47/d_2_ DECAP_INV_G11
XG4958 XI11_5/XI0/XI0_47/d__1_ XI11_5/XI0/XI0_47/d_1_ DECAP_INV_G11
XG4959 XI11_5/XI0/XI0_47/d__0_ XI11_5/XI0/XI0_47/d_0_ DECAP_INV_G11
XG4960 XI11_5/XI0/XI0_47/d_15_ XI11_5/XI0/XI0_47/d__15_ DECAP_INV_G11
XG4961 XI11_5/XI0/XI0_47/d_14_ XI11_5/XI0/XI0_47/d__14_ DECAP_INV_G11
XG4962 XI11_5/XI0/XI0_47/d_13_ XI11_5/XI0/XI0_47/d__13_ DECAP_INV_G11
XG4963 XI11_5/XI0/XI0_47/d_12_ XI11_5/XI0/XI0_47/d__12_ DECAP_INV_G11
XG4964 XI11_5/XI0/XI0_47/d_11_ XI11_5/XI0/XI0_47/d__11_ DECAP_INV_G11
XG4965 XI11_5/XI0/XI0_47/d_10_ XI11_5/XI0/XI0_47/d__10_ DECAP_INV_G11
XG4966 XI11_5/XI0/XI0_47/d_9_ XI11_5/XI0/XI0_47/d__9_ DECAP_INV_G11
XG4967 XI11_5/XI0/XI0_47/d_8_ XI11_5/XI0/XI0_47/d__8_ DECAP_INV_G11
XG4968 XI11_5/XI0/XI0_47/d_7_ XI11_5/XI0/XI0_47/d__7_ DECAP_INV_G11
XG4969 XI11_5/XI0/XI0_47/d_6_ XI11_5/XI0/XI0_47/d__6_ DECAP_INV_G11
XG4970 XI11_5/XI0/XI0_47/d_5_ XI11_5/XI0/XI0_47/d__5_ DECAP_INV_G11
XG4971 XI11_5/XI0/XI0_47/d_4_ XI11_5/XI0/XI0_47/d__4_ DECAP_INV_G11
XG4972 XI11_5/XI0/XI0_47/d_3_ XI11_5/XI0/XI0_47/d__3_ DECAP_INV_G11
XG4973 XI11_5/XI0/XI0_47/d_2_ XI11_5/XI0/XI0_47/d__2_ DECAP_INV_G11
XG4974 XI11_5/XI0/XI0_47/d_1_ XI11_5/XI0/XI0_47/d__1_ DECAP_INV_G11
XG4975 XI11_5/XI0/XI0_47/d_0_ XI11_5/XI0/XI0_47/d__0_ DECAP_INV_G11
XG4976 XI11_5/XI0/XI0_46/d__15_ XI11_5/XI0/XI0_46/d_15_ DECAP_INV_G11
XG4977 XI11_5/XI0/XI0_46/d__14_ XI11_5/XI0/XI0_46/d_14_ DECAP_INV_G11
XG4978 XI11_5/XI0/XI0_46/d__13_ XI11_5/XI0/XI0_46/d_13_ DECAP_INV_G11
XG4979 XI11_5/XI0/XI0_46/d__12_ XI11_5/XI0/XI0_46/d_12_ DECAP_INV_G11
XG4980 XI11_5/XI0/XI0_46/d__11_ XI11_5/XI0/XI0_46/d_11_ DECAP_INV_G11
XG4981 XI11_5/XI0/XI0_46/d__10_ XI11_5/XI0/XI0_46/d_10_ DECAP_INV_G11
XG4982 XI11_5/XI0/XI0_46/d__9_ XI11_5/XI0/XI0_46/d_9_ DECAP_INV_G11
XG4983 XI11_5/XI0/XI0_46/d__8_ XI11_5/XI0/XI0_46/d_8_ DECAP_INV_G11
XG4984 XI11_5/XI0/XI0_46/d__7_ XI11_5/XI0/XI0_46/d_7_ DECAP_INV_G11
XG4985 XI11_5/XI0/XI0_46/d__6_ XI11_5/XI0/XI0_46/d_6_ DECAP_INV_G11
XG4986 XI11_5/XI0/XI0_46/d__5_ XI11_5/XI0/XI0_46/d_5_ DECAP_INV_G11
XG4987 XI11_5/XI0/XI0_46/d__4_ XI11_5/XI0/XI0_46/d_4_ DECAP_INV_G11
XG4988 XI11_5/XI0/XI0_46/d__3_ XI11_5/XI0/XI0_46/d_3_ DECAP_INV_G11
XG4989 XI11_5/XI0/XI0_46/d__2_ XI11_5/XI0/XI0_46/d_2_ DECAP_INV_G11
XG4990 XI11_5/XI0/XI0_46/d__1_ XI11_5/XI0/XI0_46/d_1_ DECAP_INV_G11
XG4991 XI11_5/XI0/XI0_46/d__0_ XI11_5/XI0/XI0_46/d_0_ DECAP_INV_G11
XG4992 XI11_5/XI0/XI0_46/d_15_ XI11_5/XI0/XI0_46/d__15_ DECAP_INV_G11
XG4993 XI11_5/XI0/XI0_46/d_14_ XI11_5/XI0/XI0_46/d__14_ DECAP_INV_G11
XG4994 XI11_5/XI0/XI0_46/d_13_ XI11_5/XI0/XI0_46/d__13_ DECAP_INV_G11
XG4995 XI11_5/XI0/XI0_46/d_12_ XI11_5/XI0/XI0_46/d__12_ DECAP_INV_G11
XG4996 XI11_5/XI0/XI0_46/d_11_ XI11_5/XI0/XI0_46/d__11_ DECAP_INV_G11
XG4997 XI11_5/XI0/XI0_46/d_10_ XI11_5/XI0/XI0_46/d__10_ DECAP_INV_G11
XG4998 XI11_5/XI0/XI0_46/d_9_ XI11_5/XI0/XI0_46/d__9_ DECAP_INV_G11
XG4999 XI11_5/XI0/XI0_46/d_8_ XI11_5/XI0/XI0_46/d__8_ DECAP_INV_G11
XG5000 XI11_5/XI0/XI0_46/d_7_ XI11_5/XI0/XI0_46/d__7_ DECAP_INV_G11
XG5001 XI11_5/XI0/XI0_46/d_6_ XI11_5/XI0/XI0_46/d__6_ DECAP_INV_G11
XG5002 XI11_5/XI0/XI0_46/d_5_ XI11_5/XI0/XI0_46/d__5_ DECAP_INV_G11
XG5003 XI11_5/XI0/XI0_46/d_4_ XI11_5/XI0/XI0_46/d__4_ DECAP_INV_G11
XG5004 XI11_5/XI0/XI0_46/d_3_ XI11_5/XI0/XI0_46/d__3_ DECAP_INV_G11
XG5005 XI11_5/XI0/XI0_46/d_2_ XI11_5/XI0/XI0_46/d__2_ DECAP_INV_G11
XG5006 XI11_5/XI0/XI0_46/d_1_ XI11_5/XI0/XI0_46/d__1_ DECAP_INV_G11
XG5007 XI11_5/XI0/XI0_46/d_0_ XI11_5/XI0/XI0_46/d__0_ DECAP_INV_G11
XG5008 XI11_5/XI0/XI0_45/d__15_ XI11_5/XI0/XI0_45/d_15_ DECAP_INV_G11
XG5009 XI11_5/XI0/XI0_45/d__14_ XI11_5/XI0/XI0_45/d_14_ DECAP_INV_G11
XG5010 XI11_5/XI0/XI0_45/d__13_ XI11_5/XI0/XI0_45/d_13_ DECAP_INV_G11
XG5011 XI11_5/XI0/XI0_45/d__12_ XI11_5/XI0/XI0_45/d_12_ DECAP_INV_G11
XG5012 XI11_5/XI0/XI0_45/d__11_ XI11_5/XI0/XI0_45/d_11_ DECAP_INV_G11
XG5013 XI11_5/XI0/XI0_45/d__10_ XI11_5/XI0/XI0_45/d_10_ DECAP_INV_G11
XG5014 XI11_5/XI0/XI0_45/d__9_ XI11_5/XI0/XI0_45/d_9_ DECAP_INV_G11
XG5015 XI11_5/XI0/XI0_45/d__8_ XI11_5/XI0/XI0_45/d_8_ DECAP_INV_G11
XG5016 XI11_5/XI0/XI0_45/d__7_ XI11_5/XI0/XI0_45/d_7_ DECAP_INV_G11
XG5017 XI11_5/XI0/XI0_45/d__6_ XI11_5/XI0/XI0_45/d_6_ DECAP_INV_G11
XG5018 XI11_5/XI0/XI0_45/d__5_ XI11_5/XI0/XI0_45/d_5_ DECAP_INV_G11
XG5019 XI11_5/XI0/XI0_45/d__4_ XI11_5/XI0/XI0_45/d_4_ DECAP_INV_G11
XG5020 XI11_5/XI0/XI0_45/d__3_ XI11_5/XI0/XI0_45/d_3_ DECAP_INV_G11
XG5021 XI11_5/XI0/XI0_45/d__2_ XI11_5/XI0/XI0_45/d_2_ DECAP_INV_G11
XG5022 XI11_5/XI0/XI0_45/d__1_ XI11_5/XI0/XI0_45/d_1_ DECAP_INV_G11
XG5023 XI11_5/XI0/XI0_45/d__0_ XI11_5/XI0/XI0_45/d_0_ DECAP_INV_G11
XG5024 XI11_5/XI0/XI0_45/d_15_ XI11_5/XI0/XI0_45/d__15_ DECAP_INV_G11
XG5025 XI11_5/XI0/XI0_45/d_14_ XI11_5/XI0/XI0_45/d__14_ DECAP_INV_G11
XG5026 XI11_5/XI0/XI0_45/d_13_ XI11_5/XI0/XI0_45/d__13_ DECAP_INV_G11
XG5027 XI11_5/XI0/XI0_45/d_12_ XI11_5/XI0/XI0_45/d__12_ DECAP_INV_G11
XG5028 XI11_5/XI0/XI0_45/d_11_ XI11_5/XI0/XI0_45/d__11_ DECAP_INV_G11
XG5029 XI11_5/XI0/XI0_45/d_10_ XI11_5/XI0/XI0_45/d__10_ DECAP_INV_G11
XG5030 XI11_5/XI0/XI0_45/d_9_ XI11_5/XI0/XI0_45/d__9_ DECAP_INV_G11
XG5031 XI11_5/XI0/XI0_45/d_8_ XI11_5/XI0/XI0_45/d__8_ DECAP_INV_G11
XG5032 XI11_5/XI0/XI0_45/d_7_ XI11_5/XI0/XI0_45/d__7_ DECAP_INV_G11
XG5033 XI11_5/XI0/XI0_45/d_6_ XI11_5/XI0/XI0_45/d__6_ DECAP_INV_G11
XG5034 XI11_5/XI0/XI0_45/d_5_ XI11_5/XI0/XI0_45/d__5_ DECAP_INV_G11
XG5035 XI11_5/XI0/XI0_45/d_4_ XI11_5/XI0/XI0_45/d__4_ DECAP_INV_G11
XG5036 XI11_5/XI0/XI0_45/d_3_ XI11_5/XI0/XI0_45/d__3_ DECAP_INV_G11
XG5037 XI11_5/XI0/XI0_45/d_2_ XI11_5/XI0/XI0_45/d__2_ DECAP_INV_G11
XG5038 XI11_5/XI0/XI0_45/d_1_ XI11_5/XI0/XI0_45/d__1_ DECAP_INV_G11
XG5039 XI11_5/XI0/XI0_45/d_0_ XI11_5/XI0/XI0_45/d__0_ DECAP_INV_G11
XG5040 XI11_5/XI0/XI0_44/d__15_ XI11_5/XI0/XI0_44/d_15_ DECAP_INV_G11
XG5041 XI11_5/XI0/XI0_44/d__14_ XI11_5/XI0/XI0_44/d_14_ DECAP_INV_G11
XG5042 XI11_5/XI0/XI0_44/d__13_ XI11_5/XI0/XI0_44/d_13_ DECAP_INV_G11
XG5043 XI11_5/XI0/XI0_44/d__12_ XI11_5/XI0/XI0_44/d_12_ DECAP_INV_G11
XG5044 XI11_5/XI0/XI0_44/d__11_ XI11_5/XI0/XI0_44/d_11_ DECAP_INV_G11
XG5045 XI11_5/XI0/XI0_44/d__10_ XI11_5/XI0/XI0_44/d_10_ DECAP_INV_G11
XG5046 XI11_5/XI0/XI0_44/d__9_ XI11_5/XI0/XI0_44/d_9_ DECAP_INV_G11
XG5047 XI11_5/XI0/XI0_44/d__8_ XI11_5/XI0/XI0_44/d_8_ DECAP_INV_G11
XG5048 XI11_5/XI0/XI0_44/d__7_ XI11_5/XI0/XI0_44/d_7_ DECAP_INV_G11
XG5049 XI11_5/XI0/XI0_44/d__6_ XI11_5/XI0/XI0_44/d_6_ DECAP_INV_G11
XG5050 XI11_5/XI0/XI0_44/d__5_ XI11_5/XI0/XI0_44/d_5_ DECAP_INV_G11
XG5051 XI11_5/XI0/XI0_44/d__4_ XI11_5/XI0/XI0_44/d_4_ DECAP_INV_G11
XG5052 XI11_5/XI0/XI0_44/d__3_ XI11_5/XI0/XI0_44/d_3_ DECAP_INV_G11
XG5053 XI11_5/XI0/XI0_44/d__2_ XI11_5/XI0/XI0_44/d_2_ DECAP_INV_G11
XG5054 XI11_5/XI0/XI0_44/d__1_ XI11_5/XI0/XI0_44/d_1_ DECAP_INV_G11
XG5055 XI11_5/XI0/XI0_44/d__0_ XI11_5/XI0/XI0_44/d_0_ DECAP_INV_G11
XG5056 XI11_5/XI0/XI0_44/d_15_ XI11_5/XI0/XI0_44/d__15_ DECAP_INV_G11
XG5057 XI11_5/XI0/XI0_44/d_14_ XI11_5/XI0/XI0_44/d__14_ DECAP_INV_G11
XG5058 XI11_5/XI0/XI0_44/d_13_ XI11_5/XI0/XI0_44/d__13_ DECAP_INV_G11
XG5059 XI11_5/XI0/XI0_44/d_12_ XI11_5/XI0/XI0_44/d__12_ DECAP_INV_G11
XG5060 XI11_5/XI0/XI0_44/d_11_ XI11_5/XI0/XI0_44/d__11_ DECAP_INV_G11
XG5061 XI11_5/XI0/XI0_44/d_10_ XI11_5/XI0/XI0_44/d__10_ DECAP_INV_G11
XG5062 XI11_5/XI0/XI0_44/d_9_ XI11_5/XI0/XI0_44/d__9_ DECAP_INV_G11
XG5063 XI11_5/XI0/XI0_44/d_8_ XI11_5/XI0/XI0_44/d__8_ DECAP_INV_G11
XG5064 XI11_5/XI0/XI0_44/d_7_ XI11_5/XI0/XI0_44/d__7_ DECAP_INV_G11
XG5065 XI11_5/XI0/XI0_44/d_6_ XI11_5/XI0/XI0_44/d__6_ DECAP_INV_G11
XG5066 XI11_5/XI0/XI0_44/d_5_ XI11_5/XI0/XI0_44/d__5_ DECAP_INV_G11
XG5067 XI11_5/XI0/XI0_44/d_4_ XI11_5/XI0/XI0_44/d__4_ DECAP_INV_G11
XG5068 XI11_5/XI0/XI0_44/d_3_ XI11_5/XI0/XI0_44/d__3_ DECAP_INV_G11
XG5069 XI11_5/XI0/XI0_44/d_2_ XI11_5/XI0/XI0_44/d__2_ DECAP_INV_G11
XG5070 XI11_5/XI0/XI0_44/d_1_ XI11_5/XI0/XI0_44/d__1_ DECAP_INV_G11
XG5071 XI11_5/XI0/XI0_44/d_0_ XI11_5/XI0/XI0_44/d__0_ DECAP_INV_G11
XG5072 XI11_5/XI0/XI0_43/d__15_ XI11_5/XI0/XI0_43/d_15_ DECAP_INV_G11
XG5073 XI11_5/XI0/XI0_43/d__14_ XI11_5/XI0/XI0_43/d_14_ DECAP_INV_G11
XG5074 XI11_5/XI0/XI0_43/d__13_ XI11_5/XI0/XI0_43/d_13_ DECAP_INV_G11
XG5075 XI11_5/XI0/XI0_43/d__12_ XI11_5/XI0/XI0_43/d_12_ DECAP_INV_G11
XG5076 XI11_5/XI0/XI0_43/d__11_ XI11_5/XI0/XI0_43/d_11_ DECAP_INV_G11
XG5077 XI11_5/XI0/XI0_43/d__10_ XI11_5/XI0/XI0_43/d_10_ DECAP_INV_G11
XG5078 XI11_5/XI0/XI0_43/d__9_ XI11_5/XI0/XI0_43/d_9_ DECAP_INV_G11
XG5079 XI11_5/XI0/XI0_43/d__8_ XI11_5/XI0/XI0_43/d_8_ DECAP_INV_G11
XG5080 XI11_5/XI0/XI0_43/d__7_ XI11_5/XI0/XI0_43/d_7_ DECAP_INV_G11
XG5081 XI11_5/XI0/XI0_43/d__6_ XI11_5/XI0/XI0_43/d_6_ DECAP_INV_G11
XG5082 XI11_5/XI0/XI0_43/d__5_ XI11_5/XI0/XI0_43/d_5_ DECAP_INV_G11
XG5083 XI11_5/XI0/XI0_43/d__4_ XI11_5/XI0/XI0_43/d_4_ DECAP_INV_G11
XG5084 XI11_5/XI0/XI0_43/d__3_ XI11_5/XI0/XI0_43/d_3_ DECAP_INV_G11
XG5085 XI11_5/XI0/XI0_43/d__2_ XI11_5/XI0/XI0_43/d_2_ DECAP_INV_G11
XG5086 XI11_5/XI0/XI0_43/d__1_ XI11_5/XI0/XI0_43/d_1_ DECAP_INV_G11
XG5087 XI11_5/XI0/XI0_43/d__0_ XI11_5/XI0/XI0_43/d_0_ DECAP_INV_G11
XG5088 XI11_5/XI0/XI0_43/d_15_ XI11_5/XI0/XI0_43/d__15_ DECAP_INV_G11
XG5089 XI11_5/XI0/XI0_43/d_14_ XI11_5/XI0/XI0_43/d__14_ DECAP_INV_G11
XG5090 XI11_5/XI0/XI0_43/d_13_ XI11_5/XI0/XI0_43/d__13_ DECAP_INV_G11
XG5091 XI11_5/XI0/XI0_43/d_12_ XI11_5/XI0/XI0_43/d__12_ DECAP_INV_G11
XG5092 XI11_5/XI0/XI0_43/d_11_ XI11_5/XI0/XI0_43/d__11_ DECAP_INV_G11
XG5093 XI11_5/XI0/XI0_43/d_10_ XI11_5/XI0/XI0_43/d__10_ DECAP_INV_G11
XG5094 XI11_5/XI0/XI0_43/d_9_ XI11_5/XI0/XI0_43/d__9_ DECAP_INV_G11
XG5095 XI11_5/XI0/XI0_43/d_8_ XI11_5/XI0/XI0_43/d__8_ DECAP_INV_G11
XG5096 XI11_5/XI0/XI0_43/d_7_ XI11_5/XI0/XI0_43/d__7_ DECAP_INV_G11
XG5097 XI11_5/XI0/XI0_43/d_6_ XI11_5/XI0/XI0_43/d__6_ DECAP_INV_G11
XG5098 XI11_5/XI0/XI0_43/d_5_ XI11_5/XI0/XI0_43/d__5_ DECAP_INV_G11
XG5099 XI11_5/XI0/XI0_43/d_4_ XI11_5/XI0/XI0_43/d__4_ DECAP_INV_G11
XG5100 XI11_5/XI0/XI0_43/d_3_ XI11_5/XI0/XI0_43/d__3_ DECAP_INV_G11
XG5101 XI11_5/XI0/XI0_43/d_2_ XI11_5/XI0/XI0_43/d__2_ DECAP_INV_G11
XG5102 XI11_5/XI0/XI0_43/d_1_ XI11_5/XI0/XI0_43/d__1_ DECAP_INV_G11
XG5103 XI11_5/XI0/XI0_43/d_0_ XI11_5/XI0/XI0_43/d__0_ DECAP_INV_G11
XG5104 XI11_5/XI0/XI0_42/d__15_ XI11_5/XI0/XI0_42/d_15_ DECAP_INV_G11
XG5105 XI11_5/XI0/XI0_42/d__14_ XI11_5/XI0/XI0_42/d_14_ DECAP_INV_G11
XG5106 XI11_5/XI0/XI0_42/d__13_ XI11_5/XI0/XI0_42/d_13_ DECAP_INV_G11
XG5107 XI11_5/XI0/XI0_42/d__12_ XI11_5/XI0/XI0_42/d_12_ DECAP_INV_G11
XG5108 XI11_5/XI0/XI0_42/d__11_ XI11_5/XI0/XI0_42/d_11_ DECAP_INV_G11
XG5109 XI11_5/XI0/XI0_42/d__10_ XI11_5/XI0/XI0_42/d_10_ DECAP_INV_G11
XG5110 XI11_5/XI0/XI0_42/d__9_ XI11_5/XI0/XI0_42/d_9_ DECAP_INV_G11
XG5111 XI11_5/XI0/XI0_42/d__8_ XI11_5/XI0/XI0_42/d_8_ DECAP_INV_G11
XG5112 XI11_5/XI0/XI0_42/d__7_ XI11_5/XI0/XI0_42/d_7_ DECAP_INV_G11
XG5113 XI11_5/XI0/XI0_42/d__6_ XI11_5/XI0/XI0_42/d_6_ DECAP_INV_G11
XG5114 XI11_5/XI0/XI0_42/d__5_ XI11_5/XI0/XI0_42/d_5_ DECAP_INV_G11
XG5115 XI11_5/XI0/XI0_42/d__4_ XI11_5/XI0/XI0_42/d_4_ DECAP_INV_G11
XG5116 XI11_5/XI0/XI0_42/d__3_ XI11_5/XI0/XI0_42/d_3_ DECAP_INV_G11
XG5117 XI11_5/XI0/XI0_42/d__2_ XI11_5/XI0/XI0_42/d_2_ DECAP_INV_G11
XG5118 XI11_5/XI0/XI0_42/d__1_ XI11_5/XI0/XI0_42/d_1_ DECAP_INV_G11
XG5119 XI11_5/XI0/XI0_42/d__0_ XI11_5/XI0/XI0_42/d_0_ DECAP_INV_G11
XG5120 XI11_5/XI0/XI0_42/d_15_ XI11_5/XI0/XI0_42/d__15_ DECAP_INV_G11
XG5121 XI11_5/XI0/XI0_42/d_14_ XI11_5/XI0/XI0_42/d__14_ DECAP_INV_G11
XG5122 XI11_5/XI0/XI0_42/d_13_ XI11_5/XI0/XI0_42/d__13_ DECAP_INV_G11
XG5123 XI11_5/XI0/XI0_42/d_12_ XI11_5/XI0/XI0_42/d__12_ DECAP_INV_G11
XG5124 XI11_5/XI0/XI0_42/d_11_ XI11_5/XI0/XI0_42/d__11_ DECAP_INV_G11
XG5125 XI11_5/XI0/XI0_42/d_10_ XI11_5/XI0/XI0_42/d__10_ DECAP_INV_G11
XG5126 XI11_5/XI0/XI0_42/d_9_ XI11_5/XI0/XI0_42/d__9_ DECAP_INV_G11
XG5127 XI11_5/XI0/XI0_42/d_8_ XI11_5/XI0/XI0_42/d__8_ DECAP_INV_G11
XG5128 XI11_5/XI0/XI0_42/d_7_ XI11_5/XI0/XI0_42/d__7_ DECAP_INV_G11
XG5129 XI11_5/XI0/XI0_42/d_6_ XI11_5/XI0/XI0_42/d__6_ DECAP_INV_G11
XG5130 XI11_5/XI0/XI0_42/d_5_ XI11_5/XI0/XI0_42/d__5_ DECAP_INV_G11
XG5131 XI11_5/XI0/XI0_42/d_4_ XI11_5/XI0/XI0_42/d__4_ DECAP_INV_G11
XG5132 XI11_5/XI0/XI0_42/d_3_ XI11_5/XI0/XI0_42/d__3_ DECAP_INV_G11
XG5133 XI11_5/XI0/XI0_42/d_2_ XI11_5/XI0/XI0_42/d__2_ DECAP_INV_G11
XG5134 XI11_5/XI0/XI0_42/d_1_ XI11_5/XI0/XI0_42/d__1_ DECAP_INV_G11
XG5135 XI11_5/XI0/XI0_42/d_0_ XI11_5/XI0/XI0_42/d__0_ DECAP_INV_G11
XG5136 XI11_5/XI0/XI0_41/d__15_ XI11_5/XI0/XI0_41/d_15_ DECAP_INV_G11
XG5137 XI11_5/XI0/XI0_41/d__14_ XI11_5/XI0/XI0_41/d_14_ DECAP_INV_G11
XG5138 XI11_5/XI0/XI0_41/d__13_ XI11_5/XI0/XI0_41/d_13_ DECAP_INV_G11
XG5139 XI11_5/XI0/XI0_41/d__12_ XI11_5/XI0/XI0_41/d_12_ DECAP_INV_G11
XG5140 XI11_5/XI0/XI0_41/d__11_ XI11_5/XI0/XI0_41/d_11_ DECAP_INV_G11
XG5141 XI11_5/XI0/XI0_41/d__10_ XI11_5/XI0/XI0_41/d_10_ DECAP_INV_G11
XG5142 XI11_5/XI0/XI0_41/d__9_ XI11_5/XI0/XI0_41/d_9_ DECAP_INV_G11
XG5143 XI11_5/XI0/XI0_41/d__8_ XI11_5/XI0/XI0_41/d_8_ DECAP_INV_G11
XG5144 XI11_5/XI0/XI0_41/d__7_ XI11_5/XI0/XI0_41/d_7_ DECAP_INV_G11
XG5145 XI11_5/XI0/XI0_41/d__6_ XI11_5/XI0/XI0_41/d_6_ DECAP_INV_G11
XG5146 XI11_5/XI0/XI0_41/d__5_ XI11_5/XI0/XI0_41/d_5_ DECAP_INV_G11
XG5147 XI11_5/XI0/XI0_41/d__4_ XI11_5/XI0/XI0_41/d_4_ DECAP_INV_G11
XG5148 XI11_5/XI0/XI0_41/d__3_ XI11_5/XI0/XI0_41/d_3_ DECAP_INV_G11
XG5149 XI11_5/XI0/XI0_41/d__2_ XI11_5/XI0/XI0_41/d_2_ DECAP_INV_G11
XG5150 XI11_5/XI0/XI0_41/d__1_ XI11_5/XI0/XI0_41/d_1_ DECAP_INV_G11
XG5151 XI11_5/XI0/XI0_41/d__0_ XI11_5/XI0/XI0_41/d_0_ DECAP_INV_G11
XG5152 XI11_5/XI0/XI0_41/d_15_ XI11_5/XI0/XI0_41/d__15_ DECAP_INV_G11
XG5153 XI11_5/XI0/XI0_41/d_14_ XI11_5/XI0/XI0_41/d__14_ DECAP_INV_G11
XG5154 XI11_5/XI0/XI0_41/d_13_ XI11_5/XI0/XI0_41/d__13_ DECAP_INV_G11
XG5155 XI11_5/XI0/XI0_41/d_12_ XI11_5/XI0/XI0_41/d__12_ DECAP_INV_G11
XG5156 XI11_5/XI0/XI0_41/d_11_ XI11_5/XI0/XI0_41/d__11_ DECAP_INV_G11
XG5157 XI11_5/XI0/XI0_41/d_10_ XI11_5/XI0/XI0_41/d__10_ DECAP_INV_G11
XG5158 XI11_5/XI0/XI0_41/d_9_ XI11_5/XI0/XI0_41/d__9_ DECAP_INV_G11
XG5159 XI11_5/XI0/XI0_41/d_8_ XI11_5/XI0/XI0_41/d__8_ DECAP_INV_G11
XG5160 XI11_5/XI0/XI0_41/d_7_ XI11_5/XI0/XI0_41/d__7_ DECAP_INV_G11
XG5161 XI11_5/XI0/XI0_41/d_6_ XI11_5/XI0/XI0_41/d__6_ DECAP_INV_G11
XG5162 XI11_5/XI0/XI0_41/d_5_ XI11_5/XI0/XI0_41/d__5_ DECAP_INV_G11
XG5163 XI11_5/XI0/XI0_41/d_4_ XI11_5/XI0/XI0_41/d__4_ DECAP_INV_G11
XG5164 XI11_5/XI0/XI0_41/d_3_ XI11_5/XI0/XI0_41/d__3_ DECAP_INV_G11
XG5165 XI11_5/XI0/XI0_41/d_2_ XI11_5/XI0/XI0_41/d__2_ DECAP_INV_G11
XG5166 XI11_5/XI0/XI0_41/d_1_ XI11_5/XI0/XI0_41/d__1_ DECAP_INV_G11
XG5167 XI11_5/XI0/XI0_41/d_0_ XI11_5/XI0/XI0_41/d__0_ DECAP_INV_G11
XG5168 XI11_5/XI0/XI0_40/d__15_ XI11_5/XI0/XI0_40/d_15_ DECAP_INV_G11
XG5169 XI11_5/XI0/XI0_40/d__14_ XI11_5/XI0/XI0_40/d_14_ DECAP_INV_G11
XG5170 XI11_5/XI0/XI0_40/d__13_ XI11_5/XI0/XI0_40/d_13_ DECAP_INV_G11
XG5171 XI11_5/XI0/XI0_40/d__12_ XI11_5/XI0/XI0_40/d_12_ DECAP_INV_G11
XG5172 XI11_5/XI0/XI0_40/d__11_ XI11_5/XI0/XI0_40/d_11_ DECAP_INV_G11
XG5173 XI11_5/XI0/XI0_40/d__10_ XI11_5/XI0/XI0_40/d_10_ DECAP_INV_G11
XG5174 XI11_5/XI0/XI0_40/d__9_ XI11_5/XI0/XI0_40/d_9_ DECAP_INV_G11
XG5175 XI11_5/XI0/XI0_40/d__8_ XI11_5/XI0/XI0_40/d_8_ DECAP_INV_G11
XG5176 XI11_5/XI0/XI0_40/d__7_ XI11_5/XI0/XI0_40/d_7_ DECAP_INV_G11
XG5177 XI11_5/XI0/XI0_40/d__6_ XI11_5/XI0/XI0_40/d_6_ DECAP_INV_G11
XG5178 XI11_5/XI0/XI0_40/d__5_ XI11_5/XI0/XI0_40/d_5_ DECAP_INV_G11
XG5179 XI11_5/XI0/XI0_40/d__4_ XI11_5/XI0/XI0_40/d_4_ DECAP_INV_G11
XG5180 XI11_5/XI0/XI0_40/d__3_ XI11_5/XI0/XI0_40/d_3_ DECAP_INV_G11
XG5181 XI11_5/XI0/XI0_40/d__2_ XI11_5/XI0/XI0_40/d_2_ DECAP_INV_G11
XG5182 XI11_5/XI0/XI0_40/d__1_ XI11_5/XI0/XI0_40/d_1_ DECAP_INV_G11
XG5183 XI11_5/XI0/XI0_40/d__0_ XI11_5/XI0/XI0_40/d_0_ DECAP_INV_G11
XG5184 XI11_5/XI0/XI0_40/d_15_ XI11_5/XI0/XI0_40/d__15_ DECAP_INV_G11
XG5185 XI11_5/XI0/XI0_40/d_14_ XI11_5/XI0/XI0_40/d__14_ DECAP_INV_G11
XG5186 XI11_5/XI0/XI0_40/d_13_ XI11_5/XI0/XI0_40/d__13_ DECAP_INV_G11
XG5187 XI11_5/XI0/XI0_40/d_12_ XI11_5/XI0/XI0_40/d__12_ DECAP_INV_G11
XG5188 XI11_5/XI0/XI0_40/d_11_ XI11_5/XI0/XI0_40/d__11_ DECAP_INV_G11
XG5189 XI11_5/XI0/XI0_40/d_10_ XI11_5/XI0/XI0_40/d__10_ DECAP_INV_G11
XG5190 XI11_5/XI0/XI0_40/d_9_ XI11_5/XI0/XI0_40/d__9_ DECAP_INV_G11
XG5191 XI11_5/XI0/XI0_40/d_8_ XI11_5/XI0/XI0_40/d__8_ DECAP_INV_G11
XG5192 XI11_5/XI0/XI0_40/d_7_ XI11_5/XI0/XI0_40/d__7_ DECAP_INV_G11
XG5193 XI11_5/XI0/XI0_40/d_6_ XI11_5/XI0/XI0_40/d__6_ DECAP_INV_G11
XG5194 XI11_5/XI0/XI0_40/d_5_ XI11_5/XI0/XI0_40/d__5_ DECAP_INV_G11
XG5195 XI11_5/XI0/XI0_40/d_4_ XI11_5/XI0/XI0_40/d__4_ DECAP_INV_G11
XG5196 XI11_5/XI0/XI0_40/d_3_ XI11_5/XI0/XI0_40/d__3_ DECAP_INV_G11
XG5197 XI11_5/XI0/XI0_40/d_2_ XI11_5/XI0/XI0_40/d__2_ DECAP_INV_G11
XG5198 XI11_5/XI0/XI0_40/d_1_ XI11_5/XI0/XI0_40/d__1_ DECAP_INV_G11
XG5199 XI11_5/XI0/XI0_40/d_0_ XI11_5/XI0/XI0_40/d__0_ DECAP_INV_G11
XG5200 XI11_5/XI0/XI0_39/d__15_ XI11_5/XI0/XI0_39/d_15_ DECAP_INV_G11
XG5201 XI11_5/XI0/XI0_39/d__14_ XI11_5/XI0/XI0_39/d_14_ DECAP_INV_G11
XG5202 XI11_5/XI0/XI0_39/d__13_ XI11_5/XI0/XI0_39/d_13_ DECAP_INV_G11
XG5203 XI11_5/XI0/XI0_39/d__12_ XI11_5/XI0/XI0_39/d_12_ DECAP_INV_G11
XG5204 XI11_5/XI0/XI0_39/d__11_ XI11_5/XI0/XI0_39/d_11_ DECAP_INV_G11
XG5205 XI11_5/XI0/XI0_39/d__10_ XI11_5/XI0/XI0_39/d_10_ DECAP_INV_G11
XG5206 XI11_5/XI0/XI0_39/d__9_ XI11_5/XI0/XI0_39/d_9_ DECAP_INV_G11
XG5207 XI11_5/XI0/XI0_39/d__8_ XI11_5/XI0/XI0_39/d_8_ DECAP_INV_G11
XG5208 XI11_5/XI0/XI0_39/d__7_ XI11_5/XI0/XI0_39/d_7_ DECAP_INV_G11
XG5209 XI11_5/XI0/XI0_39/d__6_ XI11_5/XI0/XI0_39/d_6_ DECAP_INV_G11
XG5210 XI11_5/XI0/XI0_39/d__5_ XI11_5/XI0/XI0_39/d_5_ DECAP_INV_G11
XG5211 XI11_5/XI0/XI0_39/d__4_ XI11_5/XI0/XI0_39/d_4_ DECAP_INV_G11
XG5212 XI11_5/XI0/XI0_39/d__3_ XI11_5/XI0/XI0_39/d_3_ DECAP_INV_G11
XG5213 XI11_5/XI0/XI0_39/d__2_ XI11_5/XI0/XI0_39/d_2_ DECAP_INV_G11
XG5214 XI11_5/XI0/XI0_39/d__1_ XI11_5/XI0/XI0_39/d_1_ DECAP_INV_G11
XG5215 XI11_5/XI0/XI0_39/d__0_ XI11_5/XI0/XI0_39/d_0_ DECAP_INV_G11
XG5216 XI11_5/XI0/XI0_39/d_15_ XI11_5/XI0/XI0_39/d__15_ DECAP_INV_G11
XG5217 XI11_5/XI0/XI0_39/d_14_ XI11_5/XI0/XI0_39/d__14_ DECAP_INV_G11
XG5218 XI11_5/XI0/XI0_39/d_13_ XI11_5/XI0/XI0_39/d__13_ DECAP_INV_G11
XG5219 XI11_5/XI0/XI0_39/d_12_ XI11_5/XI0/XI0_39/d__12_ DECAP_INV_G11
XG5220 XI11_5/XI0/XI0_39/d_11_ XI11_5/XI0/XI0_39/d__11_ DECAP_INV_G11
XG5221 XI11_5/XI0/XI0_39/d_10_ XI11_5/XI0/XI0_39/d__10_ DECAP_INV_G11
XG5222 XI11_5/XI0/XI0_39/d_9_ XI11_5/XI0/XI0_39/d__9_ DECAP_INV_G11
XG5223 XI11_5/XI0/XI0_39/d_8_ XI11_5/XI0/XI0_39/d__8_ DECAP_INV_G11
XG5224 XI11_5/XI0/XI0_39/d_7_ XI11_5/XI0/XI0_39/d__7_ DECAP_INV_G11
XG5225 XI11_5/XI0/XI0_39/d_6_ XI11_5/XI0/XI0_39/d__6_ DECAP_INV_G11
XG5226 XI11_5/XI0/XI0_39/d_5_ XI11_5/XI0/XI0_39/d__5_ DECAP_INV_G11
XG5227 XI11_5/XI0/XI0_39/d_4_ XI11_5/XI0/XI0_39/d__4_ DECAP_INV_G11
XG5228 XI11_5/XI0/XI0_39/d_3_ XI11_5/XI0/XI0_39/d__3_ DECAP_INV_G11
XG5229 XI11_5/XI0/XI0_39/d_2_ XI11_5/XI0/XI0_39/d__2_ DECAP_INV_G11
XG5230 XI11_5/XI0/XI0_39/d_1_ XI11_5/XI0/XI0_39/d__1_ DECAP_INV_G11
XG5231 XI11_5/XI0/XI0_39/d_0_ XI11_5/XI0/XI0_39/d__0_ DECAP_INV_G11
XG5232 XI11_5/XI0/XI0_38/d__15_ XI11_5/XI0/XI0_38/d_15_ DECAP_INV_G11
XG5233 XI11_5/XI0/XI0_38/d__14_ XI11_5/XI0/XI0_38/d_14_ DECAP_INV_G11
XG5234 XI11_5/XI0/XI0_38/d__13_ XI11_5/XI0/XI0_38/d_13_ DECAP_INV_G11
XG5235 XI11_5/XI0/XI0_38/d__12_ XI11_5/XI0/XI0_38/d_12_ DECAP_INV_G11
XG5236 XI11_5/XI0/XI0_38/d__11_ XI11_5/XI0/XI0_38/d_11_ DECAP_INV_G11
XG5237 XI11_5/XI0/XI0_38/d__10_ XI11_5/XI0/XI0_38/d_10_ DECAP_INV_G11
XG5238 XI11_5/XI0/XI0_38/d__9_ XI11_5/XI0/XI0_38/d_9_ DECAP_INV_G11
XG5239 XI11_5/XI0/XI0_38/d__8_ XI11_5/XI0/XI0_38/d_8_ DECAP_INV_G11
XG5240 XI11_5/XI0/XI0_38/d__7_ XI11_5/XI0/XI0_38/d_7_ DECAP_INV_G11
XG5241 XI11_5/XI0/XI0_38/d__6_ XI11_5/XI0/XI0_38/d_6_ DECAP_INV_G11
XG5242 XI11_5/XI0/XI0_38/d__5_ XI11_5/XI0/XI0_38/d_5_ DECAP_INV_G11
XG5243 XI11_5/XI0/XI0_38/d__4_ XI11_5/XI0/XI0_38/d_4_ DECAP_INV_G11
XG5244 XI11_5/XI0/XI0_38/d__3_ XI11_5/XI0/XI0_38/d_3_ DECAP_INV_G11
XG5245 XI11_5/XI0/XI0_38/d__2_ XI11_5/XI0/XI0_38/d_2_ DECAP_INV_G11
XG5246 XI11_5/XI0/XI0_38/d__1_ XI11_5/XI0/XI0_38/d_1_ DECAP_INV_G11
XG5247 XI11_5/XI0/XI0_38/d__0_ XI11_5/XI0/XI0_38/d_0_ DECAP_INV_G11
XG5248 XI11_5/XI0/XI0_38/d_15_ XI11_5/XI0/XI0_38/d__15_ DECAP_INV_G11
XG5249 XI11_5/XI0/XI0_38/d_14_ XI11_5/XI0/XI0_38/d__14_ DECAP_INV_G11
XG5250 XI11_5/XI0/XI0_38/d_13_ XI11_5/XI0/XI0_38/d__13_ DECAP_INV_G11
XG5251 XI11_5/XI0/XI0_38/d_12_ XI11_5/XI0/XI0_38/d__12_ DECAP_INV_G11
XG5252 XI11_5/XI0/XI0_38/d_11_ XI11_5/XI0/XI0_38/d__11_ DECAP_INV_G11
XG5253 XI11_5/XI0/XI0_38/d_10_ XI11_5/XI0/XI0_38/d__10_ DECAP_INV_G11
XG5254 XI11_5/XI0/XI0_38/d_9_ XI11_5/XI0/XI0_38/d__9_ DECAP_INV_G11
XG5255 XI11_5/XI0/XI0_38/d_8_ XI11_5/XI0/XI0_38/d__8_ DECAP_INV_G11
XG5256 XI11_5/XI0/XI0_38/d_7_ XI11_5/XI0/XI0_38/d__7_ DECAP_INV_G11
XG5257 XI11_5/XI0/XI0_38/d_6_ XI11_5/XI0/XI0_38/d__6_ DECAP_INV_G11
XG5258 XI11_5/XI0/XI0_38/d_5_ XI11_5/XI0/XI0_38/d__5_ DECAP_INV_G11
XG5259 XI11_5/XI0/XI0_38/d_4_ XI11_5/XI0/XI0_38/d__4_ DECAP_INV_G11
XG5260 XI11_5/XI0/XI0_38/d_3_ XI11_5/XI0/XI0_38/d__3_ DECAP_INV_G11
XG5261 XI11_5/XI0/XI0_38/d_2_ XI11_5/XI0/XI0_38/d__2_ DECAP_INV_G11
XG5262 XI11_5/XI0/XI0_38/d_1_ XI11_5/XI0/XI0_38/d__1_ DECAP_INV_G11
XG5263 XI11_5/XI0/XI0_38/d_0_ XI11_5/XI0/XI0_38/d__0_ DECAP_INV_G11
XG5264 XI11_5/XI0/XI0_37/d__15_ XI11_5/XI0/XI0_37/d_15_ DECAP_INV_G11
XG5265 XI11_5/XI0/XI0_37/d__14_ XI11_5/XI0/XI0_37/d_14_ DECAP_INV_G11
XG5266 XI11_5/XI0/XI0_37/d__13_ XI11_5/XI0/XI0_37/d_13_ DECAP_INV_G11
XG5267 XI11_5/XI0/XI0_37/d__12_ XI11_5/XI0/XI0_37/d_12_ DECAP_INV_G11
XG5268 XI11_5/XI0/XI0_37/d__11_ XI11_5/XI0/XI0_37/d_11_ DECAP_INV_G11
XG5269 XI11_5/XI0/XI0_37/d__10_ XI11_5/XI0/XI0_37/d_10_ DECAP_INV_G11
XG5270 XI11_5/XI0/XI0_37/d__9_ XI11_5/XI0/XI0_37/d_9_ DECAP_INV_G11
XG5271 XI11_5/XI0/XI0_37/d__8_ XI11_5/XI0/XI0_37/d_8_ DECAP_INV_G11
XG5272 XI11_5/XI0/XI0_37/d__7_ XI11_5/XI0/XI0_37/d_7_ DECAP_INV_G11
XG5273 XI11_5/XI0/XI0_37/d__6_ XI11_5/XI0/XI0_37/d_6_ DECAP_INV_G11
XG5274 XI11_5/XI0/XI0_37/d__5_ XI11_5/XI0/XI0_37/d_5_ DECAP_INV_G11
XG5275 XI11_5/XI0/XI0_37/d__4_ XI11_5/XI0/XI0_37/d_4_ DECAP_INV_G11
XG5276 XI11_5/XI0/XI0_37/d__3_ XI11_5/XI0/XI0_37/d_3_ DECAP_INV_G11
XG5277 XI11_5/XI0/XI0_37/d__2_ XI11_5/XI0/XI0_37/d_2_ DECAP_INV_G11
XG5278 XI11_5/XI0/XI0_37/d__1_ XI11_5/XI0/XI0_37/d_1_ DECAP_INV_G11
XG5279 XI11_5/XI0/XI0_37/d__0_ XI11_5/XI0/XI0_37/d_0_ DECAP_INV_G11
XG5280 XI11_5/XI0/XI0_37/d_15_ XI11_5/XI0/XI0_37/d__15_ DECAP_INV_G11
XG5281 XI11_5/XI0/XI0_37/d_14_ XI11_5/XI0/XI0_37/d__14_ DECAP_INV_G11
XG5282 XI11_5/XI0/XI0_37/d_13_ XI11_5/XI0/XI0_37/d__13_ DECAP_INV_G11
XG5283 XI11_5/XI0/XI0_37/d_12_ XI11_5/XI0/XI0_37/d__12_ DECAP_INV_G11
XG5284 XI11_5/XI0/XI0_37/d_11_ XI11_5/XI0/XI0_37/d__11_ DECAP_INV_G11
XG5285 XI11_5/XI0/XI0_37/d_10_ XI11_5/XI0/XI0_37/d__10_ DECAP_INV_G11
XG5286 XI11_5/XI0/XI0_37/d_9_ XI11_5/XI0/XI0_37/d__9_ DECAP_INV_G11
XG5287 XI11_5/XI0/XI0_37/d_8_ XI11_5/XI0/XI0_37/d__8_ DECAP_INV_G11
XG5288 XI11_5/XI0/XI0_37/d_7_ XI11_5/XI0/XI0_37/d__7_ DECAP_INV_G11
XG5289 XI11_5/XI0/XI0_37/d_6_ XI11_5/XI0/XI0_37/d__6_ DECAP_INV_G11
XG5290 XI11_5/XI0/XI0_37/d_5_ XI11_5/XI0/XI0_37/d__5_ DECAP_INV_G11
XG5291 XI11_5/XI0/XI0_37/d_4_ XI11_5/XI0/XI0_37/d__4_ DECAP_INV_G11
XG5292 XI11_5/XI0/XI0_37/d_3_ XI11_5/XI0/XI0_37/d__3_ DECAP_INV_G11
XG5293 XI11_5/XI0/XI0_37/d_2_ XI11_5/XI0/XI0_37/d__2_ DECAP_INV_G11
XG5294 XI11_5/XI0/XI0_37/d_1_ XI11_5/XI0/XI0_37/d__1_ DECAP_INV_G11
XG5295 XI11_5/XI0/XI0_37/d_0_ XI11_5/XI0/XI0_37/d__0_ DECAP_INV_G11
XG5296 XI11_5/XI0/XI0_36/d__15_ XI11_5/XI0/XI0_36/d_15_ DECAP_INV_G11
XG5297 XI11_5/XI0/XI0_36/d__14_ XI11_5/XI0/XI0_36/d_14_ DECAP_INV_G11
XG5298 XI11_5/XI0/XI0_36/d__13_ XI11_5/XI0/XI0_36/d_13_ DECAP_INV_G11
XG5299 XI11_5/XI0/XI0_36/d__12_ XI11_5/XI0/XI0_36/d_12_ DECAP_INV_G11
XG5300 XI11_5/XI0/XI0_36/d__11_ XI11_5/XI0/XI0_36/d_11_ DECAP_INV_G11
XG5301 XI11_5/XI0/XI0_36/d__10_ XI11_5/XI0/XI0_36/d_10_ DECAP_INV_G11
XG5302 XI11_5/XI0/XI0_36/d__9_ XI11_5/XI0/XI0_36/d_9_ DECAP_INV_G11
XG5303 XI11_5/XI0/XI0_36/d__8_ XI11_5/XI0/XI0_36/d_8_ DECAP_INV_G11
XG5304 XI11_5/XI0/XI0_36/d__7_ XI11_5/XI0/XI0_36/d_7_ DECAP_INV_G11
XG5305 XI11_5/XI0/XI0_36/d__6_ XI11_5/XI0/XI0_36/d_6_ DECAP_INV_G11
XG5306 XI11_5/XI0/XI0_36/d__5_ XI11_5/XI0/XI0_36/d_5_ DECAP_INV_G11
XG5307 XI11_5/XI0/XI0_36/d__4_ XI11_5/XI0/XI0_36/d_4_ DECAP_INV_G11
XG5308 XI11_5/XI0/XI0_36/d__3_ XI11_5/XI0/XI0_36/d_3_ DECAP_INV_G11
XG5309 XI11_5/XI0/XI0_36/d__2_ XI11_5/XI0/XI0_36/d_2_ DECAP_INV_G11
XG5310 XI11_5/XI0/XI0_36/d__1_ XI11_5/XI0/XI0_36/d_1_ DECAP_INV_G11
XG5311 XI11_5/XI0/XI0_36/d__0_ XI11_5/XI0/XI0_36/d_0_ DECAP_INV_G11
XG5312 XI11_5/XI0/XI0_36/d_15_ XI11_5/XI0/XI0_36/d__15_ DECAP_INV_G11
XG5313 XI11_5/XI0/XI0_36/d_14_ XI11_5/XI0/XI0_36/d__14_ DECAP_INV_G11
XG5314 XI11_5/XI0/XI0_36/d_13_ XI11_5/XI0/XI0_36/d__13_ DECAP_INV_G11
XG5315 XI11_5/XI0/XI0_36/d_12_ XI11_5/XI0/XI0_36/d__12_ DECAP_INV_G11
XG5316 XI11_5/XI0/XI0_36/d_11_ XI11_5/XI0/XI0_36/d__11_ DECAP_INV_G11
XG5317 XI11_5/XI0/XI0_36/d_10_ XI11_5/XI0/XI0_36/d__10_ DECAP_INV_G11
XG5318 XI11_5/XI0/XI0_36/d_9_ XI11_5/XI0/XI0_36/d__9_ DECAP_INV_G11
XG5319 XI11_5/XI0/XI0_36/d_8_ XI11_5/XI0/XI0_36/d__8_ DECAP_INV_G11
XG5320 XI11_5/XI0/XI0_36/d_7_ XI11_5/XI0/XI0_36/d__7_ DECAP_INV_G11
XG5321 XI11_5/XI0/XI0_36/d_6_ XI11_5/XI0/XI0_36/d__6_ DECAP_INV_G11
XG5322 XI11_5/XI0/XI0_36/d_5_ XI11_5/XI0/XI0_36/d__5_ DECAP_INV_G11
XG5323 XI11_5/XI0/XI0_36/d_4_ XI11_5/XI0/XI0_36/d__4_ DECAP_INV_G11
XG5324 XI11_5/XI0/XI0_36/d_3_ XI11_5/XI0/XI0_36/d__3_ DECAP_INV_G11
XG5325 XI11_5/XI0/XI0_36/d_2_ XI11_5/XI0/XI0_36/d__2_ DECAP_INV_G11
XG5326 XI11_5/XI0/XI0_36/d_1_ XI11_5/XI0/XI0_36/d__1_ DECAP_INV_G11
XG5327 XI11_5/XI0/XI0_36/d_0_ XI11_5/XI0/XI0_36/d__0_ DECAP_INV_G11
XG5328 XI11_5/XI0/XI0_35/d__15_ XI11_5/XI0/XI0_35/d_15_ DECAP_INV_G11
XG5329 XI11_5/XI0/XI0_35/d__14_ XI11_5/XI0/XI0_35/d_14_ DECAP_INV_G11
XG5330 XI11_5/XI0/XI0_35/d__13_ XI11_5/XI0/XI0_35/d_13_ DECAP_INV_G11
XG5331 XI11_5/XI0/XI0_35/d__12_ XI11_5/XI0/XI0_35/d_12_ DECAP_INV_G11
XG5332 XI11_5/XI0/XI0_35/d__11_ XI11_5/XI0/XI0_35/d_11_ DECAP_INV_G11
XG5333 XI11_5/XI0/XI0_35/d__10_ XI11_5/XI0/XI0_35/d_10_ DECAP_INV_G11
XG5334 XI11_5/XI0/XI0_35/d__9_ XI11_5/XI0/XI0_35/d_9_ DECAP_INV_G11
XG5335 XI11_5/XI0/XI0_35/d__8_ XI11_5/XI0/XI0_35/d_8_ DECAP_INV_G11
XG5336 XI11_5/XI0/XI0_35/d__7_ XI11_5/XI0/XI0_35/d_7_ DECAP_INV_G11
XG5337 XI11_5/XI0/XI0_35/d__6_ XI11_5/XI0/XI0_35/d_6_ DECAP_INV_G11
XG5338 XI11_5/XI0/XI0_35/d__5_ XI11_5/XI0/XI0_35/d_5_ DECAP_INV_G11
XG5339 XI11_5/XI0/XI0_35/d__4_ XI11_5/XI0/XI0_35/d_4_ DECAP_INV_G11
XG5340 XI11_5/XI0/XI0_35/d__3_ XI11_5/XI0/XI0_35/d_3_ DECAP_INV_G11
XG5341 XI11_5/XI0/XI0_35/d__2_ XI11_5/XI0/XI0_35/d_2_ DECAP_INV_G11
XG5342 XI11_5/XI0/XI0_35/d__1_ XI11_5/XI0/XI0_35/d_1_ DECAP_INV_G11
XG5343 XI11_5/XI0/XI0_35/d__0_ XI11_5/XI0/XI0_35/d_0_ DECAP_INV_G11
XG5344 XI11_5/XI0/XI0_35/d_15_ XI11_5/XI0/XI0_35/d__15_ DECAP_INV_G11
XG5345 XI11_5/XI0/XI0_35/d_14_ XI11_5/XI0/XI0_35/d__14_ DECAP_INV_G11
XG5346 XI11_5/XI0/XI0_35/d_13_ XI11_5/XI0/XI0_35/d__13_ DECAP_INV_G11
XG5347 XI11_5/XI0/XI0_35/d_12_ XI11_5/XI0/XI0_35/d__12_ DECAP_INV_G11
XG5348 XI11_5/XI0/XI0_35/d_11_ XI11_5/XI0/XI0_35/d__11_ DECAP_INV_G11
XG5349 XI11_5/XI0/XI0_35/d_10_ XI11_5/XI0/XI0_35/d__10_ DECAP_INV_G11
XG5350 XI11_5/XI0/XI0_35/d_9_ XI11_5/XI0/XI0_35/d__9_ DECAP_INV_G11
XG5351 XI11_5/XI0/XI0_35/d_8_ XI11_5/XI0/XI0_35/d__8_ DECAP_INV_G11
XG5352 XI11_5/XI0/XI0_35/d_7_ XI11_5/XI0/XI0_35/d__7_ DECAP_INV_G11
XG5353 XI11_5/XI0/XI0_35/d_6_ XI11_5/XI0/XI0_35/d__6_ DECAP_INV_G11
XG5354 XI11_5/XI0/XI0_35/d_5_ XI11_5/XI0/XI0_35/d__5_ DECAP_INV_G11
XG5355 XI11_5/XI0/XI0_35/d_4_ XI11_5/XI0/XI0_35/d__4_ DECAP_INV_G11
XG5356 XI11_5/XI0/XI0_35/d_3_ XI11_5/XI0/XI0_35/d__3_ DECAP_INV_G11
XG5357 XI11_5/XI0/XI0_35/d_2_ XI11_5/XI0/XI0_35/d__2_ DECAP_INV_G11
XG5358 XI11_5/XI0/XI0_35/d_1_ XI11_5/XI0/XI0_35/d__1_ DECAP_INV_G11
XG5359 XI11_5/XI0/XI0_35/d_0_ XI11_5/XI0/XI0_35/d__0_ DECAP_INV_G11
XG5360 XI11_5/XI0/XI0_34/d__15_ XI11_5/XI0/XI0_34/d_15_ DECAP_INV_G11
XG5361 XI11_5/XI0/XI0_34/d__14_ XI11_5/XI0/XI0_34/d_14_ DECAP_INV_G11
XG5362 XI11_5/XI0/XI0_34/d__13_ XI11_5/XI0/XI0_34/d_13_ DECAP_INV_G11
XG5363 XI11_5/XI0/XI0_34/d__12_ XI11_5/XI0/XI0_34/d_12_ DECAP_INV_G11
XG5364 XI11_5/XI0/XI0_34/d__11_ XI11_5/XI0/XI0_34/d_11_ DECAP_INV_G11
XG5365 XI11_5/XI0/XI0_34/d__10_ XI11_5/XI0/XI0_34/d_10_ DECAP_INV_G11
XG5366 XI11_5/XI0/XI0_34/d__9_ XI11_5/XI0/XI0_34/d_9_ DECAP_INV_G11
XG5367 XI11_5/XI0/XI0_34/d__8_ XI11_5/XI0/XI0_34/d_8_ DECAP_INV_G11
XG5368 XI11_5/XI0/XI0_34/d__7_ XI11_5/XI0/XI0_34/d_7_ DECAP_INV_G11
XG5369 XI11_5/XI0/XI0_34/d__6_ XI11_5/XI0/XI0_34/d_6_ DECAP_INV_G11
XG5370 XI11_5/XI0/XI0_34/d__5_ XI11_5/XI0/XI0_34/d_5_ DECAP_INV_G11
XG5371 XI11_5/XI0/XI0_34/d__4_ XI11_5/XI0/XI0_34/d_4_ DECAP_INV_G11
XG5372 XI11_5/XI0/XI0_34/d__3_ XI11_5/XI0/XI0_34/d_3_ DECAP_INV_G11
XG5373 XI11_5/XI0/XI0_34/d__2_ XI11_5/XI0/XI0_34/d_2_ DECAP_INV_G11
XG5374 XI11_5/XI0/XI0_34/d__1_ XI11_5/XI0/XI0_34/d_1_ DECAP_INV_G11
XG5375 XI11_5/XI0/XI0_34/d__0_ XI11_5/XI0/XI0_34/d_0_ DECAP_INV_G11
XG5376 XI11_5/XI0/XI0_34/d_15_ XI11_5/XI0/XI0_34/d__15_ DECAP_INV_G11
XG5377 XI11_5/XI0/XI0_34/d_14_ XI11_5/XI0/XI0_34/d__14_ DECAP_INV_G11
XG5378 XI11_5/XI0/XI0_34/d_13_ XI11_5/XI0/XI0_34/d__13_ DECAP_INV_G11
XG5379 XI11_5/XI0/XI0_34/d_12_ XI11_5/XI0/XI0_34/d__12_ DECAP_INV_G11
XG5380 XI11_5/XI0/XI0_34/d_11_ XI11_5/XI0/XI0_34/d__11_ DECAP_INV_G11
XG5381 XI11_5/XI0/XI0_34/d_10_ XI11_5/XI0/XI0_34/d__10_ DECAP_INV_G11
XG5382 XI11_5/XI0/XI0_34/d_9_ XI11_5/XI0/XI0_34/d__9_ DECAP_INV_G11
XG5383 XI11_5/XI0/XI0_34/d_8_ XI11_5/XI0/XI0_34/d__8_ DECAP_INV_G11
XG5384 XI11_5/XI0/XI0_34/d_7_ XI11_5/XI0/XI0_34/d__7_ DECAP_INV_G11
XG5385 XI11_5/XI0/XI0_34/d_6_ XI11_5/XI0/XI0_34/d__6_ DECAP_INV_G11
XG5386 XI11_5/XI0/XI0_34/d_5_ XI11_5/XI0/XI0_34/d__5_ DECAP_INV_G11
XG5387 XI11_5/XI0/XI0_34/d_4_ XI11_5/XI0/XI0_34/d__4_ DECAP_INV_G11
XG5388 XI11_5/XI0/XI0_34/d_3_ XI11_5/XI0/XI0_34/d__3_ DECAP_INV_G11
XG5389 XI11_5/XI0/XI0_34/d_2_ XI11_5/XI0/XI0_34/d__2_ DECAP_INV_G11
XG5390 XI11_5/XI0/XI0_34/d_1_ XI11_5/XI0/XI0_34/d__1_ DECAP_INV_G11
XG5391 XI11_5/XI0/XI0_34/d_0_ XI11_5/XI0/XI0_34/d__0_ DECAP_INV_G11
XG5392 XI11_5/XI0/XI0_33/d__15_ XI11_5/XI0/XI0_33/d_15_ DECAP_INV_G11
XG5393 XI11_5/XI0/XI0_33/d__14_ XI11_5/XI0/XI0_33/d_14_ DECAP_INV_G11
XG5394 XI11_5/XI0/XI0_33/d__13_ XI11_5/XI0/XI0_33/d_13_ DECAP_INV_G11
XG5395 XI11_5/XI0/XI0_33/d__12_ XI11_5/XI0/XI0_33/d_12_ DECAP_INV_G11
XG5396 XI11_5/XI0/XI0_33/d__11_ XI11_5/XI0/XI0_33/d_11_ DECAP_INV_G11
XG5397 XI11_5/XI0/XI0_33/d__10_ XI11_5/XI0/XI0_33/d_10_ DECAP_INV_G11
XG5398 XI11_5/XI0/XI0_33/d__9_ XI11_5/XI0/XI0_33/d_9_ DECAP_INV_G11
XG5399 XI11_5/XI0/XI0_33/d__8_ XI11_5/XI0/XI0_33/d_8_ DECAP_INV_G11
XG5400 XI11_5/XI0/XI0_33/d__7_ XI11_5/XI0/XI0_33/d_7_ DECAP_INV_G11
XG5401 XI11_5/XI0/XI0_33/d__6_ XI11_5/XI0/XI0_33/d_6_ DECAP_INV_G11
XG5402 XI11_5/XI0/XI0_33/d__5_ XI11_5/XI0/XI0_33/d_5_ DECAP_INV_G11
XG5403 XI11_5/XI0/XI0_33/d__4_ XI11_5/XI0/XI0_33/d_4_ DECAP_INV_G11
XG5404 XI11_5/XI0/XI0_33/d__3_ XI11_5/XI0/XI0_33/d_3_ DECAP_INV_G11
XG5405 XI11_5/XI0/XI0_33/d__2_ XI11_5/XI0/XI0_33/d_2_ DECAP_INV_G11
XG5406 XI11_5/XI0/XI0_33/d__1_ XI11_5/XI0/XI0_33/d_1_ DECAP_INV_G11
XG5407 XI11_5/XI0/XI0_33/d__0_ XI11_5/XI0/XI0_33/d_0_ DECAP_INV_G11
XG5408 XI11_5/XI0/XI0_33/d_15_ XI11_5/XI0/XI0_33/d__15_ DECAP_INV_G11
XG5409 XI11_5/XI0/XI0_33/d_14_ XI11_5/XI0/XI0_33/d__14_ DECAP_INV_G11
XG5410 XI11_5/XI0/XI0_33/d_13_ XI11_5/XI0/XI0_33/d__13_ DECAP_INV_G11
XG5411 XI11_5/XI0/XI0_33/d_12_ XI11_5/XI0/XI0_33/d__12_ DECAP_INV_G11
XG5412 XI11_5/XI0/XI0_33/d_11_ XI11_5/XI0/XI0_33/d__11_ DECAP_INV_G11
XG5413 XI11_5/XI0/XI0_33/d_10_ XI11_5/XI0/XI0_33/d__10_ DECAP_INV_G11
XG5414 XI11_5/XI0/XI0_33/d_9_ XI11_5/XI0/XI0_33/d__9_ DECAP_INV_G11
XG5415 XI11_5/XI0/XI0_33/d_8_ XI11_5/XI0/XI0_33/d__8_ DECAP_INV_G11
XG5416 XI11_5/XI0/XI0_33/d_7_ XI11_5/XI0/XI0_33/d__7_ DECAP_INV_G11
XG5417 XI11_5/XI0/XI0_33/d_6_ XI11_5/XI0/XI0_33/d__6_ DECAP_INV_G11
XG5418 XI11_5/XI0/XI0_33/d_5_ XI11_5/XI0/XI0_33/d__5_ DECAP_INV_G11
XG5419 XI11_5/XI0/XI0_33/d_4_ XI11_5/XI0/XI0_33/d__4_ DECAP_INV_G11
XG5420 XI11_5/XI0/XI0_33/d_3_ XI11_5/XI0/XI0_33/d__3_ DECAP_INV_G11
XG5421 XI11_5/XI0/XI0_33/d_2_ XI11_5/XI0/XI0_33/d__2_ DECAP_INV_G11
XG5422 XI11_5/XI0/XI0_33/d_1_ XI11_5/XI0/XI0_33/d__1_ DECAP_INV_G11
XG5423 XI11_5/XI0/XI0_33/d_0_ XI11_5/XI0/XI0_33/d__0_ DECAP_INV_G11
XG5424 XI11_5/XI0/XI0_32/d__15_ XI11_5/XI0/XI0_32/d_15_ DECAP_INV_G11
XG5425 XI11_5/XI0/XI0_32/d__14_ XI11_5/XI0/XI0_32/d_14_ DECAP_INV_G11
XG5426 XI11_5/XI0/XI0_32/d__13_ XI11_5/XI0/XI0_32/d_13_ DECAP_INV_G11
XG5427 XI11_5/XI0/XI0_32/d__12_ XI11_5/XI0/XI0_32/d_12_ DECAP_INV_G11
XG5428 XI11_5/XI0/XI0_32/d__11_ XI11_5/XI0/XI0_32/d_11_ DECAP_INV_G11
XG5429 XI11_5/XI0/XI0_32/d__10_ XI11_5/XI0/XI0_32/d_10_ DECAP_INV_G11
XG5430 XI11_5/XI0/XI0_32/d__9_ XI11_5/XI0/XI0_32/d_9_ DECAP_INV_G11
XG5431 XI11_5/XI0/XI0_32/d__8_ XI11_5/XI0/XI0_32/d_8_ DECAP_INV_G11
XG5432 XI11_5/XI0/XI0_32/d__7_ XI11_5/XI0/XI0_32/d_7_ DECAP_INV_G11
XG5433 XI11_5/XI0/XI0_32/d__6_ XI11_5/XI0/XI0_32/d_6_ DECAP_INV_G11
XG5434 XI11_5/XI0/XI0_32/d__5_ XI11_5/XI0/XI0_32/d_5_ DECAP_INV_G11
XG5435 XI11_5/XI0/XI0_32/d__4_ XI11_5/XI0/XI0_32/d_4_ DECAP_INV_G11
XG5436 XI11_5/XI0/XI0_32/d__3_ XI11_5/XI0/XI0_32/d_3_ DECAP_INV_G11
XG5437 XI11_5/XI0/XI0_32/d__2_ XI11_5/XI0/XI0_32/d_2_ DECAP_INV_G11
XG5438 XI11_5/XI0/XI0_32/d__1_ XI11_5/XI0/XI0_32/d_1_ DECAP_INV_G11
XG5439 XI11_5/XI0/XI0_32/d__0_ XI11_5/XI0/XI0_32/d_0_ DECAP_INV_G11
XG5440 XI11_5/XI0/XI0_32/d_15_ XI11_5/XI0/XI0_32/d__15_ DECAP_INV_G11
XG5441 XI11_5/XI0/XI0_32/d_14_ XI11_5/XI0/XI0_32/d__14_ DECAP_INV_G11
XG5442 XI11_5/XI0/XI0_32/d_13_ XI11_5/XI0/XI0_32/d__13_ DECAP_INV_G11
XG5443 XI11_5/XI0/XI0_32/d_12_ XI11_5/XI0/XI0_32/d__12_ DECAP_INV_G11
XG5444 XI11_5/XI0/XI0_32/d_11_ XI11_5/XI0/XI0_32/d__11_ DECAP_INV_G11
XG5445 XI11_5/XI0/XI0_32/d_10_ XI11_5/XI0/XI0_32/d__10_ DECAP_INV_G11
XG5446 XI11_5/XI0/XI0_32/d_9_ XI11_5/XI0/XI0_32/d__9_ DECAP_INV_G11
XG5447 XI11_5/XI0/XI0_32/d_8_ XI11_5/XI0/XI0_32/d__8_ DECAP_INV_G11
XG5448 XI11_5/XI0/XI0_32/d_7_ XI11_5/XI0/XI0_32/d__7_ DECAP_INV_G11
XG5449 XI11_5/XI0/XI0_32/d_6_ XI11_5/XI0/XI0_32/d__6_ DECAP_INV_G11
XG5450 XI11_5/XI0/XI0_32/d_5_ XI11_5/XI0/XI0_32/d__5_ DECAP_INV_G11
XG5451 XI11_5/XI0/XI0_32/d_4_ XI11_5/XI0/XI0_32/d__4_ DECAP_INV_G11
XG5452 XI11_5/XI0/XI0_32/d_3_ XI11_5/XI0/XI0_32/d__3_ DECAP_INV_G11
XG5453 XI11_5/XI0/XI0_32/d_2_ XI11_5/XI0/XI0_32/d__2_ DECAP_INV_G11
XG5454 XI11_5/XI0/XI0_32/d_1_ XI11_5/XI0/XI0_32/d__1_ DECAP_INV_G11
XG5455 XI11_5/XI0/XI0_32/d_0_ XI11_5/XI0/XI0_32/d__0_ DECAP_INV_G11
XG5456 XI11_5/XI0/XI0_31/d__15_ XI11_5/XI0/XI0_31/d_15_ DECAP_INV_G11
XG5457 XI11_5/XI0/XI0_31/d__14_ XI11_5/XI0/XI0_31/d_14_ DECAP_INV_G11
XG5458 XI11_5/XI0/XI0_31/d__13_ XI11_5/XI0/XI0_31/d_13_ DECAP_INV_G11
XG5459 XI11_5/XI0/XI0_31/d__12_ XI11_5/XI0/XI0_31/d_12_ DECAP_INV_G11
XG5460 XI11_5/XI0/XI0_31/d__11_ XI11_5/XI0/XI0_31/d_11_ DECAP_INV_G11
XG5461 XI11_5/XI0/XI0_31/d__10_ XI11_5/XI0/XI0_31/d_10_ DECAP_INV_G11
XG5462 XI11_5/XI0/XI0_31/d__9_ XI11_5/XI0/XI0_31/d_9_ DECAP_INV_G11
XG5463 XI11_5/XI0/XI0_31/d__8_ XI11_5/XI0/XI0_31/d_8_ DECAP_INV_G11
XG5464 XI11_5/XI0/XI0_31/d__7_ XI11_5/XI0/XI0_31/d_7_ DECAP_INV_G11
XG5465 XI11_5/XI0/XI0_31/d__6_ XI11_5/XI0/XI0_31/d_6_ DECAP_INV_G11
XG5466 XI11_5/XI0/XI0_31/d__5_ XI11_5/XI0/XI0_31/d_5_ DECAP_INV_G11
XG5467 XI11_5/XI0/XI0_31/d__4_ XI11_5/XI0/XI0_31/d_4_ DECAP_INV_G11
XG5468 XI11_5/XI0/XI0_31/d__3_ XI11_5/XI0/XI0_31/d_3_ DECAP_INV_G11
XG5469 XI11_5/XI0/XI0_31/d__2_ XI11_5/XI0/XI0_31/d_2_ DECAP_INV_G11
XG5470 XI11_5/XI0/XI0_31/d__1_ XI11_5/XI0/XI0_31/d_1_ DECAP_INV_G11
XG5471 XI11_5/XI0/XI0_31/d__0_ XI11_5/XI0/XI0_31/d_0_ DECAP_INV_G11
XG5472 XI11_5/XI0/XI0_31/d_15_ XI11_5/XI0/XI0_31/d__15_ DECAP_INV_G11
XG5473 XI11_5/XI0/XI0_31/d_14_ XI11_5/XI0/XI0_31/d__14_ DECAP_INV_G11
XG5474 XI11_5/XI0/XI0_31/d_13_ XI11_5/XI0/XI0_31/d__13_ DECAP_INV_G11
XG5475 XI11_5/XI0/XI0_31/d_12_ XI11_5/XI0/XI0_31/d__12_ DECAP_INV_G11
XG5476 XI11_5/XI0/XI0_31/d_11_ XI11_5/XI0/XI0_31/d__11_ DECAP_INV_G11
XG5477 XI11_5/XI0/XI0_31/d_10_ XI11_5/XI0/XI0_31/d__10_ DECAP_INV_G11
XG5478 XI11_5/XI0/XI0_31/d_9_ XI11_5/XI0/XI0_31/d__9_ DECAP_INV_G11
XG5479 XI11_5/XI0/XI0_31/d_8_ XI11_5/XI0/XI0_31/d__8_ DECAP_INV_G11
XG5480 XI11_5/XI0/XI0_31/d_7_ XI11_5/XI0/XI0_31/d__7_ DECAP_INV_G11
XG5481 XI11_5/XI0/XI0_31/d_6_ XI11_5/XI0/XI0_31/d__6_ DECAP_INV_G11
XG5482 XI11_5/XI0/XI0_31/d_5_ XI11_5/XI0/XI0_31/d__5_ DECAP_INV_G11
XG5483 XI11_5/XI0/XI0_31/d_4_ XI11_5/XI0/XI0_31/d__4_ DECAP_INV_G11
XG5484 XI11_5/XI0/XI0_31/d_3_ XI11_5/XI0/XI0_31/d__3_ DECAP_INV_G11
XG5485 XI11_5/XI0/XI0_31/d_2_ XI11_5/XI0/XI0_31/d__2_ DECAP_INV_G11
XG5486 XI11_5/XI0/XI0_31/d_1_ XI11_5/XI0/XI0_31/d__1_ DECAP_INV_G11
XG5487 XI11_5/XI0/XI0_31/d_0_ XI11_5/XI0/XI0_31/d__0_ DECAP_INV_G11
XG5488 XI11_5/XI0/XI0_30/d__15_ XI11_5/XI0/XI0_30/d_15_ DECAP_INV_G11
XG5489 XI11_5/XI0/XI0_30/d__14_ XI11_5/XI0/XI0_30/d_14_ DECAP_INV_G11
XG5490 XI11_5/XI0/XI0_30/d__13_ XI11_5/XI0/XI0_30/d_13_ DECAP_INV_G11
XG5491 XI11_5/XI0/XI0_30/d__12_ XI11_5/XI0/XI0_30/d_12_ DECAP_INV_G11
XG5492 XI11_5/XI0/XI0_30/d__11_ XI11_5/XI0/XI0_30/d_11_ DECAP_INV_G11
XG5493 XI11_5/XI0/XI0_30/d__10_ XI11_5/XI0/XI0_30/d_10_ DECAP_INV_G11
XG5494 XI11_5/XI0/XI0_30/d__9_ XI11_5/XI0/XI0_30/d_9_ DECAP_INV_G11
XG5495 XI11_5/XI0/XI0_30/d__8_ XI11_5/XI0/XI0_30/d_8_ DECAP_INV_G11
XG5496 XI11_5/XI0/XI0_30/d__7_ XI11_5/XI0/XI0_30/d_7_ DECAP_INV_G11
XG5497 XI11_5/XI0/XI0_30/d__6_ XI11_5/XI0/XI0_30/d_6_ DECAP_INV_G11
XG5498 XI11_5/XI0/XI0_30/d__5_ XI11_5/XI0/XI0_30/d_5_ DECAP_INV_G11
XG5499 XI11_5/XI0/XI0_30/d__4_ XI11_5/XI0/XI0_30/d_4_ DECAP_INV_G11
XG5500 XI11_5/XI0/XI0_30/d__3_ XI11_5/XI0/XI0_30/d_3_ DECAP_INV_G11
XG5501 XI11_5/XI0/XI0_30/d__2_ XI11_5/XI0/XI0_30/d_2_ DECAP_INV_G11
XG5502 XI11_5/XI0/XI0_30/d__1_ XI11_5/XI0/XI0_30/d_1_ DECAP_INV_G11
XG5503 XI11_5/XI0/XI0_30/d__0_ XI11_5/XI0/XI0_30/d_0_ DECAP_INV_G11
XG5504 XI11_5/XI0/XI0_30/d_15_ XI11_5/XI0/XI0_30/d__15_ DECAP_INV_G11
XG5505 XI11_5/XI0/XI0_30/d_14_ XI11_5/XI0/XI0_30/d__14_ DECAP_INV_G11
XG5506 XI11_5/XI0/XI0_30/d_13_ XI11_5/XI0/XI0_30/d__13_ DECAP_INV_G11
XG5507 XI11_5/XI0/XI0_30/d_12_ XI11_5/XI0/XI0_30/d__12_ DECAP_INV_G11
XG5508 XI11_5/XI0/XI0_30/d_11_ XI11_5/XI0/XI0_30/d__11_ DECAP_INV_G11
XG5509 XI11_5/XI0/XI0_30/d_10_ XI11_5/XI0/XI0_30/d__10_ DECAP_INV_G11
XG5510 XI11_5/XI0/XI0_30/d_9_ XI11_5/XI0/XI0_30/d__9_ DECAP_INV_G11
XG5511 XI11_5/XI0/XI0_30/d_8_ XI11_5/XI0/XI0_30/d__8_ DECAP_INV_G11
XG5512 XI11_5/XI0/XI0_30/d_7_ XI11_5/XI0/XI0_30/d__7_ DECAP_INV_G11
XG5513 XI11_5/XI0/XI0_30/d_6_ XI11_5/XI0/XI0_30/d__6_ DECAP_INV_G11
XG5514 XI11_5/XI0/XI0_30/d_5_ XI11_5/XI0/XI0_30/d__5_ DECAP_INV_G11
XG5515 XI11_5/XI0/XI0_30/d_4_ XI11_5/XI0/XI0_30/d__4_ DECAP_INV_G11
XG5516 XI11_5/XI0/XI0_30/d_3_ XI11_5/XI0/XI0_30/d__3_ DECAP_INV_G11
XG5517 XI11_5/XI0/XI0_30/d_2_ XI11_5/XI0/XI0_30/d__2_ DECAP_INV_G11
XG5518 XI11_5/XI0/XI0_30/d_1_ XI11_5/XI0/XI0_30/d__1_ DECAP_INV_G11
XG5519 XI11_5/XI0/XI0_30/d_0_ XI11_5/XI0/XI0_30/d__0_ DECAP_INV_G11
XG5520 XI11_5/XI0/XI0_29/d__15_ XI11_5/XI0/XI0_29/d_15_ DECAP_INV_G11
XG5521 XI11_5/XI0/XI0_29/d__14_ XI11_5/XI0/XI0_29/d_14_ DECAP_INV_G11
XG5522 XI11_5/XI0/XI0_29/d__13_ XI11_5/XI0/XI0_29/d_13_ DECAP_INV_G11
XG5523 XI11_5/XI0/XI0_29/d__12_ XI11_5/XI0/XI0_29/d_12_ DECAP_INV_G11
XG5524 XI11_5/XI0/XI0_29/d__11_ XI11_5/XI0/XI0_29/d_11_ DECAP_INV_G11
XG5525 XI11_5/XI0/XI0_29/d__10_ XI11_5/XI0/XI0_29/d_10_ DECAP_INV_G11
XG5526 XI11_5/XI0/XI0_29/d__9_ XI11_5/XI0/XI0_29/d_9_ DECAP_INV_G11
XG5527 XI11_5/XI0/XI0_29/d__8_ XI11_5/XI0/XI0_29/d_8_ DECAP_INV_G11
XG5528 XI11_5/XI0/XI0_29/d__7_ XI11_5/XI0/XI0_29/d_7_ DECAP_INV_G11
XG5529 XI11_5/XI0/XI0_29/d__6_ XI11_5/XI0/XI0_29/d_6_ DECAP_INV_G11
XG5530 XI11_5/XI0/XI0_29/d__5_ XI11_5/XI0/XI0_29/d_5_ DECAP_INV_G11
XG5531 XI11_5/XI0/XI0_29/d__4_ XI11_5/XI0/XI0_29/d_4_ DECAP_INV_G11
XG5532 XI11_5/XI0/XI0_29/d__3_ XI11_5/XI0/XI0_29/d_3_ DECAP_INV_G11
XG5533 XI11_5/XI0/XI0_29/d__2_ XI11_5/XI0/XI0_29/d_2_ DECAP_INV_G11
XG5534 XI11_5/XI0/XI0_29/d__1_ XI11_5/XI0/XI0_29/d_1_ DECAP_INV_G11
XG5535 XI11_5/XI0/XI0_29/d__0_ XI11_5/XI0/XI0_29/d_0_ DECAP_INV_G11
XG5536 XI11_5/XI0/XI0_29/d_15_ XI11_5/XI0/XI0_29/d__15_ DECAP_INV_G11
XG5537 XI11_5/XI0/XI0_29/d_14_ XI11_5/XI0/XI0_29/d__14_ DECAP_INV_G11
XG5538 XI11_5/XI0/XI0_29/d_13_ XI11_5/XI0/XI0_29/d__13_ DECAP_INV_G11
XG5539 XI11_5/XI0/XI0_29/d_12_ XI11_5/XI0/XI0_29/d__12_ DECAP_INV_G11
XG5540 XI11_5/XI0/XI0_29/d_11_ XI11_5/XI0/XI0_29/d__11_ DECAP_INV_G11
XG5541 XI11_5/XI0/XI0_29/d_10_ XI11_5/XI0/XI0_29/d__10_ DECAP_INV_G11
XG5542 XI11_5/XI0/XI0_29/d_9_ XI11_5/XI0/XI0_29/d__9_ DECAP_INV_G11
XG5543 XI11_5/XI0/XI0_29/d_8_ XI11_5/XI0/XI0_29/d__8_ DECAP_INV_G11
XG5544 XI11_5/XI0/XI0_29/d_7_ XI11_5/XI0/XI0_29/d__7_ DECAP_INV_G11
XG5545 XI11_5/XI0/XI0_29/d_6_ XI11_5/XI0/XI0_29/d__6_ DECAP_INV_G11
XG5546 XI11_5/XI0/XI0_29/d_5_ XI11_5/XI0/XI0_29/d__5_ DECAP_INV_G11
XG5547 XI11_5/XI0/XI0_29/d_4_ XI11_5/XI0/XI0_29/d__4_ DECAP_INV_G11
XG5548 XI11_5/XI0/XI0_29/d_3_ XI11_5/XI0/XI0_29/d__3_ DECAP_INV_G11
XG5549 XI11_5/XI0/XI0_29/d_2_ XI11_5/XI0/XI0_29/d__2_ DECAP_INV_G11
XG5550 XI11_5/XI0/XI0_29/d_1_ XI11_5/XI0/XI0_29/d__1_ DECAP_INV_G11
XG5551 XI11_5/XI0/XI0_29/d_0_ XI11_5/XI0/XI0_29/d__0_ DECAP_INV_G11
XG5552 XI11_5/XI0/XI0_28/d__15_ XI11_5/XI0/XI0_28/d_15_ DECAP_INV_G11
XG5553 XI11_5/XI0/XI0_28/d__14_ XI11_5/XI0/XI0_28/d_14_ DECAP_INV_G11
XG5554 XI11_5/XI0/XI0_28/d__13_ XI11_5/XI0/XI0_28/d_13_ DECAP_INV_G11
XG5555 XI11_5/XI0/XI0_28/d__12_ XI11_5/XI0/XI0_28/d_12_ DECAP_INV_G11
XG5556 XI11_5/XI0/XI0_28/d__11_ XI11_5/XI0/XI0_28/d_11_ DECAP_INV_G11
XG5557 XI11_5/XI0/XI0_28/d__10_ XI11_5/XI0/XI0_28/d_10_ DECAP_INV_G11
XG5558 XI11_5/XI0/XI0_28/d__9_ XI11_5/XI0/XI0_28/d_9_ DECAP_INV_G11
XG5559 XI11_5/XI0/XI0_28/d__8_ XI11_5/XI0/XI0_28/d_8_ DECAP_INV_G11
XG5560 XI11_5/XI0/XI0_28/d__7_ XI11_5/XI0/XI0_28/d_7_ DECAP_INV_G11
XG5561 XI11_5/XI0/XI0_28/d__6_ XI11_5/XI0/XI0_28/d_6_ DECAP_INV_G11
XG5562 XI11_5/XI0/XI0_28/d__5_ XI11_5/XI0/XI0_28/d_5_ DECAP_INV_G11
XG5563 XI11_5/XI0/XI0_28/d__4_ XI11_5/XI0/XI0_28/d_4_ DECAP_INV_G11
XG5564 XI11_5/XI0/XI0_28/d__3_ XI11_5/XI0/XI0_28/d_3_ DECAP_INV_G11
XG5565 XI11_5/XI0/XI0_28/d__2_ XI11_5/XI0/XI0_28/d_2_ DECAP_INV_G11
XG5566 XI11_5/XI0/XI0_28/d__1_ XI11_5/XI0/XI0_28/d_1_ DECAP_INV_G11
XG5567 XI11_5/XI0/XI0_28/d__0_ XI11_5/XI0/XI0_28/d_0_ DECAP_INV_G11
XG5568 XI11_5/XI0/XI0_28/d_15_ XI11_5/XI0/XI0_28/d__15_ DECAP_INV_G11
XG5569 XI11_5/XI0/XI0_28/d_14_ XI11_5/XI0/XI0_28/d__14_ DECAP_INV_G11
XG5570 XI11_5/XI0/XI0_28/d_13_ XI11_5/XI0/XI0_28/d__13_ DECAP_INV_G11
XG5571 XI11_5/XI0/XI0_28/d_12_ XI11_5/XI0/XI0_28/d__12_ DECAP_INV_G11
XG5572 XI11_5/XI0/XI0_28/d_11_ XI11_5/XI0/XI0_28/d__11_ DECAP_INV_G11
XG5573 XI11_5/XI0/XI0_28/d_10_ XI11_5/XI0/XI0_28/d__10_ DECAP_INV_G11
XG5574 XI11_5/XI0/XI0_28/d_9_ XI11_5/XI0/XI0_28/d__9_ DECAP_INV_G11
XG5575 XI11_5/XI0/XI0_28/d_8_ XI11_5/XI0/XI0_28/d__8_ DECAP_INV_G11
XG5576 XI11_5/XI0/XI0_28/d_7_ XI11_5/XI0/XI0_28/d__7_ DECAP_INV_G11
XG5577 XI11_5/XI0/XI0_28/d_6_ XI11_5/XI0/XI0_28/d__6_ DECAP_INV_G11
XG5578 XI11_5/XI0/XI0_28/d_5_ XI11_5/XI0/XI0_28/d__5_ DECAP_INV_G11
XG5579 XI11_5/XI0/XI0_28/d_4_ XI11_5/XI0/XI0_28/d__4_ DECAP_INV_G11
XG5580 XI11_5/XI0/XI0_28/d_3_ XI11_5/XI0/XI0_28/d__3_ DECAP_INV_G11
XG5581 XI11_5/XI0/XI0_28/d_2_ XI11_5/XI0/XI0_28/d__2_ DECAP_INV_G11
XG5582 XI11_5/XI0/XI0_28/d_1_ XI11_5/XI0/XI0_28/d__1_ DECAP_INV_G11
XG5583 XI11_5/XI0/XI0_28/d_0_ XI11_5/XI0/XI0_28/d__0_ DECAP_INV_G11
XG5584 XI11_5/XI0/XI0_27/d__15_ XI11_5/XI0/XI0_27/d_15_ DECAP_INV_G11
XG5585 XI11_5/XI0/XI0_27/d__14_ XI11_5/XI0/XI0_27/d_14_ DECAP_INV_G11
XG5586 XI11_5/XI0/XI0_27/d__13_ XI11_5/XI0/XI0_27/d_13_ DECAP_INV_G11
XG5587 XI11_5/XI0/XI0_27/d__12_ XI11_5/XI0/XI0_27/d_12_ DECAP_INV_G11
XG5588 XI11_5/XI0/XI0_27/d__11_ XI11_5/XI0/XI0_27/d_11_ DECAP_INV_G11
XG5589 XI11_5/XI0/XI0_27/d__10_ XI11_5/XI0/XI0_27/d_10_ DECAP_INV_G11
XG5590 XI11_5/XI0/XI0_27/d__9_ XI11_5/XI0/XI0_27/d_9_ DECAP_INV_G11
XG5591 XI11_5/XI0/XI0_27/d__8_ XI11_5/XI0/XI0_27/d_8_ DECAP_INV_G11
XG5592 XI11_5/XI0/XI0_27/d__7_ XI11_5/XI0/XI0_27/d_7_ DECAP_INV_G11
XG5593 XI11_5/XI0/XI0_27/d__6_ XI11_5/XI0/XI0_27/d_6_ DECAP_INV_G11
XG5594 XI11_5/XI0/XI0_27/d__5_ XI11_5/XI0/XI0_27/d_5_ DECAP_INV_G11
XG5595 XI11_5/XI0/XI0_27/d__4_ XI11_5/XI0/XI0_27/d_4_ DECAP_INV_G11
XG5596 XI11_5/XI0/XI0_27/d__3_ XI11_5/XI0/XI0_27/d_3_ DECAP_INV_G11
XG5597 XI11_5/XI0/XI0_27/d__2_ XI11_5/XI0/XI0_27/d_2_ DECAP_INV_G11
XG5598 XI11_5/XI0/XI0_27/d__1_ XI11_5/XI0/XI0_27/d_1_ DECAP_INV_G11
XG5599 XI11_5/XI0/XI0_27/d__0_ XI11_5/XI0/XI0_27/d_0_ DECAP_INV_G11
XG5600 XI11_5/XI0/XI0_27/d_15_ XI11_5/XI0/XI0_27/d__15_ DECAP_INV_G11
XG5601 XI11_5/XI0/XI0_27/d_14_ XI11_5/XI0/XI0_27/d__14_ DECAP_INV_G11
XG5602 XI11_5/XI0/XI0_27/d_13_ XI11_5/XI0/XI0_27/d__13_ DECAP_INV_G11
XG5603 XI11_5/XI0/XI0_27/d_12_ XI11_5/XI0/XI0_27/d__12_ DECAP_INV_G11
XG5604 XI11_5/XI0/XI0_27/d_11_ XI11_5/XI0/XI0_27/d__11_ DECAP_INV_G11
XG5605 XI11_5/XI0/XI0_27/d_10_ XI11_5/XI0/XI0_27/d__10_ DECAP_INV_G11
XG5606 XI11_5/XI0/XI0_27/d_9_ XI11_5/XI0/XI0_27/d__9_ DECAP_INV_G11
XG5607 XI11_5/XI0/XI0_27/d_8_ XI11_5/XI0/XI0_27/d__8_ DECAP_INV_G11
XG5608 XI11_5/XI0/XI0_27/d_7_ XI11_5/XI0/XI0_27/d__7_ DECAP_INV_G11
XG5609 XI11_5/XI0/XI0_27/d_6_ XI11_5/XI0/XI0_27/d__6_ DECAP_INV_G11
XG5610 XI11_5/XI0/XI0_27/d_5_ XI11_5/XI0/XI0_27/d__5_ DECAP_INV_G11
XG5611 XI11_5/XI0/XI0_27/d_4_ XI11_5/XI0/XI0_27/d__4_ DECAP_INV_G11
XG5612 XI11_5/XI0/XI0_27/d_3_ XI11_5/XI0/XI0_27/d__3_ DECAP_INV_G11
XG5613 XI11_5/XI0/XI0_27/d_2_ XI11_5/XI0/XI0_27/d__2_ DECAP_INV_G11
XG5614 XI11_5/XI0/XI0_27/d_1_ XI11_5/XI0/XI0_27/d__1_ DECAP_INV_G11
XG5615 XI11_5/XI0/XI0_27/d_0_ XI11_5/XI0/XI0_27/d__0_ DECAP_INV_G11
XG5616 XI11_5/XI0/XI0_26/d__15_ XI11_5/XI0/XI0_26/d_15_ DECAP_INV_G11
XG5617 XI11_5/XI0/XI0_26/d__14_ XI11_5/XI0/XI0_26/d_14_ DECAP_INV_G11
XG5618 XI11_5/XI0/XI0_26/d__13_ XI11_5/XI0/XI0_26/d_13_ DECAP_INV_G11
XG5619 XI11_5/XI0/XI0_26/d__12_ XI11_5/XI0/XI0_26/d_12_ DECAP_INV_G11
XG5620 XI11_5/XI0/XI0_26/d__11_ XI11_5/XI0/XI0_26/d_11_ DECAP_INV_G11
XG5621 XI11_5/XI0/XI0_26/d__10_ XI11_5/XI0/XI0_26/d_10_ DECAP_INV_G11
XG5622 XI11_5/XI0/XI0_26/d__9_ XI11_5/XI0/XI0_26/d_9_ DECAP_INV_G11
XG5623 XI11_5/XI0/XI0_26/d__8_ XI11_5/XI0/XI0_26/d_8_ DECAP_INV_G11
XG5624 XI11_5/XI0/XI0_26/d__7_ XI11_5/XI0/XI0_26/d_7_ DECAP_INV_G11
XG5625 XI11_5/XI0/XI0_26/d__6_ XI11_5/XI0/XI0_26/d_6_ DECAP_INV_G11
XG5626 XI11_5/XI0/XI0_26/d__5_ XI11_5/XI0/XI0_26/d_5_ DECAP_INV_G11
XG5627 XI11_5/XI0/XI0_26/d__4_ XI11_5/XI0/XI0_26/d_4_ DECAP_INV_G11
XG5628 XI11_5/XI0/XI0_26/d__3_ XI11_5/XI0/XI0_26/d_3_ DECAP_INV_G11
XG5629 XI11_5/XI0/XI0_26/d__2_ XI11_5/XI0/XI0_26/d_2_ DECAP_INV_G11
XG5630 XI11_5/XI0/XI0_26/d__1_ XI11_5/XI0/XI0_26/d_1_ DECAP_INV_G11
XG5631 XI11_5/XI0/XI0_26/d__0_ XI11_5/XI0/XI0_26/d_0_ DECAP_INV_G11
XG5632 XI11_5/XI0/XI0_26/d_15_ XI11_5/XI0/XI0_26/d__15_ DECAP_INV_G11
XG5633 XI11_5/XI0/XI0_26/d_14_ XI11_5/XI0/XI0_26/d__14_ DECAP_INV_G11
XG5634 XI11_5/XI0/XI0_26/d_13_ XI11_5/XI0/XI0_26/d__13_ DECAP_INV_G11
XG5635 XI11_5/XI0/XI0_26/d_12_ XI11_5/XI0/XI0_26/d__12_ DECAP_INV_G11
XG5636 XI11_5/XI0/XI0_26/d_11_ XI11_5/XI0/XI0_26/d__11_ DECAP_INV_G11
XG5637 XI11_5/XI0/XI0_26/d_10_ XI11_5/XI0/XI0_26/d__10_ DECAP_INV_G11
XG5638 XI11_5/XI0/XI0_26/d_9_ XI11_5/XI0/XI0_26/d__9_ DECAP_INV_G11
XG5639 XI11_5/XI0/XI0_26/d_8_ XI11_5/XI0/XI0_26/d__8_ DECAP_INV_G11
XG5640 XI11_5/XI0/XI0_26/d_7_ XI11_5/XI0/XI0_26/d__7_ DECAP_INV_G11
XG5641 XI11_5/XI0/XI0_26/d_6_ XI11_5/XI0/XI0_26/d__6_ DECAP_INV_G11
XG5642 XI11_5/XI0/XI0_26/d_5_ XI11_5/XI0/XI0_26/d__5_ DECAP_INV_G11
XG5643 XI11_5/XI0/XI0_26/d_4_ XI11_5/XI0/XI0_26/d__4_ DECAP_INV_G11
XG5644 XI11_5/XI0/XI0_26/d_3_ XI11_5/XI0/XI0_26/d__3_ DECAP_INV_G11
XG5645 XI11_5/XI0/XI0_26/d_2_ XI11_5/XI0/XI0_26/d__2_ DECAP_INV_G11
XG5646 XI11_5/XI0/XI0_26/d_1_ XI11_5/XI0/XI0_26/d__1_ DECAP_INV_G11
XG5647 XI11_5/XI0/XI0_26/d_0_ XI11_5/XI0/XI0_26/d__0_ DECAP_INV_G11
XG5648 XI11_5/XI0/XI0_25/d__15_ XI11_5/XI0/XI0_25/d_15_ DECAP_INV_G11
XG5649 XI11_5/XI0/XI0_25/d__14_ XI11_5/XI0/XI0_25/d_14_ DECAP_INV_G11
XG5650 XI11_5/XI0/XI0_25/d__13_ XI11_5/XI0/XI0_25/d_13_ DECAP_INV_G11
XG5651 XI11_5/XI0/XI0_25/d__12_ XI11_5/XI0/XI0_25/d_12_ DECAP_INV_G11
XG5652 XI11_5/XI0/XI0_25/d__11_ XI11_5/XI0/XI0_25/d_11_ DECAP_INV_G11
XG5653 XI11_5/XI0/XI0_25/d__10_ XI11_5/XI0/XI0_25/d_10_ DECAP_INV_G11
XG5654 XI11_5/XI0/XI0_25/d__9_ XI11_5/XI0/XI0_25/d_9_ DECAP_INV_G11
XG5655 XI11_5/XI0/XI0_25/d__8_ XI11_5/XI0/XI0_25/d_8_ DECAP_INV_G11
XG5656 XI11_5/XI0/XI0_25/d__7_ XI11_5/XI0/XI0_25/d_7_ DECAP_INV_G11
XG5657 XI11_5/XI0/XI0_25/d__6_ XI11_5/XI0/XI0_25/d_6_ DECAP_INV_G11
XG5658 XI11_5/XI0/XI0_25/d__5_ XI11_5/XI0/XI0_25/d_5_ DECAP_INV_G11
XG5659 XI11_5/XI0/XI0_25/d__4_ XI11_5/XI0/XI0_25/d_4_ DECAP_INV_G11
XG5660 XI11_5/XI0/XI0_25/d__3_ XI11_5/XI0/XI0_25/d_3_ DECAP_INV_G11
XG5661 XI11_5/XI0/XI0_25/d__2_ XI11_5/XI0/XI0_25/d_2_ DECAP_INV_G11
XG5662 XI11_5/XI0/XI0_25/d__1_ XI11_5/XI0/XI0_25/d_1_ DECAP_INV_G11
XG5663 XI11_5/XI0/XI0_25/d__0_ XI11_5/XI0/XI0_25/d_0_ DECAP_INV_G11
XG5664 XI11_5/XI0/XI0_25/d_15_ XI11_5/XI0/XI0_25/d__15_ DECAP_INV_G11
XG5665 XI11_5/XI0/XI0_25/d_14_ XI11_5/XI0/XI0_25/d__14_ DECAP_INV_G11
XG5666 XI11_5/XI0/XI0_25/d_13_ XI11_5/XI0/XI0_25/d__13_ DECAP_INV_G11
XG5667 XI11_5/XI0/XI0_25/d_12_ XI11_5/XI0/XI0_25/d__12_ DECAP_INV_G11
XG5668 XI11_5/XI0/XI0_25/d_11_ XI11_5/XI0/XI0_25/d__11_ DECAP_INV_G11
XG5669 XI11_5/XI0/XI0_25/d_10_ XI11_5/XI0/XI0_25/d__10_ DECAP_INV_G11
XG5670 XI11_5/XI0/XI0_25/d_9_ XI11_5/XI0/XI0_25/d__9_ DECAP_INV_G11
XG5671 XI11_5/XI0/XI0_25/d_8_ XI11_5/XI0/XI0_25/d__8_ DECAP_INV_G11
XG5672 XI11_5/XI0/XI0_25/d_7_ XI11_5/XI0/XI0_25/d__7_ DECAP_INV_G11
XG5673 XI11_5/XI0/XI0_25/d_6_ XI11_5/XI0/XI0_25/d__6_ DECAP_INV_G11
XG5674 XI11_5/XI0/XI0_25/d_5_ XI11_5/XI0/XI0_25/d__5_ DECAP_INV_G11
XG5675 XI11_5/XI0/XI0_25/d_4_ XI11_5/XI0/XI0_25/d__4_ DECAP_INV_G11
XG5676 XI11_5/XI0/XI0_25/d_3_ XI11_5/XI0/XI0_25/d__3_ DECAP_INV_G11
XG5677 XI11_5/XI0/XI0_25/d_2_ XI11_5/XI0/XI0_25/d__2_ DECAP_INV_G11
XG5678 XI11_5/XI0/XI0_25/d_1_ XI11_5/XI0/XI0_25/d__1_ DECAP_INV_G11
XG5679 XI11_5/XI0/XI0_25/d_0_ XI11_5/XI0/XI0_25/d__0_ DECAP_INV_G11
XG5680 XI11_5/XI0/XI0_24/d__15_ XI11_5/XI0/XI0_24/d_15_ DECAP_INV_G11
XG5681 XI11_5/XI0/XI0_24/d__14_ XI11_5/XI0/XI0_24/d_14_ DECAP_INV_G11
XG5682 XI11_5/XI0/XI0_24/d__13_ XI11_5/XI0/XI0_24/d_13_ DECAP_INV_G11
XG5683 XI11_5/XI0/XI0_24/d__12_ XI11_5/XI0/XI0_24/d_12_ DECAP_INV_G11
XG5684 XI11_5/XI0/XI0_24/d__11_ XI11_5/XI0/XI0_24/d_11_ DECAP_INV_G11
XG5685 XI11_5/XI0/XI0_24/d__10_ XI11_5/XI0/XI0_24/d_10_ DECAP_INV_G11
XG5686 XI11_5/XI0/XI0_24/d__9_ XI11_5/XI0/XI0_24/d_9_ DECAP_INV_G11
XG5687 XI11_5/XI0/XI0_24/d__8_ XI11_5/XI0/XI0_24/d_8_ DECAP_INV_G11
XG5688 XI11_5/XI0/XI0_24/d__7_ XI11_5/XI0/XI0_24/d_7_ DECAP_INV_G11
XG5689 XI11_5/XI0/XI0_24/d__6_ XI11_5/XI0/XI0_24/d_6_ DECAP_INV_G11
XG5690 XI11_5/XI0/XI0_24/d__5_ XI11_5/XI0/XI0_24/d_5_ DECAP_INV_G11
XG5691 XI11_5/XI0/XI0_24/d__4_ XI11_5/XI0/XI0_24/d_4_ DECAP_INV_G11
XG5692 XI11_5/XI0/XI0_24/d__3_ XI11_5/XI0/XI0_24/d_3_ DECAP_INV_G11
XG5693 XI11_5/XI0/XI0_24/d__2_ XI11_5/XI0/XI0_24/d_2_ DECAP_INV_G11
XG5694 XI11_5/XI0/XI0_24/d__1_ XI11_5/XI0/XI0_24/d_1_ DECAP_INV_G11
XG5695 XI11_5/XI0/XI0_24/d__0_ XI11_5/XI0/XI0_24/d_0_ DECAP_INV_G11
XG5696 XI11_5/XI0/XI0_24/d_15_ XI11_5/XI0/XI0_24/d__15_ DECAP_INV_G11
XG5697 XI11_5/XI0/XI0_24/d_14_ XI11_5/XI0/XI0_24/d__14_ DECAP_INV_G11
XG5698 XI11_5/XI0/XI0_24/d_13_ XI11_5/XI0/XI0_24/d__13_ DECAP_INV_G11
XG5699 XI11_5/XI0/XI0_24/d_12_ XI11_5/XI0/XI0_24/d__12_ DECAP_INV_G11
XG5700 XI11_5/XI0/XI0_24/d_11_ XI11_5/XI0/XI0_24/d__11_ DECAP_INV_G11
XG5701 XI11_5/XI0/XI0_24/d_10_ XI11_5/XI0/XI0_24/d__10_ DECAP_INV_G11
XG5702 XI11_5/XI0/XI0_24/d_9_ XI11_5/XI0/XI0_24/d__9_ DECAP_INV_G11
XG5703 XI11_5/XI0/XI0_24/d_8_ XI11_5/XI0/XI0_24/d__8_ DECAP_INV_G11
XG5704 XI11_5/XI0/XI0_24/d_7_ XI11_5/XI0/XI0_24/d__7_ DECAP_INV_G11
XG5705 XI11_5/XI0/XI0_24/d_6_ XI11_5/XI0/XI0_24/d__6_ DECAP_INV_G11
XG5706 XI11_5/XI0/XI0_24/d_5_ XI11_5/XI0/XI0_24/d__5_ DECAP_INV_G11
XG5707 XI11_5/XI0/XI0_24/d_4_ XI11_5/XI0/XI0_24/d__4_ DECAP_INV_G11
XG5708 XI11_5/XI0/XI0_24/d_3_ XI11_5/XI0/XI0_24/d__3_ DECAP_INV_G11
XG5709 XI11_5/XI0/XI0_24/d_2_ XI11_5/XI0/XI0_24/d__2_ DECAP_INV_G11
XG5710 XI11_5/XI0/XI0_24/d_1_ XI11_5/XI0/XI0_24/d__1_ DECAP_INV_G11
XG5711 XI11_5/XI0/XI0_24/d_0_ XI11_5/XI0/XI0_24/d__0_ DECAP_INV_G11
XG5712 XI11_5/XI0/XI0_23/d__15_ XI11_5/XI0/XI0_23/d_15_ DECAP_INV_G11
XG5713 XI11_5/XI0/XI0_23/d__14_ XI11_5/XI0/XI0_23/d_14_ DECAP_INV_G11
XG5714 XI11_5/XI0/XI0_23/d__13_ XI11_5/XI0/XI0_23/d_13_ DECAP_INV_G11
XG5715 XI11_5/XI0/XI0_23/d__12_ XI11_5/XI0/XI0_23/d_12_ DECAP_INV_G11
XG5716 XI11_5/XI0/XI0_23/d__11_ XI11_5/XI0/XI0_23/d_11_ DECAP_INV_G11
XG5717 XI11_5/XI0/XI0_23/d__10_ XI11_5/XI0/XI0_23/d_10_ DECAP_INV_G11
XG5718 XI11_5/XI0/XI0_23/d__9_ XI11_5/XI0/XI0_23/d_9_ DECAP_INV_G11
XG5719 XI11_5/XI0/XI0_23/d__8_ XI11_5/XI0/XI0_23/d_8_ DECAP_INV_G11
XG5720 XI11_5/XI0/XI0_23/d__7_ XI11_5/XI0/XI0_23/d_7_ DECAP_INV_G11
XG5721 XI11_5/XI0/XI0_23/d__6_ XI11_5/XI0/XI0_23/d_6_ DECAP_INV_G11
XG5722 XI11_5/XI0/XI0_23/d__5_ XI11_5/XI0/XI0_23/d_5_ DECAP_INV_G11
XG5723 XI11_5/XI0/XI0_23/d__4_ XI11_5/XI0/XI0_23/d_4_ DECAP_INV_G11
XG5724 XI11_5/XI0/XI0_23/d__3_ XI11_5/XI0/XI0_23/d_3_ DECAP_INV_G11
XG5725 XI11_5/XI0/XI0_23/d__2_ XI11_5/XI0/XI0_23/d_2_ DECAP_INV_G11
XG5726 XI11_5/XI0/XI0_23/d__1_ XI11_5/XI0/XI0_23/d_1_ DECAP_INV_G11
XG5727 XI11_5/XI0/XI0_23/d__0_ XI11_5/XI0/XI0_23/d_0_ DECAP_INV_G11
XG5728 XI11_5/XI0/XI0_23/d_15_ XI11_5/XI0/XI0_23/d__15_ DECAP_INV_G11
XG5729 XI11_5/XI0/XI0_23/d_14_ XI11_5/XI0/XI0_23/d__14_ DECAP_INV_G11
XG5730 XI11_5/XI0/XI0_23/d_13_ XI11_5/XI0/XI0_23/d__13_ DECAP_INV_G11
XG5731 XI11_5/XI0/XI0_23/d_12_ XI11_5/XI0/XI0_23/d__12_ DECAP_INV_G11
XG5732 XI11_5/XI0/XI0_23/d_11_ XI11_5/XI0/XI0_23/d__11_ DECAP_INV_G11
XG5733 XI11_5/XI0/XI0_23/d_10_ XI11_5/XI0/XI0_23/d__10_ DECAP_INV_G11
XG5734 XI11_5/XI0/XI0_23/d_9_ XI11_5/XI0/XI0_23/d__9_ DECAP_INV_G11
XG5735 XI11_5/XI0/XI0_23/d_8_ XI11_5/XI0/XI0_23/d__8_ DECAP_INV_G11
XG5736 XI11_5/XI0/XI0_23/d_7_ XI11_5/XI0/XI0_23/d__7_ DECAP_INV_G11
XG5737 XI11_5/XI0/XI0_23/d_6_ XI11_5/XI0/XI0_23/d__6_ DECAP_INV_G11
XG5738 XI11_5/XI0/XI0_23/d_5_ XI11_5/XI0/XI0_23/d__5_ DECAP_INV_G11
XG5739 XI11_5/XI0/XI0_23/d_4_ XI11_5/XI0/XI0_23/d__4_ DECAP_INV_G11
XG5740 XI11_5/XI0/XI0_23/d_3_ XI11_5/XI0/XI0_23/d__3_ DECAP_INV_G11
XG5741 XI11_5/XI0/XI0_23/d_2_ XI11_5/XI0/XI0_23/d__2_ DECAP_INV_G11
XG5742 XI11_5/XI0/XI0_23/d_1_ XI11_5/XI0/XI0_23/d__1_ DECAP_INV_G11
XG5743 XI11_5/XI0/XI0_23/d_0_ XI11_5/XI0/XI0_23/d__0_ DECAP_INV_G11
XG5744 XI11_5/XI0/XI0_22/d__15_ XI11_5/XI0/XI0_22/d_15_ DECAP_INV_G11
XG5745 XI11_5/XI0/XI0_22/d__14_ XI11_5/XI0/XI0_22/d_14_ DECAP_INV_G11
XG5746 XI11_5/XI0/XI0_22/d__13_ XI11_5/XI0/XI0_22/d_13_ DECAP_INV_G11
XG5747 XI11_5/XI0/XI0_22/d__12_ XI11_5/XI0/XI0_22/d_12_ DECAP_INV_G11
XG5748 XI11_5/XI0/XI0_22/d__11_ XI11_5/XI0/XI0_22/d_11_ DECAP_INV_G11
XG5749 XI11_5/XI0/XI0_22/d__10_ XI11_5/XI0/XI0_22/d_10_ DECAP_INV_G11
XG5750 XI11_5/XI0/XI0_22/d__9_ XI11_5/XI0/XI0_22/d_9_ DECAP_INV_G11
XG5751 XI11_5/XI0/XI0_22/d__8_ XI11_5/XI0/XI0_22/d_8_ DECAP_INV_G11
XG5752 XI11_5/XI0/XI0_22/d__7_ XI11_5/XI0/XI0_22/d_7_ DECAP_INV_G11
XG5753 XI11_5/XI0/XI0_22/d__6_ XI11_5/XI0/XI0_22/d_6_ DECAP_INV_G11
XG5754 XI11_5/XI0/XI0_22/d__5_ XI11_5/XI0/XI0_22/d_5_ DECAP_INV_G11
XG5755 XI11_5/XI0/XI0_22/d__4_ XI11_5/XI0/XI0_22/d_4_ DECAP_INV_G11
XG5756 XI11_5/XI0/XI0_22/d__3_ XI11_5/XI0/XI0_22/d_3_ DECAP_INV_G11
XG5757 XI11_5/XI0/XI0_22/d__2_ XI11_5/XI0/XI0_22/d_2_ DECAP_INV_G11
XG5758 XI11_5/XI0/XI0_22/d__1_ XI11_5/XI0/XI0_22/d_1_ DECAP_INV_G11
XG5759 XI11_5/XI0/XI0_22/d__0_ XI11_5/XI0/XI0_22/d_0_ DECAP_INV_G11
XG5760 XI11_5/XI0/XI0_22/d_15_ XI11_5/XI0/XI0_22/d__15_ DECAP_INV_G11
XG5761 XI11_5/XI0/XI0_22/d_14_ XI11_5/XI0/XI0_22/d__14_ DECAP_INV_G11
XG5762 XI11_5/XI0/XI0_22/d_13_ XI11_5/XI0/XI0_22/d__13_ DECAP_INV_G11
XG5763 XI11_5/XI0/XI0_22/d_12_ XI11_5/XI0/XI0_22/d__12_ DECAP_INV_G11
XG5764 XI11_5/XI0/XI0_22/d_11_ XI11_5/XI0/XI0_22/d__11_ DECAP_INV_G11
XG5765 XI11_5/XI0/XI0_22/d_10_ XI11_5/XI0/XI0_22/d__10_ DECAP_INV_G11
XG5766 XI11_5/XI0/XI0_22/d_9_ XI11_5/XI0/XI0_22/d__9_ DECAP_INV_G11
XG5767 XI11_5/XI0/XI0_22/d_8_ XI11_5/XI0/XI0_22/d__8_ DECAP_INV_G11
XG5768 XI11_5/XI0/XI0_22/d_7_ XI11_5/XI0/XI0_22/d__7_ DECAP_INV_G11
XG5769 XI11_5/XI0/XI0_22/d_6_ XI11_5/XI0/XI0_22/d__6_ DECAP_INV_G11
XG5770 XI11_5/XI0/XI0_22/d_5_ XI11_5/XI0/XI0_22/d__5_ DECAP_INV_G11
XG5771 XI11_5/XI0/XI0_22/d_4_ XI11_5/XI0/XI0_22/d__4_ DECAP_INV_G11
XG5772 XI11_5/XI0/XI0_22/d_3_ XI11_5/XI0/XI0_22/d__3_ DECAP_INV_G11
XG5773 XI11_5/XI0/XI0_22/d_2_ XI11_5/XI0/XI0_22/d__2_ DECAP_INV_G11
XG5774 XI11_5/XI0/XI0_22/d_1_ XI11_5/XI0/XI0_22/d__1_ DECAP_INV_G11
XG5775 XI11_5/XI0/XI0_22/d_0_ XI11_5/XI0/XI0_22/d__0_ DECAP_INV_G11
XG5776 XI11_5/XI0/XI0_21/d__15_ XI11_5/XI0/XI0_21/d_15_ DECAP_INV_G11
XG5777 XI11_5/XI0/XI0_21/d__14_ XI11_5/XI0/XI0_21/d_14_ DECAP_INV_G11
XG5778 XI11_5/XI0/XI0_21/d__13_ XI11_5/XI0/XI0_21/d_13_ DECAP_INV_G11
XG5779 XI11_5/XI0/XI0_21/d__12_ XI11_5/XI0/XI0_21/d_12_ DECAP_INV_G11
XG5780 XI11_5/XI0/XI0_21/d__11_ XI11_5/XI0/XI0_21/d_11_ DECAP_INV_G11
XG5781 XI11_5/XI0/XI0_21/d__10_ XI11_5/XI0/XI0_21/d_10_ DECAP_INV_G11
XG5782 XI11_5/XI0/XI0_21/d__9_ XI11_5/XI0/XI0_21/d_9_ DECAP_INV_G11
XG5783 XI11_5/XI0/XI0_21/d__8_ XI11_5/XI0/XI0_21/d_8_ DECAP_INV_G11
XG5784 XI11_5/XI0/XI0_21/d__7_ XI11_5/XI0/XI0_21/d_7_ DECAP_INV_G11
XG5785 XI11_5/XI0/XI0_21/d__6_ XI11_5/XI0/XI0_21/d_6_ DECAP_INV_G11
XG5786 XI11_5/XI0/XI0_21/d__5_ XI11_5/XI0/XI0_21/d_5_ DECAP_INV_G11
XG5787 XI11_5/XI0/XI0_21/d__4_ XI11_5/XI0/XI0_21/d_4_ DECAP_INV_G11
XG5788 XI11_5/XI0/XI0_21/d__3_ XI11_5/XI0/XI0_21/d_3_ DECAP_INV_G11
XG5789 XI11_5/XI0/XI0_21/d__2_ XI11_5/XI0/XI0_21/d_2_ DECAP_INV_G11
XG5790 XI11_5/XI0/XI0_21/d__1_ XI11_5/XI0/XI0_21/d_1_ DECAP_INV_G11
XG5791 XI11_5/XI0/XI0_21/d__0_ XI11_5/XI0/XI0_21/d_0_ DECAP_INV_G11
XG5792 XI11_5/XI0/XI0_21/d_15_ XI11_5/XI0/XI0_21/d__15_ DECAP_INV_G11
XG5793 XI11_5/XI0/XI0_21/d_14_ XI11_5/XI0/XI0_21/d__14_ DECAP_INV_G11
XG5794 XI11_5/XI0/XI0_21/d_13_ XI11_5/XI0/XI0_21/d__13_ DECAP_INV_G11
XG5795 XI11_5/XI0/XI0_21/d_12_ XI11_5/XI0/XI0_21/d__12_ DECAP_INV_G11
XG5796 XI11_5/XI0/XI0_21/d_11_ XI11_5/XI0/XI0_21/d__11_ DECAP_INV_G11
XG5797 XI11_5/XI0/XI0_21/d_10_ XI11_5/XI0/XI0_21/d__10_ DECAP_INV_G11
XG5798 XI11_5/XI0/XI0_21/d_9_ XI11_5/XI0/XI0_21/d__9_ DECAP_INV_G11
XG5799 XI11_5/XI0/XI0_21/d_8_ XI11_5/XI0/XI0_21/d__8_ DECAP_INV_G11
XG5800 XI11_5/XI0/XI0_21/d_7_ XI11_5/XI0/XI0_21/d__7_ DECAP_INV_G11
XG5801 XI11_5/XI0/XI0_21/d_6_ XI11_5/XI0/XI0_21/d__6_ DECAP_INV_G11
XG5802 XI11_5/XI0/XI0_21/d_5_ XI11_5/XI0/XI0_21/d__5_ DECAP_INV_G11
XG5803 XI11_5/XI0/XI0_21/d_4_ XI11_5/XI0/XI0_21/d__4_ DECAP_INV_G11
XG5804 XI11_5/XI0/XI0_21/d_3_ XI11_5/XI0/XI0_21/d__3_ DECAP_INV_G11
XG5805 XI11_5/XI0/XI0_21/d_2_ XI11_5/XI0/XI0_21/d__2_ DECAP_INV_G11
XG5806 XI11_5/XI0/XI0_21/d_1_ XI11_5/XI0/XI0_21/d__1_ DECAP_INV_G11
XG5807 XI11_5/XI0/XI0_21/d_0_ XI11_5/XI0/XI0_21/d__0_ DECAP_INV_G11
XG5808 XI11_5/XI0/XI0_20/d__15_ XI11_5/XI0/XI0_20/d_15_ DECAP_INV_G11
XG5809 XI11_5/XI0/XI0_20/d__14_ XI11_5/XI0/XI0_20/d_14_ DECAP_INV_G11
XG5810 XI11_5/XI0/XI0_20/d__13_ XI11_5/XI0/XI0_20/d_13_ DECAP_INV_G11
XG5811 XI11_5/XI0/XI0_20/d__12_ XI11_5/XI0/XI0_20/d_12_ DECAP_INV_G11
XG5812 XI11_5/XI0/XI0_20/d__11_ XI11_5/XI0/XI0_20/d_11_ DECAP_INV_G11
XG5813 XI11_5/XI0/XI0_20/d__10_ XI11_5/XI0/XI0_20/d_10_ DECAP_INV_G11
XG5814 XI11_5/XI0/XI0_20/d__9_ XI11_5/XI0/XI0_20/d_9_ DECAP_INV_G11
XG5815 XI11_5/XI0/XI0_20/d__8_ XI11_5/XI0/XI0_20/d_8_ DECAP_INV_G11
XG5816 XI11_5/XI0/XI0_20/d__7_ XI11_5/XI0/XI0_20/d_7_ DECAP_INV_G11
XG5817 XI11_5/XI0/XI0_20/d__6_ XI11_5/XI0/XI0_20/d_6_ DECAP_INV_G11
XG5818 XI11_5/XI0/XI0_20/d__5_ XI11_5/XI0/XI0_20/d_5_ DECAP_INV_G11
XG5819 XI11_5/XI0/XI0_20/d__4_ XI11_5/XI0/XI0_20/d_4_ DECAP_INV_G11
XG5820 XI11_5/XI0/XI0_20/d__3_ XI11_5/XI0/XI0_20/d_3_ DECAP_INV_G11
XG5821 XI11_5/XI0/XI0_20/d__2_ XI11_5/XI0/XI0_20/d_2_ DECAP_INV_G11
XG5822 XI11_5/XI0/XI0_20/d__1_ XI11_5/XI0/XI0_20/d_1_ DECAP_INV_G11
XG5823 XI11_5/XI0/XI0_20/d__0_ XI11_5/XI0/XI0_20/d_0_ DECAP_INV_G11
XG5824 XI11_5/XI0/XI0_20/d_15_ XI11_5/XI0/XI0_20/d__15_ DECAP_INV_G11
XG5825 XI11_5/XI0/XI0_20/d_14_ XI11_5/XI0/XI0_20/d__14_ DECAP_INV_G11
XG5826 XI11_5/XI0/XI0_20/d_13_ XI11_5/XI0/XI0_20/d__13_ DECAP_INV_G11
XG5827 XI11_5/XI0/XI0_20/d_12_ XI11_5/XI0/XI0_20/d__12_ DECAP_INV_G11
XG5828 XI11_5/XI0/XI0_20/d_11_ XI11_5/XI0/XI0_20/d__11_ DECAP_INV_G11
XG5829 XI11_5/XI0/XI0_20/d_10_ XI11_5/XI0/XI0_20/d__10_ DECAP_INV_G11
XG5830 XI11_5/XI0/XI0_20/d_9_ XI11_5/XI0/XI0_20/d__9_ DECAP_INV_G11
XG5831 XI11_5/XI0/XI0_20/d_8_ XI11_5/XI0/XI0_20/d__8_ DECAP_INV_G11
XG5832 XI11_5/XI0/XI0_20/d_7_ XI11_5/XI0/XI0_20/d__7_ DECAP_INV_G11
XG5833 XI11_5/XI0/XI0_20/d_6_ XI11_5/XI0/XI0_20/d__6_ DECAP_INV_G11
XG5834 XI11_5/XI0/XI0_20/d_5_ XI11_5/XI0/XI0_20/d__5_ DECAP_INV_G11
XG5835 XI11_5/XI0/XI0_20/d_4_ XI11_5/XI0/XI0_20/d__4_ DECAP_INV_G11
XG5836 XI11_5/XI0/XI0_20/d_3_ XI11_5/XI0/XI0_20/d__3_ DECAP_INV_G11
XG5837 XI11_5/XI0/XI0_20/d_2_ XI11_5/XI0/XI0_20/d__2_ DECAP_INV_G11
XG5838 XI11_5/XI0/XI0_20/d_1_ XI11_5/XI0/XI0_20/d__1_ DECAP_INV_G11
XG5839 XI11_5/XI0/XI0_20/d_0_ XI11_5/XI0/XI0_20/d__0_ DECAP_INV_G11
XG5840 XI11_5/XI0/XI0_19/d__15_ XI11_5/XI0/XI0_19/d_15_ DECAP_INV_G11
XG5841 XI11_5/XI0/XI0_19/d__14_ XI11_5/XI0/XI0_19/d_14_ DECAP_INV_G11
XG5842 XI11_5/XI0/XI0_19/d__13_ XI11_5/XI0/XI0_19/d_13_ DECAP_INV_G11
XG5843 XI11_5/XI0/XI0_19/d__12_ XI11_5/XI0/XI0_19/d_12_ DECAP_INV_G11
XG5844 XI11_5/XI0/XI0_19/d__11_ XI11_5/XI0/XI0_19/d_11_ DECAP_INV_G11
XG5845 XI11_5/XI0/XI0_19/d__10_ XI11_5/XI0/XI0_19/d_10_ DECAP_INV_G11
XG5846 XI11_5/XI0/XI0_19/d__9_ XI11_5/XI0/XI0_19/d_9_ DECAP_INV_G11
XG5847 XI11_5/XI0/XI0_19/d__8_ XI11_5/XI0/XI0_19/d_8_ DECAP_INV_G11
XG5848 XI11_5/XI0/XI0_19/d__7_ XI11_5/XI0/XI0_19/d_7_ DECAP_INV_G11
XG5849 XI11_5/XI0/XI0_19/d__6_ XI11_5/XI0/XI0_19/d_6_ DECAP_INV_G11
XG5850 XI11_5/XI0/XI0_19/d__5_ XI11_5/XI0/XI0_19/d_5_ DECAP_INV_G11
XG5851 XI11_5/XI0/XI0_19/d__4_ XI11_5/XI0/XI0_19/d_4_ DECAP_INV_G11
XG5852 XI11_5/XI0/XI0_19/d__3_ XI11_5/XI0/XI0_19/d_3_ DECAP_INV_G11
XG5853 XI11_5/XI0/XI0_19/d__2_ XI11_5/XI0/XI0_19/d_2_ DECAP_INV_G11
XG5854 XI11_5/XI0/XI0_19/d__1_ XI11_5/XI0/XI0_19/d_1_ DECAP_INV_G11
XG5855 XI11_5/XI0/XI0_19/d__0_ XI11_5/XI0/XI0_19/d_0_ DECAP_INV_G11
XG5856 XI11_5/XI0/XI0_19/d_15_ XI11_5/XI0/XI0_19/d__15_ DECAP_INV_G11
XG5857 XI11_5/XI0/XI0_19/d_14_ XI11_5/XI0/XI0_19/d__14_ DECAP_INV_G11
XG5858 XI11_5/XI0/XI0_19/d_13_ XI11_5/XI0/XI0_19/d__13_ DECAP_INV_G11
XG5859 XI11_5/XI0/XI0_19/d_12_ XI11_5/XI0/XI0_19/d__12_ DECAP_INV_G11
XG5860 XI11_5/XI0/XI0_19/d_11_ XI11_5/XI0/XI0_19/d__11_ DECAP_INV_G11
XG5861 XI11_5/XI0/XI0_19/d_10_ XI11_5/XI0/XI0_19/d__10_ DECAP_INV_G11
XG5862 XI11_5/XI0/XI0_19/d_9_ XI11_5/XI0/XI0_19/d__9_ DECAP_INV_G11
XG5863 XI11_5/XI0/XI0_19/d_8_ XI11_5/XI0/XI0_19/d__8_ DECAP_INV_G11
XG5864 XI11_5/XI0/XI0_19/d_7_ XI11_5/XI0/XI0_19/d__7_ DECAP_INV_G11
XG5865 XI11_5/XI0/XI0_19/d_6_ XI11_5/XI0/XI0_19/d__6_ DECAP_INV_G11
XG5866 XI11_5/XI0/XI0_19/d_5_ XI11_5/XI0/XI0_19/d__5_ DECAP_INV_G11
XG5867 XI11_5/XI0/XI0_19/d_4_ XI11_5/XI0/XI0_19/d__4_ DECAP_INV_G11
XG5868 XI11_5/XI0/XI0_19/d_3_ XI11_5/XI0/XI0_19/d__3_ DECAP_INV_G11
XG5869 XI11_5/XI0/XI0_19/d_2_ XI11_5/XI0/XI0_19/d__2_ DECAP_INV_G11
XG5870 XI11_5/XI0/XI0_19/d_1_ XI11_5/XI0/XI0_19/d__1_ DECAP_INV_G11
XG5871 XI11_5/XI0/XI0_19/d_0_ XI11_5/XI0/XI0_19/d__0_ DECAP_INV_G11
XG5872 XI11_5/XI0/XI0_18/d__15_ XI11_5/XI0/XI0_18/d_15_ DECAP_INV_G11
XG5873 XI11_5/XI0/XI0_18/d__14_ XI11_5/XI0/XI0_18/d_14_ DECAP_INV_G11
XG5874 XI11_5/XI0/XI0_18/d__13_ XI11_5/XI0/XI0_18/d_13_ DECAP_INV_G11
XG5875 XI11_5/XI0/XI0_18/d__12_ XI11_5/XI0/XI0_18/d_12_ DECAP_INV_G11
XG5876 XI11_5/XI0/XI0_18/d__11_ XI11_5/XI0/XI0_18/d_11_ DECAP_INV_G11
XG5877 XI11_5/XI0/XI0_18/d__10_ XI11_5/XI0/XI0_18/d_10_ DECAP_INV_G11
XG5878 XI11_5/XI0/XI0_18/d__9_ XI11_5/XI0/XI0_18/d_9_ DECAP_INV_G11
XG5879 XI11_5/XI0/XI0_18/d__8_ XI11_5/XI0/XI0_18/d_8_ DECAP_INV_G11
XG5880 XI11_5/XI0/XI0_18/d__7_ XI11_5/XI0/XI0_18/d_7_ DECAP_INV_G11
XG5881 XI11_5/XI0/XI0_18/d__6_ XI11_5/XI0/XI0_18/d_6_ DECAP_INV_G11
XG5882 XI11_5/XI0/XI0_18/d__5_ XI11_5/XI0/XI0_18/d_5_ DECAP_INV_G11
XG5883 XI11_5/XI0/XI0_18/d__4_ XI11_5/XI0/XI0_18/d_4_ DECAP_INV_G11
XG5884 XI11_5/XI0/XI0_18/d__3_ XI11_5/XI0/XI0_18/d_3_ DECAP_INV_G11
XG5885 XI11_5/XI0/XI0_18/d__2_ XI11_5/XI0/XI0_18/d_2_ DECAP_INV_G11
XG5886 XI11_5/XI0/XI0_18/d__1_ XI11_5/XI0/XI0_18/d_1_ DECAP_INV_G11
XG5887 XI11_5/XI0/XI0_18/d__0_ XI11_5/XI0/XI0_18/d_0_ DECAP_INV_G11
XG5888 XI11_5/XI0/XI0_18/d_15_ XI11_5/XI0/XI0_18/d__15_ DECAP_INV_G11
XG5889 XI11_5/XI0/XI0_18/d_14_ XI11_5/XI0/XI0_18/d__14_ DECAP_INV_G11
XG5890 XI11_5/XI0/XI0_18/d_13_ XI11_5/XI0/XI0_18/d__13_ DECAP_INV_G11
XG5891 XI11_5/XI0/XI0_18/d_12_ XI11_5/XI0/XI0_18/d__12_ DECAP_INV_G11
XG5892 XI11_5/XI0/XI0_18/d_11_ XI11_5/XI0/XI0_18/d__11_ DECAP_INV_G11
XG5893 XI11_5/XI0/XI0_18/d_10_ XI11_5/XI0/XI0_18/d__10_ DECAP_INV_G11
XG5894 XI11_5/XI0/XI0_18/d_9_ XI11_5/XI0/XI0_18/d__9_ DECAP_INV_G11
XG5895 XI11_5/XI0/XI0_18/d_8_ XI11_5/XI0/XI0_18/d__8_ DECAP_INV_G11
XG5896 XI11_5/XI0/XI0_18/d_7_ XI11_5/XI0/XI0_18/d__7_ DECAP_INV_G11
XG5897 XI11_5/XI0/XI0_18/d_6_ XI11_5/XI0/XI0_18/d__6_ DECAP_INV_G11
XG5898 XI11_5/XI0/XI0_18/d_5_ XI11_5/XI0/XI0_18/d__5_ DECAP_INV_G11
XG5899 XI11_5/XI0/XI0_18/d_4_ XI11_5/XI0/XI0_18/d__4_ DECAP_INV_G11
XG5900 XI11_5/XI0/XI0_18/d_3_ XI11_5/XI0/XI0_18/d__3_ DECAP_INV_G11
XG5901 XI11_5/XI0/XI0_18/d_2_ XI11_5/XI0/XI0_18/d__2_ DECAP_INV_G11
XG5902 XI11_5/XI0/XI0_18/d_1_ XI11_5/XI0/XI0_18/d__1_ DECAP_INV_G11
XG5903 XI11_5/XI0/XI0_18/d_0_ XI11_5/XI0/XI0_18/d__0_ DECAP_INV_G11
XG5904 XI11_5/XI0/XI0_17/d__15_ XI11_5/XI0/XI0_17/d_15_ DECAP_INV_G11
XG5905 XI11_5/XI0/XI0_17/d__14_ XI11_5/XI0/XI0_17/d_14_ DECAP_INV_G11
XG5906 XI11_5/XI0/XI0_17/d__13_ XI11_5/XI0/XI0_17/d_13_ DECAP_INV_G11
XG5907 XI11_5/XI0/XI0_17/d__12_ XI11_5/XI0/XI0_17/d_12_ DECAP_INV_G11
XG5908 XI11_5/XI0/XI0_17/d__11_ XI11_5/XI0/XI0_17/d_11_ DECAP_INV_G11
XG5909 XI11_5/XI0/XI0_17/d__10_ XI11_5/XI0/XI0_17/d_10_ DECAP_INV_G11
XG5910 XI11_5/XI0/XI0_17/d__9_ XI11_5/XI0/XI0_17/d_9_ DECAP_INV_G11
XG5911 XI11_5/XI0/XI0_17/d__8_ XI11_5/XI0/XI0_17/d_8_ DECAP_INV_G11
XG5912 XI11_5/XI0/XI0_17/d__7_ XI11_5/XI0/XI0_17/d_7_ DECAP_INV_G11
XG5913 XI11_5/XI0/XI0_17/d__6_ XI11_5/XI0/XI0_17/d_6_ DECAP_INV_G11
XG5914 XI11_5/XI0/XI0_17/d__5_ XI11_5/XI0/XI0_17/d_5_ DECAP_INV_G11
XG5915 XI11_5/XI0/XI0_17/d__4_ XI11_5/XI0/XI0_17/d_4_ DECAP_INV_G11
XG5916 XI11_5/XI0/XI0_17/d__3_ XI11_5/XI0/XI0_17/d_3_ DECAP_INV_G11
XG5917 XI11_5/XI0/XI0_17/d__2_ XI11_5/XI0/XI0_17/d_2_ DECAP_INV_G11
XG5918 XI11_5/XI0/XI0_17/d__1_ XI11_5/XI0/XI0_17/d_1_ DECAP_INV_G11
XG5919 XI11_5/XI0/XI0_17/d__0_ XI11_5/XI0/XI0_17/d_0_ DECAP_INV_G11
XG5920 XI11_5/XI0/XI0_17/d_15_ XI11_5/XI0/XI0_17/d__15_ DECAP_INV_G11
XG5921 XI11_5/XI0/XI0_17/d_14_ XI11_5/XI0/XI0_17/d__14_ DECAP_INV_G11
XG5922 XI11_5/XI0/XI0_17/d_13_ XI11_5/XI0/XI0_17/d__13_ DECAP_INV_G11
XG5923 XI11_5/XI0/XI0_17/d_12_ XI11_5/XI0/XI0_17/d__12_ DECAP_INV_G11
XG5924 XI11_5/XI0/XI0_17/d_11_ XI11_5/XI0/XI0_17/d__11_ DECAP_INV_G11
XG5925 XI11_5/XI0/XI0_17/d_10_ XI11_5/XI0/XI0_17/d__10_ DECAP_INV_G11
XG5926 XI11_5/XI0/XI0_17/d_9_ XI11_5/XI0/XI0_17/d__9_ DECAP_INV_G11
XG5927 XI11_5/XI0/XI0_17/d_8_ XI11_5/XI0/XI0_17/d__8_ DECAP_INV_G11
XG5928 XI11_5/XI0/XI0_17/d_7_ XI11_5/XI0/XI0_17/d__7_ DECAP_INV_G11
XG5929 XI11_5/XI0/XI0_17/d_6_ XI11_5/XI0/XI0_17/d__6_ DECAP_INV_G11
XG5930 XI11_5/XI0/XI0_17/d_5_ XI11_5/XI0/XI0_17/d__5_ DECAP_INV_G11
XG5931 XI11_5/XI0/XI0_17/d_4_ XI11_5/XI0/XI0_17/d__4_ DECAP_INV_G11
XG5932 XI11_5/XI0/XI0_17/d_3_ XI11_5/XI0/XI0_17/d__3_ DECAP_INV_G11
XG5933 XI11_5/XI0/XI0_17/d_2_ XI11_5/XI0/XI0_17/d__2_ DECAP_INV_G11
XG5934 XI11_5/XI0/XI0_17/d_1_ XI11_5/XI0/XI0_17/d__1_ DECAP_INV_G11
XG5935 XI11_5/XI0/XI0_17/d_0_ XI11_5/XI0/XI0_17/d__0_ DECAP_INV_G11
XG5936 XI11_5/XI0/XI0_16/d__15_ XI11_5/XI0/XI0_16/d_15_ DECAP_INV_G11
XG5937 XI11_5/XI0/XI0_16/d__14_ XI11_5/XI0/XI0_16/d_14_ DECAP_INV_G11
XG5938 XI11_5/XI0/XI0_16/d__13_ XI11_5/XI0/XI0_16/d_13_ DECAP_INV_G11
XG5939 XI11_5/XI0/XI0_16/d__12_ XI11_5/XI0/XI0_16/d_12_ DECAP_INV_G11
XG5940 XI11_5/XI0/XI0_16/d__11_ XI11_5/XI0/XI0_16/d_11_ DECAP_INV_G11
XG5941 XI11_5/XI0/XI0_16/d__10_ XI11_5/XI0/XI0_16/d_10_ DECAP_INV_G11
XG5942 XI11_5/XI0/XI0_16/d__9_ XI11_5/XI0/XI0_16/d_9_ DECAP_INV_G11
XG5943 XI11_5/XI0/XI0_16/d__8_ XI11_5/XI0/XI0_16/d_8_ DECAP_INV_G11
XG5944 XI11_5/XI0/XI0_16/d__7_ XI11_5/XI0/XI0_16/d_7_ DECAP_INV_G11
XG5945 XI11_5/XI0/XI0_16/d__6_ XI11_5/XI0/XI0_16/d_6_ DECAP_INV_G11
XG5946 XI11_5/XI0/XI0_16/d__5_ XI11_5/XI0/XI0_16/d_5_ DECAP_INV_G11
XG5947 XI11_5/XI0/XI0_16/d__4_ XI11_5/XI0/XI0_16/d_4_ DECAP_INV_G11
XG5948 XI11_5/XI0/XI0_16/d__3_ XI11_5/XI0/XI0_16/d_3_ DECAP_INV_G11
XG5949 XI11_5/XI0/XI0_16/d__2_ XI11_5/XI0/XI0_16/d_2_ DECAP_INV_G11
XG5950 XI11_5/XI0/XI0_16/d__1_ XI11_5/XI0/XI0_16/d_1_ DECAP_INV_G11
XG5951 XI11_5/XI0/XI0_16/d__0_ XI11_5/XI0/XI0_16/d_0_ DECAP_INV_G11
XG5952 XI11_5/XI0/XI0_16/d_15_ XI11_5/XI0/XI0_16/d__15_ DECAP_INV_G11
XG5953 XI11_5/XI0/XI0_16/d_14_ XI11_5/XI0/XI0_16/d__14_ DECAP_INV_G11
XG5954 XI11_5/XI0/XI0_16/d_13_ XI11_5/XI0/XI0_16/d__13_ DECAP_INV_G11
XG5955 XI11_5/XI0/XI0_16/d_12_ XI11_5/XI0/XI0_16/d__12_ DECAP_INV_G11
XG5956 XI11_5/XI0/XI0_16/d_11_ XI11_5/XI0/XI0_16/d__11_ DECAP_INV_G11
XG5957 XI11_5/XI0/XI0_16/d_10_ XI11_5/XI0/XI0_16/d__10_ DECAP_INV_G11
XG5958 XI11_5/XI0/XI0_16/d_9_ XI11_5/XI0/XI0_16/d__9_ DECAP_INV_G11
XG5959 XI11_5/XI0/XI0_16/d_8_ XI11_5/XI0/XI0_16/d__8_ DECAP_INV_G11
XG5960 XI11_5/XI0/XI0_16/d_7_ XI11_5/XI0/XI0_16/d__7_ DECAP_INV_G11
XG5961 XI11_5/XI0/XI0_16/d_6_ XI11_5/XI0/XI0_16/d__6_ DECAP_INV_G11
XG5962 XI11_5/XI0/XI0_16/d_5_ XI11_5/XI0/XI0_16/d__5_ DECAP_INV_G11
XG5963 XI11_5/XI0/XI0_16/d_4_ XI11_5/XI0/XI0_16/d__4_ DECAP_INV_G11
XG5964 XI11_5/XI0/XI0_16/d_3_ XI11_5/XI0/XI0_16/d__3_ DECAP_INV_G11
XG5965 XI11_5/XI0/XI0_16/d_2_ XI11_5/XI0/XI0_16/d__2_ DECAP_INV_G11
XG5966 XI11_5/XI0/XI0_16/d_1_ XI11_5/XI0/XI0_16/d__1_ DECAP_INV_G11
XG5967 XI11_5/XI0/XI0_16/d_0_ XI11_5/XI0/XI0_16/d__0_ DECAP_INV_G11
XG5968 XI11_5/XI0/XI0_15/d__15_ XI11_5/XI0/XI0_15/d_15_ DECAP_INV_G11
XG5969 XI11_5/XI0/XI0_15/d__14_ XI11_5/XI0/XI0_15/d_14_ DECAP_INV_G11
XG5970 XI11_5/XI0/XI0_15/d__13_ XI11_5/XI0/XI0_15/d_13_ DECAP_INV_G11
XG5971 XI11_5/XI0/XI0_15/d__12_ XI11_5/XI0/XI0_15/d_12_ DECAP_INV_G11
XG5972 XI11_5/XI0/XI0_15/d__11_ XI11_5/XI0/XI0_15/d_11_ DECAP_INV_G11
XG5973 XI11_5/XI0/XI0_15/d__10_ XI11_5/XI0/XI0_15/d_10_ DECAP_INV_G11
XG5974 XI11_5/XI0/XI0_15/d__9_ XI11_5/XI0/XI0_15/d_9_ DECAP_INV_G11
XG5975 XI11_5/XI0/XI0_15/d__8_ XI11_5/XI0/XI0_15/d_8_ DECAP_INV_G11
XG5976 XI11_5/XI0/XI0_15/d__7_ XI11_5/XI0/XI0_15/d_7_ DECAP_INV_G11
XG5977 XI11_5/XI0/XI0_15/d__6_ XI11_5/XI0/XI0_15/d_6_ DECAP_INV_G11
XG5978 XI11_5/XI0/XI0_15/d__5_ XI11_5/XI0/XI0_15/d_5_ DECAP_INV_G11
XG5979 XI11_5/XI0/XI0_15/d__4_ XI11_5/XI0/XI0_15/d_4_ DECAP_INV_G11
XG5980 XI11_5/XI0/XI0_15/d__3_ XI11_5/XI0/XI0_15/d_3_ DECAP_INV_G11
XG5981 XI11_5/XI0/XI0_15/d__2_ XI11_5/XI0/XI0_15/d_2_ DECAP_INV_G11
XG5982 XI11_5/XI0/XI0_15/d__1_ XI11_5/XI0/XI0_15/d_1_ DECAP_INV_G11
XG5983 XI11_5/XI0/XI0_15/d__0_ XI11_5/XI0/XI0_15/d_0_ DECAP_INV_G11
XG5984 XI11_5/XI0/XI0_15/d_15_ XI11_5/XI0/XI0_15/d__15_ DECAP_INV_G11
XG5985 XI11_5/XI0/XI0_15/d_14_ XI11_5/XI0/XI0_15/d__14_ DECAP_INV_G11
XG5986 XI11_5/XI0/XI0_15/d_13_ XI11_5/XI0/XI0_15/d__13_ DECAP_INV_G11
XG5987 XI11_5/XI0/XI0_15/d_12_ XI11_5/XI0/XI0_15/d__12_ DECAP_INV_G11
XG5988 XI11_5/XI0/XI0_15/d_11_ XI11_5/XI0/XI0_15/d__11_ DECAP_INV_G11
XG5989 XI11_5/XI0/XI0_15/d_10_ XI11_5/XI0/XI0_15/d__10_ DECAP_INV_G11
XG5990 XI11_5/XI0/XI0_15/d_9_ XI11_5/XI0/XI0_15/d__9_ DECAP_INV_G11
XG5991 XI11_5/XI0/XI0_15/d_8_ XI11_5/XI0/XI0_15/d__8_ DECAP_INV_G11
XG5992 XI11_5/XI0/XI0_15/d_7_ XI11_5/XI0/XI0_15/d__7_ DECAP_INV_G11
XG5993 XI11_5/XI0/XI0_15/d_6_ XI11_5/XI0/XI0_15/d__6_ DECAP_INV_G11
XG5994 XI11_5/XI0/XI0_15/d_5_ XI11_5/XI0/XI0_15/d__5_ DECAP_INV_G11
XG5995 XI11_5/XI0/XI0_15/d_4_ XI11_5/XI0/XI0_15/d__4_ DECAP_INV_G11
XG5996 XI11_5/XI0/XI0_15/d_3_ XI11_5/XI0/XI0_15/d__3_ DECAP_INV_G11
XG5997 XI11_5/XI0/XI0_15/d_2_ XI11_5/XI0/XI0_15/d__2_ DECAP_INV_G11
XG5998 XI11_5/XI0/XI0_15/d_1_ XI11_5/XI0/XI0_15/d__1_ DECAP_INV_G11
XG5999 XI11_5/XI0/XI0_15/d_0_ XI11_5/XI0/XI0_15/d__0_ DECAP_INV_G11
XG6000 XI11_5/XI0/XI0_14/d__15_ XI11_5/XI0/XI0_14/d_15_ DECAP_INV_G11
XG6001 XI11_5/XI0/XI0_14/d__14_ XI11_5/XI0/XI0_14/d_14_ DECAP_INV_G11
XG6002 XI11_5/XI0/XI0_14/d__13_ XI11_5/XI0/XI0_14/d_13_ DECAP_INV_G11
XG6003 XI11_5/XI0/XI0_14/d__12_ XI11_5/XI0/XI0_14/d_12_ DECAP_INV_G11
XG6004 XI11_5/XI0/XI0_14/d__11_ XI11_5/XI0/XI0_14/d_11_ DECAP_INV_G11
XG6005 XI11_5/XI0/XI0_14/d__10_ XI11_5/XI0/XI0_14/d_10_ DECAP_INV_G11
XG6006 XI11_5/XI0/XI0_14/d__9_ XI11_5/XI0/XI0_14/d_9_ DECAP_INV_G11
XG6007 XI11_5/XI0/XI0_14/d__8_ XI11_5/XI0/XI0_14/d_8_ DECAP_INV_G11
XG6008 XI11_5/XI0/XI0_14/d__7_ XI11_5/XI0/XI0_14/d_7_ DECAP_INV_G11
XG6009 XI11_5/XI0/XI0_14/d__6_ XI11_5/XI0/XI0_14/d_6_ DECAP_INV_G11
XG6010 XI11_5/XI0/XI0_14/d__5_ XI11_5/XI0/XI0_14/d_5_ DECAP_INV_G11
XG6011 XI11_5/XI0/XI0_14/d__4_ XI11_5/XI0/XI0_14/d_4_ DECAP_INV_G11
XG6012 XI11_5/XI0/XI0_14/d__3_ XI11_5/XI0/XI0_14/d_3_ DECAP_INV_G11
XG6013 XI11_5/XI0/XI0_14/d__2_ XI11_5/XI0/XI0_14/d_2_ DECAP_INV_G11
XG6014 XI11_5/XI0/XI0_14/d__1_ XI11_5/XI0/XI0_14/d_1_ DECAP_INV_G11
XG6015 XI11_5/XI0/XI0_14/d__0_ XI11_5/XI0/XI0_14/d_0_ DECAP_INV_G11
XG6016 XI11_5/XI0/XI0_14/d_15_ XI11_5/XI0/XI0_14/d__15_ DECAP_INV_G11
XG6017 XI11_5/XI0/XI0_14/d_14_ XI11_5/XI0/XI0_14/d__14_ DECAP_INV_G11
XG6018 XI11_5/XI0/XI0_14/d_13_ XI11_5/XI0/XI0_14/d__13_ DECAP_INV_G11
XG6019 XI11_5/XI0/XI0_14/d_12_ XI11_5/XI0/XI0_14/d__12_ DECAP_INV_G11
XG6020 XI11_5/XI0/XI0_14/d_11_ XI11_5/XI0/XI0_14/d__11_ DECAP_INV_G11
XG6021 XI11_5/XI0/XI0_14/d_10_ XI11_5/XI0/XI0_14/d__10_ DECAP_INV_G11
XG6022 XI11_5/XI0/XI0_14/d_9_ XI11_5/XI0/XI0_14/d__9_ DECAP_INV_G11
XG6023 XI11_5/XI0/XI0_14/d_8_ XI11_5/XI0/XI0_14/d__8_ DECAP_INV_G11
XG6024 XI11_5/XI0/XI0_14/d_7_ XI11_5/XI0/XI0_14/d__7_ DECAP_INV_G11
XG6025 XI11_5/XI0/XI0_14/d_6_ XI11_5/XI0/XI0_14/d__6_ DECAP_INV_G11
XG6026 XI11_5/XI0/XI0_14/d_5_ XI11_5/XI0/XI0_14/d__5_ DECAP_INV_G11
XG6027 XI11_5/XI0/XI0_14/d_4_ XI11_5/XI0/XI0_14/d__4_ DECAP_INV_G11
XG6028 XI11_5/XI0/XI0_14/d_3_ XI11_5/XI0/XI0_14/d__3_ DECAP_INV_G11
XG6029 XI11_5/XI0/XI0_14/d_2_ XI11_5/XI0/XI0_14/d__2_ DECAP_INV_G11
XG6030 XI11_5/XI0/XI0_14/d_1_ XI11_5/XI0/XI0_14/d__1_ DECAP_INV_G11
XG6031 XI11_5/XI0/XI0_14/d_0_ XI11_5/XI0/XI0_14/d__0_ DECAP_INV_G11
XG6032 XI11_5/XI0/XI0_13/d__15_ XI11_5/XI0/XI0_13/d_15_ DECAP_INV_G11
XG6033 XI11_5/XI0/XI0_13/d__14_ XI11_5/XI0/XI0_13/d_14_ DECAP_INV_G11
XG6034 XI11_5/XI0/XI0_13/d__13_ XI11_5/XI0/XI0_13/d_13_ DECAP_INV_G11
XG6035 XI11_5/XI0/XI0_13/d__12_ XI11_5/XI0/XI0_13/d_12_ DECAP_INV_G11
XG6036 XI11_5/XI0/XI0_13/d__11_ XI11_5/XI0/XI0_13/d_11_ DECAP_INV_G11
XG6037 XI11_5/XI0/XI0_13/d__10_ XI11_5/XI0/XI0_13/d_10_ DECAP_INV_G11
XG6038 XI11_5/XI0/XI0_13/d__9_ XI11_5/XI0/XI0_13/d_9_ DECAP_INV_G11
XG6039 XI11_5/XI0/XI0_13/d__8_ XI11_5/XI0/XI0_13/d_8_ DECAP_INV_G11
XG6040 XI11_5/XI0/XI0_13/d__7_ XI11_5/XI0/XI0_13/d_7_ DECAP_INV_G11
XG6041 XI11_5/XI0/XI0_13/d__6_ XI11_5/XI0/XI0_13/d_6_ DECAP_INV_G11
XG6042 XI11_5/XI0/XI0_13/d__5_ XI11_5/XI0/XI0_13/d_5_ DECAP_INV_G11
XG6043 XI11_5/XI0/XI0_13/d__4_ XI11_5/XI0/XI0_13/d_4_ DECAP_INV_G11
XG6044 XI11_5/XI0/XI0_13/d__3_ XI11_5/XI0/XI0_13/d_3_ DECAP_INV_G11
XG6045 XI11_5/XI0/XI0_13/d__2_ XI11_5/XI0/XI0_13/d_2_ DECAP_INV_G11
XG6046 XI11_5/XI0/XI0_13/d__1_ XI11_5/XI0/XI0_13/d_1_ DECAP_INV_G11
XG6047 XI11_5/XI0/XI0_13/d__0_ XI11_5/XI0/XI0_13/d_0_ DECAP_INV_G11
XG6048 XI11_5/XI0/XI0_13/d_15_ XI11_5/XI0/XI0_13/d__15_ DECAP_INV_G11
XG6049 XI11_5/XI0/XI0_13/d_14_ XI11_5/XI0/XI0_13/d__14_ DECAP_INV_G11
XG6050 XI11_5/XI0/XI0_13/d_13_ XI11_5/XI0/XI0_13/d__13_ DECAP_INV_G11
XG6051 XI11_5/XI0/XI0_13/d_12_ XI11_5/XI0/XI0_13/d__12_ DECAP_INV_G11
XG6052 XI11_5/XI0/XI0_13/d_11_ XI11_5/XI0/XI0_13/d__11_ DECAP_INV_G11
XG6053 XI11_5/XI0/XI0_13/d_10_ XI11_5/XI0/XI0_13/d__10_ DECAP_INV_G11
XG6054 XI11_5/XI0/XI0_13/d_9_ XI11_5/XI0/XI0_13/d__9_ DECAP_INV_G11
XG6055 XI11_5/XI0/XI0_13/d_8_ XI11_5/XI0/XI0_13/d__8_ DECAP_INV_G11
XG6056 XI11_5/XI0/XI0_13/d_7_ XI11_5/XI0/XI0_13/d__7_ DECAP_INV_G11
XG6057 XI11_5/XI0/XI0_13/d_6_ XI11_5/XI0/XI0_13/d__6_ DECAP_INV_G11
XG6058 XI11_5/XI0/XI0_13/d_5_ XI11_5/XI0/XI0_13/d__5_ DECAP_INV_G11
XG6059 XI11_5/XI0/XI0_13/d_4_ XI11_5/XI0/XI0_13/d__4_ DECAP_INV_G11
XG6060 XI11_5/XI0/XI0_13/d_3_ XI11_5/XI0/XI0_13/d__3_ DECAP_INV_G11
XG6061 XI11_5/XI0/XI0_13/d_2_ XI11_5/XI0/XI0_13/d__2_ DECAP_INV_G11
XG6062 XI11_5/XI0/XI0_13/d_1_ XI11_5/XI0/XI0_13/d__1_ DECAP_INV_G11
XG6063 XI11_5/XI0/XI0_13/d_0_ XI11_5/XI0/XI0_13/d__0_ DECAP_INV_G11
XG6064 XI11_5/XI0/XI0_12/d__15_ XI11_5/XI0/XI0_12/d_15_ DECAP_INV_G11
XG6065 XI11_5/XI0/XI0_12/d__14_ XI11_5/XI0/XI0_12/d_14_ DECAP_INV_G11
XG6066 XI11_5/XI0/XI0_12/d__13_ XI11_5/XI0/XI0_12/d_13_ DECAP_INV_G11
XG6067 XI11_5/XI0/XI0_12/d__12_ XI11_5/XI0/XI0_12/d_12_ DECAP_INV_G11
XG6068 XI11_5/XI0/XI0_12/d__11_ XI11_5/XI0/XI0_12/d_11_ DECAP_INV_G11
XG6069 XI11_5/XI0/XI0_12/d__10_ XI11_5/XI0/XI0_12/d_10_ DECAP_INV_G11
XG6070 XI11_5/XI0/XI0_12/d__9_ XI11_5/XI0/XI0_12/d_9_ DECAP_INV_G11
XG6071 XI11_5/XI0/XI0_12/d__8_ XI11_5/XI0/XI0_12/d_8_ DECAP_INV_G11
XG6072 XI11_5/XI0/XI0_12/d__7_ XI11_5/XI0/XI0_12/d_7_ DECAP_INV_G11
XG6073 XI11_5/XI0/XI0_12/d__6_ XI11_5/XI0/XI0_12/d_6_ DECAP_INV_G11
XG6074 XI11_5/XI0/XI0_12/d__5_ XI11_5/XI0/XI0_12/d_5_ DECAP_INV_G11
XG6075 XI11_5/XI0/XI0_12/d__4_ XI11_5/XI0/XI0_12/d_4_ DECAP_INV_G11
XG6076 XI11_5/XI0/XI0_12/d__3_ XI11_5/XI0/XI0_12/d_3_ DECAP_INV_G11
XG6077 XI11_5/XI0/XI0_12/d__2_ XI11_5/XI0/XI0_12/d_2_ DECAP_INV_G11
XG6078 XI11_5/XI0/XI0_12/d__1_ XI11_5/XI0/XI0_12/d_1_ DECAP_INV_G11
XG6079 XI11_5/XI0/XI0_12/d__0_ XI11_5/XI0/XI0_12/d_0_ DECAP_INV_G11
XG6080 XI11_5/XI0/XI0_12/d_15_ XI11_5/XI0/XI0_12/d__15_ DECAP_INV_G11
XG6081 XI11_5/XI0/XI0_12/d_14_ XI11_5/XI0/XI0_12/d__14_ DECAP_INV_G11
XG6082 XI11_5/XI0/XI0_12/d_13_ XI11_5/XI0/XI0_12/d__13_ DECAP_INV_G11
XG6083 XI11_5/XI0/XI0_12/d_12_ XI11_5/XI0/XI0_12/d__12_ DECAP_INV_G11
XG6084 XI11_5/XI0/XI0_12/d_11_ XI11_5/XI0/XI0_12/d__11_ DECAP_INV_G11
XG6085 XI11_5/XI0/XI0_12/d_10_ XI11_5/XI0/XI0_12/d__10_ DECAP_INV_G11
XG6086 XI11_5/XI0/XI0_12/d_9_ XI11_5/XI0/XI0_12/d__9_ DECAP_INV_G11
XG6087 XI11_5/XI0/XI0_12/d_8_ XI11_5/XI0/XI0_12/d__8_ DECAP_INV_G11
XG6088 XI11_5/XI0/XI0_12/d_7_ XI11_5/XI0/XI0_12/d__7_ DECAP_INV_G11
XG6089 XI11_5/XI0/XI0_12/d_6_ XI11_5/XI0/XI0_12/d__6_ DECAP_INV_G11
XG6090 XI11_5/XI0/XI0_12/d_5_ XI11_5/XI0/XI0_12/d__5_ DECAP_INV_G11
XG6091 XI11_5/XI0/XI0_12/d_4_ XI11_5/XI0/XI0_12/d__4_ DECAP_INV_G11
XG6092 XI11_5/XI0/XI0_12/d_3_ XI11_5/XI0/XI0_12/d__3_ DECAP_INV_G11
XG6093 XI11_5/XI0/XI0_12/d_2_ XI11_5/XI0/XI0_12/d__2_ DECAP_INV_G11
XG6094 XI11_5/XI0/XI0_12/d_1_ XI11_5/XI0/XI0_12/d__1_ DECAP_INV_G11
XG6095 XI11_5/XI0/XI0_12/d_0_ XI11_5/XI0/XI0_12/d__0_ DECAP_INV_G11
XG6096 XI11_5/XI0/XI0_11/d__15_ XI11_5/XI0/XI0_11/d_15_ DECAP_INV_G11
XG6097 XI11_5/XI0/XI0_11/d__14_ XI11_5/XI0/XI0_11/d_14_ DECAP_INV_G11
XG6098 XI11_5/XI0/XI0_11/d__13_ XI11_5/XI0/XI0_11/d_13_ DECAP_INV_G11
XG6099 XI11_5/XI0/XI0_11/d__12_ XI11_5/XI0/XI0_11/d_12_ DECAP_INV_G11
XG6100 XI11_5/XI0/XI0_11/d__11_ XI11_5/XI0/XI0_11/d_11_ DECAP_INV_G11
XG6101 XI11_5/XI0/XI0_11/d__10_ XI11_5/XI0/XI0_11/d_10_ DECAP_INV_G11
XG6102 XI11_5/XI0/XI0_11/d__9_ XI11_5/XI0/XI0_11/d_9_ DECAP_INV_G11
XG6103 XI11_5/XI0/XI0_11/d__8_ XI11_5/XI0/XI0_11/d_8_ DECAP_INV_G11
XG6104 XI11_5/XI0/XI0_11/d__7_ XI11_5/XI0/XI0_11/d_7_ DECAP_INV_G11
XG6105 XI11_5/XI0/XI0_11/d__6_ XI11_5/XI0/XI0_11/d_6_ DECAP_INV_G11
XG6106 XI11_5/XI0/XI0_11/d__5_ XI11_5/XI0/XI0_11/d_5_ DECAP_INV_G11
XG6107 XI11_5/XI0/XI0_11/d__4_ XI11_5/XI0/XI0_11/d_4_ DECAP_INV_G11
XG6108 XI11_5/XI0/XI0_11/d__3_ XI11_5/XI0/XI0_11/d_3_ DECAP_INV_G11
XG6109 XI11_5/XI0/XI0_11/d__2_ XI11_5/XI0/XI0_11/d_2_ DECAP_INV_G11
XG6110 XI11_5/XI0/XI0_11/d__1_ XI11_5/XI0/XI0_11/d_1_ DECAP_INV_G11
XG6111 XI11_5/XI0/XI0_11/d__0_ XI11_5/XI0/XI0_11/d_0_ DECAP_INV_G11
XG6112 XI11_5/XI0/XI0_11/d_15_ XI11_5/XI0/XI0_11/d__15_ DECAP_INV_G11
XG6113 XI11_5/XI0/XI0_11/d_14_ XI11_5/XI0/XI0_11/d__14_ DECAP_INV_G11
XG6114 XI11_5/XI0/XI0_11/d_13_ XI11_5/XI0/XI0_11/d__13_ DECAP_INV_G11
XG6115 XI11_5/XI0/XI0_11/d_12_ XI11_5/XI0/XI0_11/d__12_ DECAP_INV_G11
XG6116 XI11_5/XI0/XI0_11/d_11_ XI11_5/XI0/XI0_11/d__11_ DECAP_INV_G11
XG6117 XI11_5/XI0/XI0_11/d_10_ XI11_5/XI0/XI0_11/d__10_ DECAP_INV_G11
XG6118 XI11_5/XI0/XI0_11/d_9_ XI11_5/XI0/XI0_11/d__9_ DECAP_INV_G11
XG6119 XI11_5/XI0/XI0_11/d_8_ XI11_5/XI0/XI0_11/d__8_ DECAP_INV_G11
XG6120 XI11_5/XI0/XI0_11/d_7_ XI11_5/XI0/XI0_11/d__7_ DECAP_INV_G11
XG6121 XI11_5/XI0/XI0_11/d_6_ XI11_5/XI0/XI0_11/d__6_ DECAP_INV_G11
XG6122 XI11_5/XI0/XI0_11/d_5_ XI11_5/XI0/XI0_11/d__5_ DECAP_INV_G11
XG6123 XI11_5/XI0/XI0_11/d_4_ XI11_5/XI0/XI0_11/d__4_ DECAP_INV_G11
XG6124 XI11_5/XI0/XI0_11/d_3_ XI11_5/XI0/XI0_11/d__3_ DECAP_INV_G11
XG6125 XI11_5/XI0/XI0_11/d_2_ XI11_5/XI0/XI0_11/d__2_ DECAP_INV_G11
XG6126 XI11_5/XI0/XI0_11/d_1_ XI11_5/XI0/XI0_11/d__1_ DECAP_INV_G11
XG6127 XI11_5/XI0/XI0_11/d_0_ XI11_5/XI0/XI0_11/d__0_ DECAP_INV_G11
XG6128 XI11_5/XI0/XI0_10/d__15_ XI11_5/XI0/XI0_10/d_15_ DECAP_INV_G11
XG6129 XI11_5/XI0/XI0_10/d__14_ XI11_5/XI0/XI0_10/d_14_ DECAP_INV_G11
XG6130 XI11_5/XI0/XI0_10/d__13_ XI11_5/XI0/XI0_10/d_13_ DECAP_INV_G11
XG6131 XI11_5/XI0/XI0_10/d__12_ XI11_5/XI0/XI0_10/d_12_ DECAP_INV_G11
XG6132 XI11_5/XI0/XI0_10/d__11_ XI11_5/XI0/XI0_10/d_11_ DECAP_INV_G11
XG6133 XI11_5/XI0/XI0_10/d__10_ XI11_5/XI0/XI0_10/d_10_ DECAP_INV_G11
XG6134 XI11_5/XI0/XI0_10/d__9_ XI11_5/XI0/XI0_10/d_9_ DECAP_INV_G11
XG6135 XI11_5/XI0/XI0_10/d__8_ XI11_5/XI0/XI0_10/d_8_ DECAP_INV_G11
XG6136 XI11_5/XI0/XI0_10/d__7_ XI11_5/XI0/XI0_10/d_7_ DECAP_INV_G11
XG6137 XI11_5/XI0/XI0_10/d__6_ XI11_5/XI0/XI0_10/d_6_ DECAP_INV_G11
XG6138 XI11_5/XI0/XI0_10/d__5_ XI11_5/XI0/XI0_10/d_5_ DECAP_INV_G11
XG6139 XI11_5/XI0/XI0_10/d__4_ XI11_5/XI0/XI0_10/d_4_ DECAP_INV_G11
XG6140 XI11_5/XI0/XI0_10/d__3_ XI11_5/XI0/XI0_10/d_3_ DECAP_INV_G11
XG6141 XI11_5/XI0/XI0_10/d__2_ XI11_5/XI0/XI0_10/d_2_ DECAP_INV_G11
XG6142 XI11_5/XI0/XI0_10/d__1_ XI11_5/XI0/XI0_10/d_1_ DECAP_INV_G11
XG6143 XI11_5/XI0/XI0_10/d__0_ XI11_5/XI0/XI0_10/d_0_ DECAP_INV_G11
XG6144 XI11_5/XI0/XI0_10/d_15_ XI11_5/XI0/XI0_10/d__15_ DECAP_INV_G11
XG6145 XI11_5/XI0/XI0_10/d_14_ XI11_5/XI0/XI0_10/d__14_ DECAP_INV_G11
XG6146 XI11_5/XI0/XI0_10/d_13_ XI11_5/XI0/XI0_10/d__13_ DECAP_INV_G11
XG6147 XI11_5/XI0/XI0_10/d_12_ XI11_5/XI0/XI0_10/d__12_ DECAP_INV_G11
XG6148 XI11_5/XI0/XI0_10/d_11_ XI11_5/XI0/XI0_10/d__11_ DECAP_INV_G11
XG6149 XI11_5/XI0/XI0_10/d_10_ XI11_5/XI0/XI0_10/d__10_ DECAP_INV_G11
XG6150 XI11_5/XI0/XI0_10/d_9_ XI11_5/XI0/XI0_10/d__9_ DECAP_INV_G11
XG6151 XI11_5/XI0/XI0_10/d_8_ XI11_5/XI0/XI0_10/d__8_ DECAP_INV_G11
XG6152 XI11_5/XI0/XI0_10/d_7_ XI11_5/XI0/XI0_10/d__7_ DECAP_INV_G11
XG6153 XI11_5/XI0/XI0_10/d_6_ XI11_5/XI0/XI0_10/d__6_ DECAP_INV_G11
XG6154 XI11_5/XI0/XI0_10/d_5_ XI11_5/XI0/XI0_10/d__5_ DECAP_INV_G11
XG6155 XI11_5/XI0/XI0_10/d_4_ XI11_5/XI0/XI0_10/d__4_ DECAP_INV_G11
XG6156 XI11_5/XI0/XI0_10/d_3_ XI11_5/XI0/XI0_10/d__3_ DECAP_INV_G11
XG6157 XI11_5/XI0/XI0_10/d_2_ XI11_5/XI0/XI0_10/d__2_ DECAP_INV_G11
XG6158 XI11_5/XI0/XI0_10/d_1_ XI11_5/XI0/XI0_10/d__1_ DECAP_INV_G11
XG6159 XI11_5/XI0/XI0_10/d_0_ XI11_5/XI0/XI0_10/d__0_ DECAP_INV_G11
XG6160 XI11_5/XI0/XI0_9/d__15_ XI11_5/XI0/XI0_9/d_15_ DECAP_INV_G11
XG6161 XI11_5/XI0/XI0_9/d__14_ XI11_5/XI0/XI0_9/d_14_ DECAP_INV_G11
XG6162 XI11_5/XI0/XI0_9/d__13_ XI11_5/XI0/XI0_9/d_13_ DECAP_INV_G11
XG6163 XI11_5/XI0/XI0_9/d__12_ XI11_5/XI0/XI0_9/d_12_ DECAP_INV_G11
XG6164 XI11_5/XI0/XI0_9/d__11_ XI11_5/XI0/XI0_9/d_11_ DECAP_INV_G11
XG6165 XI11_5/XI0/XI0_9/d__10_ XI11_5/XI0/XI0_9/d_10_ DECAP_INV_G11
XG6166 XI11_5/XI0/XI0_9/d__9_ XI11_5/XI0/XI0_9/d_9_ DECAP_INV_G11
XG6167 XI11_5/XI0/XI0_9/d__8_ XI11_5/XI0/XI0_9/d_8_ DECAP_INV_G11
XG6168 XI11_5/XI0/XI0_9/d__7_ XI11_5/XI0/XI0_9/d_7_ DECAP_INV_G11
XG6169 XI11_5/XI0/XI0_9/d__6_ XI11_5/XI0/XI0_9/d_6_ DECAP_INV_G11
XG6170 XI11_5/XI0/XI0_9/d__5_ XI11_5/XI0/XI0_9/d_5_ DECAP_INV_G11
XG6171 XI11_5/XI0/XI0_9/d__4_ XI11_5/XI0/XI0_9/d_4_ DECAP_INV_G11
XG6172 XI11_5/XI0/XI0_9/d__3_ XI11_5/XI0/XI0_9/d_3_ DECAP_INV_G11
XG6173 XI11_5/XI0/XI0_9/d__2_ XI11_5/XI0/XI0_9/d_2_ DECAP_INV_G11
XG6174 XI11_5/XI0/XI0_9/d__1_ XI11_5/XI0/XI0_9/d_1_ DECAP_INV_G11
XG6175 XI11_5/XI0/XI0_9/d__0_ XI11_5/XI0/XI0_9/d_0_ DECAP_INV_G11
XG6176 XI11_5/XI0/XI0_9/d_15_ XI11_5/XI0/XI0_9/d__15_ DECAP_INV_G11
XG6177 XI11_5/XI0/XI0_9/d_14_ XI11_5/XI0/XI0_9/d__14_ DECAP_INV_G11
XG6178 XI11_5/XI0/XI0_9/d_13_ XI11_5/XI0/XI0_9/d__13_ DECAP_INV_G11
XG6179 XI11_5/XI0/XI0_9/d_12_ XI11_5/XI0/XI0_9/d__12_ DECAP_INV_G11
XG6180 XI11_5/XI0/XI0_9/d_11_ XI11_5/XI0/XI0_9/d__11_ DECAP_INV_G11
XG6181 XI11_5/XI0/XI0_9/d_10_ XI11_5/XI0/XI0_9/d__10_ DECAP_INV_G11
XG6182 XI11_5/XI0/XI0_9/d_9_ XI11_5/XI0/XI0_9/d__9_ DECAP_INV_G11
XG6183 XI11_5/XI0/XI0_9/d_8_ XI11_5/XI0/XI0_9/d__8_ DECAP_INV_G11
XG6184 XI11_5/XI0/XI0_9/d_7_ XI11_5/XI0/XI0_9/d__7_ DECAP_INV_G11
XG6185 XI11_5/XI0/XI0_9/d_6_ XI11_5/XI0/XI0_9/d__6_ DECAP_INV_G11
XG6186 XI11_5/XI0/XI0_9/d_5_ XI11_5/XI0/XI0_9/d__5_ DECAP_INV_G11
XG6187 XI11_5/XI0/XI0_9/d_4_ XI11_5/XI0/XI0_9/d__4_ DECAP_INV_G11
XG6188 XI11_5/XI0/XI0_9/d_3_ XI11_5/XI0/XI0_9/d__3_ DECAP_INV_G11
XG6189 XI11_5/XI0/XI0_9/d_2_ XI11_5/XI0/XI0_9/d__2_ DECAP_INV_G11
XG6190 XI11_5/XI0/XI0_9/d_1_ XI11_5/XI0/XI0_9/d__1_ DECAP_INV_G11
XG6191 XI11_5/XI0/XI0_9/d_0_ XI11_5/XI0/XI0_9/d__0_ DECAP_INV_G11
XG6192 XI11_5/XI0/XI0_8/d__15_ XI11_5/XI0/XI0_8/d_15_ DECAP_INV_G11
XG6193 XI11_5/XI0/XI0_8/d__14_ XI11_5/XI0/XI0_8/d_14_ DECAP_INV_G11
XG6194 XI11_5/XI0/XI0_8/d__13_ XI11_5/XI0/XI0_8/d_13_ DECAP_INV_G11
XG6195 XI11_5/XI0/XI0_8/d__12_ XI11_5/XI0/XI0_8/d_12_ DECAP_INV_G11
XG6196 XI11_5/XI0/XI0_8/d__11_ XI11_5/XI0/XI0_8/d_11_ DECAP_INV_G11
XG6197 XI11_5/XI0/XI0_8/d__10_ XI11_5/XI0/XI0_8/d_10_ DECAP_INV_G11
XG6198 XI11_5/XI0/XI0_8/d__9_ XI11_5/XI0/XI0_8/d_9_ DECAP_INV_G11
XG6199 XI11_5/XI0/XI0_8/d__8_ XI11_5/XI0/XI0_8/d_8_ DECAP_INV_G11
XG6200 XI11_5/XI0/XI0_8/d__7_ XI11_5/XI0/XI0_8/d_7_ DECAP_INV_G11
XG6201 XI11_5/XI0/XI0_8/d__6_ XI11_5/XI0/XI0_8/d_6_ DECAP_INV_G11
XG6202 XI11_5/XI0/XI0_8/d__5_ XI11_5/XI0/XI0_8/d_5_ DECAP_INV_G11
XG6203 XI11_5/XI0/XI0_8/d__4_ XI11_5/XI0/XI0_8/d_4_ DECAP_INV_G11
XG6204 XI11_5/XI0/XI0_8/d__3_ XI11_5/XI0/XI0_8/d_3_ DECAP_INV_G11
XG6205 XI11_5/XI0/XI0_8/d__2_ XI11_5/XI0/XI0_8/d_2_ DECAP_INV_G11
XG6206 XI11_5/XI0/XI0_8/d__1_ XI11_5/XI0/XI0_8/d_1_ DECAP_INV_G11
XG6207 XI11_5/XI0/XI0_8/d__0_ XI11_5/XI0/XI0_8/d_0_ DECAP_INV_G11
XG6208 XI11_5/XI0/XI0_8/d_15_ XI11_5/XI0/XI0_8/d__15_ DECAP_INV_G11
XG6209 XI11_5/XI0/XI0_8/d_14_ XI11_5/XI0/XI0_8/d__14_ DECAP_INV_G11
XG6210 XI11_5/XI0/XI0_8/d_13_ XI11_5/XI0/XI0_8/d__13_ DECAP_INV_G11
XG6211 XI11_5/XI0/XI0_8/d_12_ XI11_5/XI0/XI0_8/d__12_ DECAP_INV_G11
XG6212 XI11_5/XI0/XI0_8/d_11_ XI11_5/XI0/XI0_8/d__11_ DECAP_INV_G11
XG6213 XI11_5/XI0/XI0_8/d_10_ XI11_5/XI0/XI0_8/d__10_ DECAP_INV_G11
XG6214 XI11_5/XI0/XI0_8/d_9_ XI11_5/XI0/XI0_8/d__9_ DECAP_INV_G11
XG6215 XI11_5/XI0/XI0_8/d_8_ XI11_5/XI0/XI0_8/d__8_ DECAP_INV_G11
XG6216 XI11_5/XI0/XI0_8/d_7_ XI11_5/XI0/XI0_8/d__7_ DECAP_INV_G11
XG6217 XI11_5/XI0/XI0_8/d_6_ XI11_5/XI0/XI0_8/d__6_ DECAP_INV_G11
XG6218 XI11_5/XI0/XI0_8/d_5_ XI11_5/XI0/XI0_8/d__5_ DECAP_INV_G11
XG6219 XI11_5/XI0/XI0_8/d_4_ XI11_5/XI0/XI0_8/d__4_ DECAP_INV_G11
XG6220 XI11_5/XI0/XI0_8/d_3_ XI11_5/XI0/XI0_8/d__3_ DECAP_INV_G11
XG6221 XI11_5/XI0/XI0_8/d_2_ XI11_5/XI0/XI0_8/d__2_ DECAP_INV_G11
XG6222 XI11_5/XI0/XI0_8/d_1_ XI11_5/XI0/XI0_8/d__1_ DECAP_INV_G11
XG6223 XI11_5/XI0/XI0_8/d_0_ XI11_5/XI0/XI0_8/d__0_ DECAP_INV_G11
XG6224 XI11_5/XI0/XI0_7/d__15_ XI11_5/XI0/XI0_7/d_15_ DECAP_INV_G11
XG6225 XI11_5/XI0/XI0_7/d__14_ XI11_5/XI0/XI0_7/d_14_ DECAP_INV_G11
XG6226 XI11_5/XI0/XI0_7/d__13_ XI11_5/XI0/XI0_7/d_13_ DECAP_INV_G11
XG6227 XI11_5/XI0/XI0_7/d__12_ XI11_5/XI0/XI0_7/d_12_ DECAP_INV_G11
XG6228 XI11_5/XI0/XI0_7/d__11_ XI11_5/XI0/XI0_7/d_11_ DECAP_INV_G11
XG6229 XI11_5/XI0/XI0_7/d__10_ XI11_5/XI0/XI0_7/d_10_ DECAP_INV_G11
XG6230 XI11_5/XI0/XI0_7/d__9_ XI11_5/XI0/XI0_7/d_9_ DECAP_INV_G11
XG6231 XI11_5/XI0/XI0_7/d__8_ XI11_5/XI0/XI0_7/d_8_ DECAP_INV_G11
XG6232 XI11_5/XI0/XI0_7/d__7_ XI11_5/XI0/XI0_7/d_7_ DECAP_INV_G11
XG6233 XI11_5/XI0/XI0_7/d__6_ XI11_5/XI0/XI0_7/d_6_ DECAP_INV_G11
XG6234 XI11_5/XI0/XI0_7/d__5_ XI11_5/XI0/XI0_7/d_5_ DECAP_INV_G11
XG6235 XI11_5/XI0/XI0_7/d__4_ XI11_5/XI0/XI0_7/d_4_ DECAP_INV_G11
XG6236 XI11_5/XI0/XI0_7/d__3_ XI11_5/XI0/XI0_7/d_3_ DECAP_INV_G11
XG6237 XI11_5/XI0/XI0_7/d__2_ XI11_5/XI0/XI0_7/d_2_ DECAP_INV_G11
XG6238 XI11_5/XI0/XI0_7/d__1_ XI11_5/XI0/XI0_7/d_1_ DECAP_INV_G11
XG6239 XI11_5/XI0/XI0_7/d__0_ XI11_5/XI0/XI0_7/d_0_ DECAP_INV_G11
XG6240 XI11_5/XI0/XI0_7/d_15_ XI11_5/XI0/XI0_7/d__15_ DECAP_INV_G11
XG6241 XI11_5/XI0/XI0_7/d_14_ XI11_5/XI0/XI0_7/d__14_ DECAP_INV_G11
XG6242 XI11_5/XI0/XI0_7/d_13_ XI11_5/XI0/XI0_7/d__13_ DECAP_INV_G11
XG6243 XI11_5/XI0/XI0_7/d_12_ XI11_5/XI0/XI0_7/d__12_ DECAP_INV_G11
XG6244 XI11_5/XI0/XI0_7/d_11_ XI11_5/XI0/XI0_7/d__11_ DECAP_INV_G11
XG6245 XI11_5/XI0/XI0_7/d_10_ XI11_5/XI0/XI0_7/d__10_ DECAP_INV_G11
XG6246 XI11_5/XI0/XI0_7/d_9_ XI11_5/XI0/XI0_7/d__9_ DECAP_INV_G11
XG6247 XI11_5/XI0/XI0_7/d_8_ XI11_5/XI0/XI0_7/d__8_ DECAP_INV_G11
XG6248 XI11_5/XI0/XI0_7/d_7_ XI11_5/XI0/XI0_7/d__7_ DECAP_INV_G11
XG6249 XI11_5/XI0/XI0_7/d_6_ XI11_5/XI0/XI0_7/d__6_ DECAP_INV_G11
XG6250 XI11_5/XI0/XI0_7/d_5_ XI11_5/XI0/XI0_7/d__5_ DECAP_INV_G11
XG6251 XI11_5/XI0/XI0_7/d_4_ XI11_5/XI0/XI0_7/d__4_ DECAP_INV_G11
XG6252 XI11_5/XI0/XI0_7/d_3_ XI11_5/XI0/XI0_7/d__3_ DECAP_INV_G11
XG6253 XI11_5/XI0/XI0_7/d_2_ XI11_5/XI0/XI0_7/d__2_ DECAP_INV_G11
XG6254 XI11_5/XI0/XI0_7/d_1_ XI11_5/XI0/XI0_7/d__1_ DECAP_INV_G11
XG6255 XI11_5/XI0/XI0_7/d_0_ XI11_5/XI0/XI0_7/d__0_ DECAP_INV_G11
XG6256 XI11_5/XI0/XI0_6/d__15_ XI11_5/XI0/XI0_6/d_15_ DECAP_INV_G11
XG6257 XI11_5/XI0/XI0_6/d__14_ XI11_5/XI0/XI0_6/d_14_ DECAP_INV_G11
XG6258 XI11_5/XI0/XI0_6/d__13_ XI11_5/XI0/XI0_6/d_13_ DECAP_INV_G11
XG6259 XI11_5/XI0/XI0_6/d__12_ XI11_5/XI0/XI0_6/d_12_ DECAP_INV_G11
XG6260 XI11_5/XI0/XI0_6/d__11_ XI11_5/XI0/XI0_6/d_11_ DECAP_INV_G11
XG6261 XI11_5/XI0/XI0_6/d__10_ XI11_5/XI0/XI0_6/d_10_ DECAP_INV_G11
XG6262 XI11_5/XI0/XI0_6/d__9_ XI11_5/XI0/XI0_6/d_9_ DECAP_INV_G11
XG6263 XI11_5/XI0/XI0_6/d__8_ XI11_5/XI0/XI0_6/d_8_ DECAP_INV_G11
XG6264 XI11_5/XI0/XI0_6/d__7_ XI11_5/XI0/XI0_6/d_7_ DECAP_INV_G11
XG6265 XI11_5/XI0/XI0_6/d__6_ XI11_5/XI0/XI0_6/d_6_ DECAP_INV_G11
XG6266 XI11_5/XI0/XI0_6/d__5_ XI11_5/XI0/XI0_6/d_5_ DECAP_INV_G11
XG6267 XI11_5/XI0/XI0_6/d__4_ XI11_5/XI0/XI0_6/d_4_ DECAP_INV_G11
XG6268 XI11_5/XI0/XI0_6/d__3_ XI11_5/XI0/XI0_6/d_3_ DECAP_INV_G11
XG6269 XI11_5/XI0/XI0_6/d__2_ XI11_5/XI0/XI0_6/d_2_ DECAP_INV_G11
XG6270 XI11_5/XI0/XI0_6/d__1_ XI11_5/XI0/XI0_6/d_1_ DECAP_INV_G11
XG6271 XI11_5/XI0/XI0_6/d__0_ XI11_5/XI0/XI0_6/d_0_ DECAP_INV_G11
XG6272 XI11_5/XI0/XI0_6/d_15_ XI11_5/XI0/XI0_6/d__15_ DECAP_INV_G11
XG6273 XI11_5/XI0/XI0_6/d_14_ XI11_5/XI0/XI0_6/d__14_ DECAP_INV_G11
XG6274 XI11_5/XI0/XI0_6/d_13_ XI11_5/XI0/XI0_6/d__13_ DECAP_INV_G11
XG6275 XI11_5/XI0/XI0_6/d_12_ XI11_5/XI0/XI0_6/d__12_ DECAP_INV_G11
XG6276 XI11_5/XI0/XI0_6/d_11_ XI11_5/XI0/XI0_6/d__11_ DECAP_INV_G11
XG6277 XI11_5/XI0/XI0_6/d_10_ XI11_5/XI0/XI0_6/d__10_ DECAP_INV_G11
XG6278 XI11_5/XI0/XI0_6/d_9_ XI11_5/XI0/XI0_6/d__9_ DECAP_INV_G11
XG6279 XI11_5/XI0/XI0_6/d_8_ XI11_5/XI0/XI0_6/d__8_ DECAP_INV_G11
XG6280 XI11_5/XI0/XI0_6/d_7_ XI11_5/XI0/XI0_6/d__7_ DECAP_INV_G11
XG6281 XI11_5/XI0/XI0_6/d_6_ XI11_5/XI0/XI0_6/d__6_ DECAP_INV_G11
XG6282 XI11_5/XI0/XI0_6/d_5_ XI11_5/XI0/XI0_6/d__5_ DECAP_INV_G11
XG6283 XI11_5/XI0/XI0_6/d_4_ XI11_5/XI0/XI0_6/d__4_ DECAP_INV_G11
XG6284 XI11_5/XI0/XI0_6/d_3_ XI11_5/XI0/XI0_6/d__3_ DECAP_INV_G11
XG6285 XI11_5/XI0/XI0_6/d_2_ XI11_5/XI0/XI0_6/d__2_ DECAP_INV_G11
XG6286 XI11_5/XI0/XI0_6/d_1_ XI11_5/XI0/XI0_6/d__1_ DECAP_INV_G11
XG6287 XI11_5/XI0/XI0_6/d_0_ XI11_5/XI0/XI0_6/d__0_ DECAP_INV_G11
XG6288 XI11_5/XI0/XI0_5/d__15_ XI11_5/XI0/XI0_5/d_15_ DECAP_INV_G11
XG6289 XI11_5/XI0/XI0_5/d__14_ XI11_5/XI0/XI0_5/d_14_ DECAP_INV_G11
XG6290 XI11_5/XI0/XI0_5/d__13_ XI11_5/XI0/XI0_5/d_13_ DECAP_INV_G11
XG6291 XI11_5/XI0/XI0_5/d__12_ XI11_5/XI0/XI0_5/d_12_ DECAP_INV_G11
XG6292 XI11_5/XI0/XI0_5/d__11_ XI11_5/XI0/XI0_5/d_11_ DECAP_INV_G11
XG6293 XI11_5/XI0/XI0_5/d__10_ XI11_5/XI0/XI0_5/d_10_ DECAP_INV_G11
XG6294 XI11_5/XI0/XI0_5/d__9_ XI11_5/XI0/XI0_5/d_9_ DECAP_INV_G11
XG6295 XI11_5/XI0/XI0_5/d__8_ XI11_5/XI0/XI0_5/d_8_ DECAP_INV_G11
XG6296 XI11_5/XI0/XI0_5/d__7_ XI11_5/XI0/XI0_5/d_7_ DECAP_INV_G11
XG6297 XI11_5/XI0/XI0_5/d__6_ XI11_5/XI0/XI0_5/d_6_ DECAP_INV_G11
XG6298 XI11_5/XI0/XI0_5/d__5_ XI11_5/XI0/XI0_5/d_5_ DECAP_INV_G11
XG6299 XI11_5/XI0/XI0_5/d__4_ XI11_5/XI0/XI0_5/d_4_ DECAP_INV_G11
XG6300 XI11_5/XI0/XI0_5/d__3_ XI11_5/XI0/XI0_5/d_3_ DECAP_INV_G11
XG6301 XI11_5/XI0/XI0_5/d__2_ XI11_5/XI0/XI0_5/d_2_ DECAP_INV_G11
XG6302 XI11_5/XI0/XI0_5/d__1_ XI11_5/XI0/XI0_5/d_1_ DECAP_INV_G11
XG6303 XI11_5/XI0/XI0_5/d__0_ XI11_5/XI0/XI0_5/d_0_ DECAP_INV_G11
XG6304 XI11_5/XI0/XI0_5/d_15_ XI11_5/XI0/XI0_5/d__15_ DECAP_INV_G11
XG6305 XI11_5/XI0/XI0_5/d_14_ XI11_5/XI0/XI0_5/d__14_ DECAP_INV_G11
XG6306 XI11_5/XI0/XI0_5/d_13_ XI11_5/XI0/XI0_5/d__13_ DECAP_INV_G11
XG6307 XI11_5/XI0/XI0_5/d_12_ XI11_5/XI0/XI0_5/d__12_ DECAP_INV_G11
XG6308 XI11_5/XI0/XI0_5/d_11_ XI11_5/XI0/XI0_5/d__11_ DECAP_INV_G11
XG6309 XI11_5/XI0/XI0_5/d_10_ XI11_5/XI0/XI0_5/d__10_ DECAP_INV_G11
XG6310 XI11_5/XI0/XI0_5/d_9_ XI11_5/XI0/XI0_5/d__9_ DECAP_INV_G11
XG6311 XI11_5/XI0/XI0_5/d_8_ XI11_5/XI0/XI0_5/d__8_ DECAP_INV_G11
XG6312 XI11_5/XI0/XI0_5/d_7_ XI11_5/XI0/XI0_5/d__7_ DECAP_INV_G11
XG6313 XI11_5/XI0/XI0_5/d_6_ XI11_5/XI0/XI0_5/d__6_ DECAP_INV_G11
XG6314 XI11_5/XI0/XI0_5/d_5_ XI11_5/XI0/XI0_5/d__5_ DECAP_INV_G11
XG6315 XI11_5/XI0/XI0_5/d_4_ XI11_5/XI0/XI0_5/d__4_ DECAP_INV_G11
XG6316 XI11_5/XI0/XI0_5/d_3_ XI11_5/XI0/XI0_5/d__3_ DECAP_INV_G11
XG6317 XI11_5/XI0/XI0_5/d_2_ XI11_5/XI0/XI0_5/d__2_ DECAP_INV_G11
XG6318 XI11_5/XI0/XI0_5/d_1_ XI11_5/XI0/XI0_5/d__1_ DECAP_INV_G11
XG6319 XI11_5/XI0/XI0_5/d_0_ XI11_5/XI0/XI0_5/d__0_ DECAP_INV_G11
XG6320 XI11_5/XI0/XI0_4/d__15_ XI11_5/XI0/XI0_4/d_15_ DECAP_INV_G11
XG6321 XI11_5/XI0/XI0_4/d__14_ XI11_5/XI0/XI0_4/d_14_ DECAP_INV_G11
XG6322 XI11_5/XI0/XI0_4/d__13_ XI11_5/XI0/XI0_4/d_13_ DECAP_INV_G11
XG6323 XI11_5/XI0/XI0_4/d__12_ XI11_5/XI0/XI0_4/d_12_ DECAP_INV_G11
XG6324 XI11_5/XI0/XI0_4/d__11_ XI11_5/XI0/XI0_4/d_11_ DECAP_INV_G11
XG6325 XI11_5/XI0/XI0_4/d__10_ XI11_5/XI0/XI0_4/d_10_ DECAP_INV_G11
XG6326 XI11_5/XI0/XI0_4/d__9_ XI11_5/XI0/XI0_4/d_9_ DECAP_INV_G11
XG6327 XI11_5/XI0/XI0_4/d__8_ XI11_5/XI0/XI0_4/d_8_ DECAP_INV_G11
XG6328 XI11_5/XI0/XI0_4/d__7_ XI11_5/XI0/XI0_4/d_7_ DECAP_INV_G11
XG6329 XI11_5/XI0/XI0_4/d__6_ XI11_5/XI0/XI0_4/d_6_ DECAP_INV_G11
XG6330 XI11_5/XI0/XI0_4/d__5_ XI11_5/XI0/XI0_4/d_5_ DECAP_INV_G11
XG6331 XI11_5/XI0/XI0_4/d__4_ XI11_5/XI0/XI0_4/d_4_ DECAP_INV_G11
XG6332 XI11_5/XI0/XI0_4/d__3_ XI11_5/XI0/XI0_4/d_3_ DECAP_INV_G11
XG6333 XI11_5/XI0/XI0_4/d__2_ XI11_5/XI0/XI0_4/d_2_ DECAP_INV_G11
XG6334 XI11_5/XI0/XI0_4/d__1_ XI11_5/XI0/XI0_4/d_1_ DECAP_INV_G11
XG6335 XI11_5/XI0/XI0_4/d__0_ XI11_5/XI0/XI0_4/d_0_ DECAP_INV_G11
XG6336 XI11_5/XI0/XI0_4/d_15_ XI11_5/XI0/XI0_4/d__15_ DECAP_INV_G11
XG6337 XI11_5/XI0/XI0_4/d_14_ XI11_5/XI0/XI0_4/d__14_ DECAP_INV_G11
XG6338 XI11_5/XI0/XI0_4/d_13_ XI11_5/XI0/XI0_4/d__13_ DECAP_INV_G11
XG6339 XI11_5/XI0/XI0_4/d_12_ XI11_5/XI0/XI0_4/d__12_ DECAP_INV_G11
XG6340 XI11_5/XI0/XI0_4/d_11_ XI11_5/XI0/XI0_4/d__11_ DECAP_INV_G11
XG6341 XI11_5/XI0/XI0_4/d_10_ XI11_5/XI0/XI0_4/d__10_ DECAP_INV_G11
XG6342 XI11_5/XI0/XI0_4/d_9_ XI11_5/XI0/XI0_4/d__9_ DECAP_INV_G11
XG6343 XI11_5/XI0/XI0_4/d_8_ XI11_5/XI0/XI0_4/d__8_ DECAP_INV_G11
XG6344 XI11_5/XI0/XI0_4/d_7_ XI11_5/XI0/XI0_4/d__7_ DECAP_INV_G11
XG6345 XI11_5/XI0/XI0_4/d_6_ XI11_5/XI0/XI0_4/d__6_ DECAP_INV_G11
XG6346 XI11_5/XI0/XI0_4/d_5_ XI11_5/XI0/XI0_4/d__5_ DECAP_INV_G11
XG6347 XI11_5/XI0/XI0_4/d_4_ XI11_5/XI0/XI0_4/d__4_ DECAP_INV_G11
XG6348 XI11_5/XI0/XI0_4/d_3_ XI11_5/XI0/XI0_4/d__3_ DECAP_INV_G11
XG6349 XI11_5/XI0/XI0_4/d_2_ XI11_5/XI0/XI0_4/d__2_ DECAP_INV_G11
XG6350 XI11_5/XI0/XI0_4/d_1_ XI11_5/XI0/XI0_4/d__1_ DECAP_INV_G11
XG6351 XI11_5/XI0/XI0_4/d_0_ XI11_5/XI0/XI0_4/d__0_ DECAP_INV_G11
XG6352 XI11_5/XI0/XI0_3/d__15_ XI11_5/XI0/XI0_3/d_15_ DECAP_INV_G11
XG6353 XI11_5/XI0/XI0_3/d__14_ XI11_5/XI0/XI0_3/d_14_ DECAP_INV_G11
XG6354 XI11_5/XI0/XI0_3/d__13_ XI11_5/XI0/XI0_3/d_13_ DECAP_INV_G11
XG6355 XI11_5/XI0/XI0_3/d__12_ XI11_5/XI0/XI0_3/d_12_ DECAP_INV_G11
XG6356 XI11_5/XI0/XI0_3/d__11_ XI11_5/XI0/XI0_3/d_11_ DECAP_INV_G11
XG6357 XI11_5/XI0/XI0_3/d__10_ XI11_5/XI0/XI0_3/d_10_ DECAP_INV_G11
XG6358 XI11_5/XI0/XI0_3/d__9_ XI11_5/XI0/XI0_3/d_9_ DECAP_INV_G11
XG6359 XI11_5/XI0/XI0_3/d__8_ XI11_5/XI0/XI0_3/d_8_ DECAP_INV_G11
XG6360 XI11_5/XI0/XI0_3/d__7_ XI11_5/XI0/XI0_3/d_7_ DECAP_INV_G11
XG6361 XI11_5/XI0/XI0_3/d__6_ XI11_5/XI0/XI0_3/d_6_ DECAP_INV_G11
XG6362 XI11_5/XI0/XI0_3/d__5_ XI11_5/XI0/XI0_3/d_5_ DECAP_INV_G11
XG6363 XI11_5/XI0/XI0_3/d__4_ XI11_5/XI0/XI0_3/d_4_ DECAP_INV_G11
XG6364 XI11_5/XI0/XI0_3/d__3_ XI11_5/XI0/XI0_3/d_3_ DECAP_INV_G11
XG6365 XI11_5/XI0/XI0_3/d__2_ XI11_5/XI0/XI0_3/d_2_ DECAP_INV_G11
XG6366 XI11_5/XI0/XI0_3/d__1_ XI11_5/XI0/XI0_3/d_1_ DECAP_INV_G11
XG6367 XI11_5/XI0/XI0_3/d__0_ XI11_5/XI0/XI0_3/d_0_ DECAP_INV_G11
XG6368 XI11_5/XI0/XI0_3/d_15_ XI11_5/XI0/XI0_3/d__15_ DECAP_INV_G11
XG6369 XI11_5/XI0/XI0_3/d_14_ XI11_5/XI0/XI0_3/d__14_ DECAP_INV_G11
XG6370 XI11_5/XI0/XI0_3/d_13_ XI11_5/XI0/XI0_3/d__13_ DECAP_INV_G11
XG6371 XI11_5/XI0/XI0_3/d_12_ XI11_5/XI0/XI0_3/d__12_ DECAP_INV_G11
XG6372 XI11_5/XI0/XI0_3/d_11_ XI11_5/XI0/XI0_3/d__11_ DECAP_INV_G11
XG6373 XI11_5/XI0/XI0_3/d_10_ XI11_5/XI0/XI0_3/d__10_ DECAP_INV_G11
XG6374 XI11_5/XI0/XI0_3/d_9_ XI11_5/XI0/XI0_3/d__9_ DECAP_INV_G11
XG6375 XI11_5/XI0/XI0_3/d_8_ XI11_5/XI0/XI0_3/d__8_ DECAP_INV_G11
XG6376 XI11_5/XI0/XI0_3/d_7_ XI11_5/XI0/XI0_3/d__7_ DECAP_INV_G11
XG6377 XI11_5/XI0/XI0_3/d_6_ XI11_5/XI0/XI0_3/d__6_ DECAP_INV_G11
XG6378 XI11_5/XI0/XI0_3/d_5_ XI11_5/XI0/XI0_3/d__5_ DECAP_INV_G11
XG6379 XI11_5/XI0/XI0_3/d_4_ XI11_5/XI0/XI0_3/d__4_ DECAP_INV_G11
XG6380 XI11_5/XI0/XI0_3/d_3_ XI11_5/XI0/XI0_3/d__3_ DECAP_INV_G11
XG6381 XI11_5/XI0/XI0_3/d_2_ XI11_5/XI0/XI0_3/d__2_ DECAP_INV_G11
XG6382 XI11_5/XI0/XI0_3/d_1_ XI11_5/XI0/XI0_3/d__1_ DECAP_INV_G11
XG6383 XI11_5/XI0/XI0_3/d_0_ XI11_5/XI0/XI0_3/d__0_ DECAP_INV_G11
XG6384 XI11_5/XI0/XI0_2/d__15_ XI11_5/XI0/XI0_2/d_15_ DECAP_INV_G11
XG6385 XI11_5/XI0/XI0_2/d__14_ XI11_5/XI0/XI0_2/d_14_ DECAP_INV_G11
XG6386 XI11_5/XI0/XI0_2/d__13_ XI11_5/XI0/XI0_2/d_13_ DECAP_INV_G11
XG6387 XI11_5/XI0/XI0_2/d__12_ XI11_5/XI0/XI0_2/d_12_ DECAP_INV_G11
XG6388 XI11_5/XI0/XI0_2/d__11_ XI11_5/XI0/XI0_2/d_11_ DECAP_INV_G11
XG6389 XI11_5/XI0/XI0_2/d__10_ XI11_5/XI0/XI0_2/d_10_ DECAP_INV_G11
XG6390 XI11_5/XI0/XI0_2/d__9_ XI11_5/XI0/XI0_2/d_9_ DECAP_INV_G11
XG6391 XI11_5/XI0/XI0_2/d__8_ XI11_5/XI0/XI0_2/d_8_ DECAP_INV_G11
XG6392 XI11_5/XI0/XI0_2/d__7_ XI11_5/XI0/XI0_2/d_7_ DECAP_INV_G11
XG6393 XI11_5/XI0/XI0_2/d__6_ XI11_5/XI0/XI0_2/d_6_ DECAP_INV_G11
XG6394 XI11_5/XI0/XI0_2/d__5_ XI11_5/XI0/XI0_2/d_5_ DECAP_INV_G11
XG6395 XI11_5/XI0/XI0_2/d__4_ XI11_5/XI0/XI0_2/d_4_ DECAP_INV_G11
XG6396 XI11_5/XI0/XI0_2/d__3_ XI11_5/XI0/XI0_2/d_3_ DECAP_INV_G11
XG6397 XI11_5/XI0/XI0_2/d__2_ XI11_5/XI0/XI0_2/d_2_ DECAP_INV_G11
XG6398 XI11_5/XI0/XI0_2/d__1_ XI11_5/XI0/XI0_2/d_1_ DECAP_INV_G11
XG6399 XI11_5/XI0/XI0_2/d__0_ XI11_5/XI0/XI0_2/d_0_ DECAP_INV_G11
XG6400 XI11_5/XI0/XI0_2/d_15_ XI11_5/XI0/XI0_2/d__15_ DECAP_INV_G11
XG6401 XI11_5/XI0/XI0_2/d_14_ XI11_5/XI0/XI0_2/d__14_ DECAP_INV_G11
XG6402 XI11_5/XI0/XI0_2/d_13_ XI11_5/XI0/XI0_2/d__13_ DECAP_INV_G11
XG6403 XI11_5/XI0/XI0_2/d_12_ XI11_5/XI0/XI0_2/d__12_ DECAP_INV_G11
XG6404 XI11_5/XI0/XI0_2/d_11_ XI11_5/XI0/XI0_2/d__11_ DECAP_INV_G11
XG6405 XI11_5/XI0/XI0_2/d_10_ XI11_5/XI0/XI0_2/d__10_ DECAP_INV_G11
XG6406 XI11_5/XI0/XI0_2/d_9_ XI11_5/XI0/XI0_2/d__9_ DECAP_INV_G11
XG6407 XI11_5/XI0/XI0_2/d_8_ XI11_5/XI0/XI0_2/d__8_ DECAP_INV_G11
XG6408 XI11_5/XI0/XI0_2/d_7_ XI11_5/XI0/XI0_2/d__7_ DECAP_INV_G11
XG6409 XI11_5/XI0/XI0_2/d_6_ XI11_5/XI0/XI0_2/d__6_ DECAP_INV_G11
XG6410 XI11_5/XI0/XI0_2/d_5_ XI11_5/XI0/XI0_2/d__5_ DECAP_INV_G11
XG6411 XI11_5/XI0/XI0_2/d_4_ XI11_5/XI0/XI0_2/d__4_ DECAP_INV_G11
XG6412 XI11_5/XI0/XI0_2/d_3_ XI11_5/XI0/XI0_2/d__3_ DECAP_INV_G11
XG6413 XI11_5/XI0/XI0_2/d_2_ XI11_5/XI0/XI0_2/d__2_ DECAP_INV_G11
XG6414 XI11_5/XI0/XI0_2/d_1_ XI11_5/XI0/XI0_2/d__1_ DECAP_INV_G11
XG6415 XI11_5/XI0/XI0_2/d_0_ XI11_5/XI0/XI0_2/d__0_ DECAP_INV_G11
XG6416 XI11_5/XI0/XI0_1/d__15_ XI11_5/XI0/XI0_1/d_15_ DECAP_INV_G11
XG6417 XI11_5/XI0/XI0_1/d__14_ XI11_5/XI0/XI0_1/d_14_ DECAP_INV_G11
XG6418 XI11_5/XI0/XI0_1/d__13_ XI11_5/XI0/XI0_1/d_13_ DECAP_INV_G11
XG6419 XI11_5/XI0/XI0_1/d__12_ XI11_5/XI0/XI0_1/d_12_ DECAP_INV_G11
XG6420 XI11_5/XI0/XI0_1/d__11_ XI11_5/XI0/XI0_1/d_11_ DECAP_INV_G11
XG6421 XI11_5/XI0/XI0_1/d__10_ XI11_5/XI0/XI0_1/d_10_ DECAP_INV_G11
XG6422 XI11_5/XI0/XI0_1/d__9_ XI11_5/XI0/XI0_1/d_9_ DECAP_INV_G11
XG6423 XI11_5/XI0/XI0_1/d__8_ XI11_5/XI0/XI0_1/d_8_ DECAP_INV_G11
XG6424 XI11_5/XI0/XI0_1/d__7_ XI11_5/XI0/XI0_1/d_7_ DECAP_INV_G11
XG6425 XI11_5/XI0/XI0_1/d__6_ XI11_5/XI0/XI0_1/d_6_ DECAP_INV_G11
XG6426 XI11_5/XI0/XI0_1/d__5_ XI11_5/XI0/XI0_1/d_5_ DECAP_INV_G11
XG6427 XI11_5/XI0/XI0_1/d__4_ XI11_5/XI0/XI0_1/d_4_ DECAP_INV_G11
XG6428 XI11_5/XI0/XI0_1/d__3_ XI11_5/XI0/XI0_1/d_3_ DECAP_INV_G11
XG6429 XI11_5/XI0/XI0_1/d__2_ XI11_5/XI0/XI0_1/d_2_ DECAP_INV_G11
XG6430 XI11_5/XI0/XI0_1/d__1_ XI11_5/XI0/XI0_1/d_1_ DECAP_INV_G11
XG6431 XI11_5/XI0/XI0_1/d__0_ XI11_5/XI0/XI0_1/d_0_ DECAP_INV_G11
XG6432 XI11_5/XI0/XI0_1/d_15_ XI11_5/XI0/XI0_1/d__15_ DECAP_INV_G11
XG6433 XI11_5/XI0/XI0_1/d_14_ XI11_5/XI0/XI0_1/d__14_ DECAP_INV_G11
XG6434 XI11_5/XI0/XI0_1/d_13_ XI11_5/XI0/XI0_1/d__13_ DECAP_INV_G11
XG6435 XI11_5/XI0/XI0_1/d_12_ XI11_5/XI0/XI0_1/d__12_ DECAP_INV_G11
XG6436 XI11_5/XI0/XI0_1/d_11_ XI11_5/XI0/XI0_1/d__11_ DECAP_INV_G11
XG6437 XI11_5/XI0/XI0_1/d_10_ XI11_5/XI0/XI0_1/d__10_ DECAP_INV_G11
XG6438 XI11_5/XI0/XI0_1/d_9_ XI11_5/XI0/XI0_1/d__9_ DECAP_INV_G11
XG6439 XI11_5/XI0/XI0_1/d_8_ XI11_5/XI0/XI0_1/d__8_ DECAP_INV_G11
XG6440 XI11_5/XI0/XI0_1/d_7_ XI11_5/XI0/XI0_1/d__7_ DECAP_INV_G11
XG6441 XI11_5/XI0/XI0_1/d_6_ XI11_5/XI0/XI0_1/d__6_ DECAP_INV_G11
XG6442 XI11_5/XI0/XI0_1/d_5_ XI11_5/XI0/XI0_1/d__5_ DECAP_INV_G11
XG6443 XI11_5/XI0/XI0_1/d_4_ XI11_5/XI0/XI0_1/d__4_ DECAP_INV_G11
XG6444 XI11_5/XI0/XI0_1/d_3_ XI11_5/XI0/XI0_1/d__3_ DECAP_INV_G11
XG6445 XI11_5/XI0/XI0_1/d_2_ XI11_5/XI0/XI0_1/d__2_ DECAP_INV_G11
XG6446 XI11_5/XI0/XI0_1/d_1_ XI11_5/XI0/XI0_1/d__1_ DECAP_INV_G11
XG6447 XI11_5/XI0/XI0_1/d_0_ XI11_5/XI0/XI0_1/d__0_ DECAP_INV_G11
XG6448 XI11_5/XI0/XI0_0/d__15_ XI11_5/XI0/XI0_0/d_15_ DECAP_INV_G11
XG6449 XI11_5/XI0/XI0_0/d__14_ XI11_5/XI0/XI0_0/d_14_ DECAP_INV_G11
XG6450 XI11_5/XI0/XI0_0/d__13_ XI11_5/XI0/XI0_0/d_13_ DECAP_INV_G11
XG6451 XI11_5/XI0/XI0_0/d__12_ XI11_5/XI0/XI0_0/d_12_ DECAP_INV_G11
XG6452 XI11_5/XI0/XI0_0/d__11_ XI11_5/XI0/XI0_0/d_11_ DECAP_INV_G11
XG6453 XI11_5/XI0/XI0_0/d__10_ XI11_5/XI0/XI0_0/d_10_ DECAP_INV_G11
XG6454 XI11_5/XI0/XI0_0/d__9_ XI11_5/XI0/XI0_0/d_9_ DECAP_INV_G11
XG6455 XI11_5/XI0/XI0_0/d__8_ XI11_5/XI0/XI0_0/d_8_ DECAP_INV_G11
XG6456 XI11_5/XI0/XI0_0/d__7_ XI11_5/XI0/XI0_0/d_7_ DECAP_INV_G11
XG6457 XI11_5/XI0/XI0_0/d__6_ XI11_5/XI0/XI0_0/d_6_ DECAP_INV_G11
XG6458 XI11_5/XI0/XI0_0/d__5_ XI11_5/XI0/XI0_0/d_5_ DECAP_INV_G11
XG6459 XI11_5/XI0/XI0_0/d__4_ XI11_5/XI0/XI0_0/d_4_ DECAP_INV_G11
XG6460 XI11_5/XI0/XI0_0/d__3_ XI11_5/XI0/XI0_0/d_3_ DECAP_INV_G11
XG6461 XI11_5/XI0/XI0_0/d__2_ XI11_5/XI0/XI0_0/d_2_ DECAP_INV_G11
XG6462 XI11_5/XI0/XI0_0/d__1_ XI11_5/XI0/XI0_0/d_1_ DECAP_INV_G11
XG6463 XI11_5/XI0/XI0_0/d__0_ XI11_5/XI0/XI0_0/d_0_ DECAP_INV_G11
XG6464 XI11_5/XI0/XI0_0/d_15_ XI11_5/XI0/XI0_0/d__15_ DECAP_INV_G11
XG6465 XI11_5/XI0/XI0_0/d_14_ XI11_5/XI0/XI0_0/d__14_ DECAP_INV_G11
XG6466 XI11_5/XI0/XI0_0/d_13_ XI11_5/XI0/XI0_0/d__13_ DECAP_INV_G11
XG6467 XI11_5/XI0/XI0_0/d_12_ XI11_5/XI0/XI0_0/d__12_ DECAP_INV_G11
XG6468 XI11_5/XI0/XI0_0/d_11_ XI11_5/XI0/XI0_0/d__11_ DECAP_INV_G11
XG6469 XI11_5/XI0/XI0_0/d_10_ XI11_5/XI0/XI0_0/d__10_ DECAP_INV_G11
XG6470 XI11_5/XI0/XI0_0/d_9_ XI11_5/XI0/XI0_0/d__9_ DECAP_INV_G11
XG6471 XI11_5/XI0/XI0_0/d_8_ XI11_5/XI0/XI0_0/d__8_ DECAP_INV_G11
XG6472 XI11_5/XI0/XI0_0/d_7_ XI11_5/XI0/XI0_0/d__7_ DECAP_INV_G11
XG6473 XI11_5/XI0/XI0_0/d_6_ XI11_5/XI0/XI0_0/d__6_ DECAP_INV_G11
XG6474 XI11_5/XI0/XI0_0/d_5_ XI11_5/XI0/XI0_0/d__5_ DECAP_INV_G11
XG6475 XI11_5/XI0/XI0_0/d_4_ XI11_5/XI0/XI0_0/d__4_ DECAP_INV_G11
XG6476 XI11_5/XI0/XI0_0/d_3_ XI11_5/XI0/XI0_0/d__3_ DECAP_INV_G11
XG6477 XI11_5/XI0/XI0_0/d_2_ XI11_5/XI0/XI0_0/d__2_ DECAP_INV_G11
XG6478 XI11_5/XI0/XI0_0/d_1_ XI11_5/XI0/XI0_0/d__1_ DECAP_INV_G11
XG6479 XI11_5/XI0/XI0_0/d_0_ XI11_5/XI0/XI0_0/d__0_ DECAP_INV_G11
XG6480 XI11_4/XI3/net17 XI11_4/XI3/net5 DECAP_INV_G7
XG6481 XI11_4/XI3/net5 XI11_4/preck DECAP_INV_G8
XG6482 sck_bar XI11_4/XI3/net018 DECAP_INV_G9
XG6483 XI11_4/XI3/net018 XI11_4/XI3/net012 DECAP_INV_G9
XG6484 XI11_4/XI3/net014 XI11_4/XI3/net7 DECAP_INV_G9
XG6485 XI11_4/XI3/net012 XI11_4/XI3/net014 DECAP_INV_G9
XG6486 XI11_4/XI4/net063 XI11_4/XI4/net0112 DECAP_INV_G10
XG6487 XI11_4/XI4/net26 XI11_4/XI4/net089 DECAP_INV_G10
XG6488 XI11_4/XI4/data_out XI11_4/XI4/data_out_ DECAP_INV_G10
XG6489 XI11_4/XI4/net20 XI11_4/XI4/net0103 DECAP_INV_G10
XG6490 XI11_4/net12 XI11_4/XI4/net32 DECAP_INV_G7
XG6491 XI11_4/net9 XI11_4/XI4/net52 DECAP_INV_G7
XG6492 XI11_4/XI4/data_out_ XI11_4/XI4/data_out DECAP_INV_G10
XG6493 XI11_4/XI0/XI0_63/d__15_ XI11_4/XI0/XI0_63/d_15_ DECAP_INV_G11
XG6494 XI11_4/XI0/XI0_63/d__14_ XI11_4/XI0/XI0_63/d_14_ DECAP_INV_G11
XG6495 XI11_4/XI0/XI0_63/d__13_ XI11_4/XI0/XI0_63/d_13_ DECAP_INV_G11
XG6496 XI11_4/XI0/XI0_63/d__12_ XI11_4/XI0/XI0_63/d_12_ DECAP_INV_G11
XG6497 XI11_4/XI0/XI0_63/d__11_ XI11_4/XI0/XI0_63/d_11_ DECAP_INV_G11
XG6498 XI11_4/XI0/XI0_63/d__10_ XI11_4/XI0/XI0_63/d_10_ DECAP_INV_G11
XG6499 XI11_4/XI0/XI0_63/d__9_ XI11_4/XI0/XI0_63/d_9_ DECAP_INV_G11
XG6500 XI11_4/XI0/XI0_63/d__8_ XI11_4/XI0/XI0_63/d_8_ DECAP_INV_G11
XG6501 XI11_4/XI0/XI0_63/d__7_ XI11_4/XI0/XI0_63/d_7_ DECAP_INV_G11
XG6502 XI11_4/XI0/XI0_63/d__6_ XI11_4/XI0/XI0_63/d_6_ DECAP_INV_G11
XG6503 XI11_4/XI0/XI0_63/d__5_ XI11_4/XI0/XI0_63/d_5_ DECAP_INV_G11
XG6504 XI11_4/XI0/XI0_63/d__4_ XI11_4/XI0/XI0_63/d_4_ DECAP_INV_G11
XG6505 XI11_4/XI0/XI0_63/d__3_ XI11_4/XI0/XI0_63/d_3_ DECAP_INV_G11
XG6506 XI11_4/XI0/XI0_63/d__2_ XI11_4/XI0/XI0_63/d_2_ DECAP_INV_G11
XG6507 XI11_4/XI0/XI0_63/d__1_ XI11_4/XI0/XI0_63/d_1_ DECAP_INV_G11
XG6508 XI11_4/XI0/XI0_63/d__0_ XI11_4/XI0/XI0_63/d_0_ DECAP_INV_G11
XG6509 XI11_4/XI0/XI0_63/d_15_ XI11_4/XI0/XI0_63/d__15_ DECAP_INV_G11
XG6510 XI11_4/XI0/XI0_63/d_14_ XI11_4/XI0/XI0_63/d__14_ DECAP_INV_G11
XG6511 XI11_4/XI0/XI0_63/d_13_ XI11_4/XI0/XI0_63/d__13_ DECAP_INV_G11
XG6512 XI11_4/XI0/XI0_63/d_12_ XI11_4/XI0/XI0_63/d__12_ DECAP_INV_G11
XG6513 XI11_4/XI0/XI0_63/d_11_ XI11_4/XI0/XI0_63/d__11_ DECAP_INV_G11
XG6514 XI11_4/XI0/XI0_63/d_10_ XI11_4/XI0/XI0_63/d__10_ DECAP_INV_G11
XG6515 XI11_4/XI0/XI0_63/d_9_ XI11_4/XI0/XI0_63/d__9_ DECAP_INV_G11
XG6516 XI11_4/XI0/XI0_63/d_8_ XI11_4/XI0/XI0_63/d__8_ DECAP_INV_G11
XG6517 XI11_4/XI0/XI0_63/d_7_ XI11_4/XI0/XI0_63/d__7_ DECAP_INV_G11
XG6518 XI11_4/XI0/XI0_63/d_6_ XI11_4/XI0/XI0_63/d__6_ DECAP_INV_G11
XG6519 XI11_4/XI0/XI0_63/d_5_ XI11_4/XI0/XI0_63/d__5_ DECAP_INV_G11
XG6520 XI11_4/XI0/XI0_63/d_4_ XI11_4/XI0/XI0_63/d__4_ DECAP_INV_G11
XG6521 XI11_4/XI0/XI0_63/d_3_ XI11_4/XI0/XI0_63/d__3_ DECAP_INV_G11
XG6522 XI11_4/XI0/XI0_63/d_2_ XI11_4/XI0/XI0_63/d__2_ DECAP_INV_G11
XG6523 XI11_4/XI0/XI0_63/d_1_ XI11_4/XI0/XI0_63/d__1_ DECAP_INV_G11
XG6524 XI11_4/XI0/XI0_63/d_0_ XI11_4/XI0/XI0_63/d__0_ DECAP_INV_G11
XG6525 XI11_4/XI0/XI0_62/d__15_ XI11_4/XI0/XI0_62/d_15_ DECAP_INV_G11
XG6526 XI11_4/XI0/XI0_62/d__14_ XI11_4/XI0/XI0_62/d_14_ DECAP_INV_G11
XG6527 XI11_4/XI0/XI0_62/d__13_ XI11_4/XI0/XI0_62/d_13_ DECAP_INV_G11
XG6528 XI11_4/XI0/XI0_62/d__12_ XI11_4/XI0/XI0_62/d_12_ DECAP_INV_G11
XG6529 XI11_4/XI0/XI0_62/d__11_ XI11_4/XI0/XI0_62/d_11_ DECAP_INV_G11
XG6530 XI11_4/XI0/XI0_62/d__10_ XI11_4/XI0/XI0_62/d_10_ DECAP_INV_G11
XG6531 XI11_4/XI0/XI0_62/d__9_ XI11_4/XI0/XI0_62/d_9_ DECAP_INV_G11
XG6532 XI11_4/XI0/XI0_62/d__8_ XI11_4/XI0/XI0_62/d_8_ DECAP_INV_G11
XG6533 XI11_4/XI0/XI0_62/d__7_ XI11_4/XI0/XI0_62/d_7_ DECAP_INV_G11
XG6534 XI11_4/XI0/XI0_62/d__6_ XI11_4/XI0/XI0_62/d_6_ DECAP_INV_G11
XG6535 XI11_4/XI0/XI0_62/d__5_ XI11_4/XI0/XI0_62/d_5_ DECAP_INV_G11
XG6536 XI11_4/XI0/XI0_62/d__4_ XI11_4/XI0/XI0_62/d_4_ DECAP_INV_G11
XG6537 XI11_4/XI0/XI0_62/d__3_ XI11_4/XI0/XI0_62/d_3_ DECAP_INV_G11
XG6538 XI11_4/XI0/XI0_62/d__2_ XI11_4/XI0/XI0_62/d_2_ DECAP_INV_G11
XG6539 XI11_4/XI0/XI0_62/d__1_ XI11_4/XI0/XI0_62/d_1_ DECAP_INV_G11
XG6540 XI11_4/XI0/XI0_62/d__0_ XI11_4/XI0/XI0_62/d_0_ DECAP_INV_G11
XG6541 XI11_4/XI0/XI0_62/d_15_ XI11_4/XI0/XI0_62/d__15_ DECAP_INV_G11
XG6542 XI11_4/XI0/XI0_62/d_14_ XI11_4/XI0/XI0_62/d__14_ DECAP_INV_G11
XG6543 XI11_4/XI0/XI0_62/d_13_ XI11_4/XI0/XI0_62/d__13_ DECAP_INV_G11
XG6544 XI11_4/XI0/XI0_62/d_12_ XI11_4/XI0/XI0_62/d__12_ DECAP_INV_G11
XG6545 XI11_4/XI0/XI0_62/d_11_ XI11_4/XI0/XI0_62/d__11_ DECAP_INV_G11
XG6546 XI11_4/XI0/XI0_62/d_10_ XI11_4/XI0/XI0_62/d__10_ DECAP_INV_G11
XG6547 XI11_4/XI0/XI0_62/d_9_ XI11_4/XI0/XI0_62/d__9_ DECAP_INV_G11
XG6548 XI11_4/XI0/XI0_62/d_8_ XI11_4/XI0/XI0_62/d__8_ DECAP_INV_G11
XG6549 XI11_4/XI0/XI0_62/d_7_ XI11_4/XI0/XI0_62/d__7_ DECAP_INV_G11
XG6550 XI11_4/XI0/XI0_62/d_6_ XI11_4/XI0/XI0_62/d__6_ DECAP_INV_G11
XG6551 XI11_4/XI0/XI0_62/d_5_ XI11_4/XI0/XI0_62/d__5_ DECAP_INV_G11
XG6552 XI11_4/XI0/XI0_62/d_4_ XI11_4/XI0/XI0_62/d__4_ DECAP_INV_G11
XG6553 XI11_4/XI0/XI0_62/d_3_ XI11_4/XI0/XI0_62/d__3_ DECAP_INV_G11
XG6554 XI11_4/XI0/XI0_62/d_2_ XI11_4/XI0/XI0_62/d__2_ DECAP_INV_G11
XG6555 XI11_4/XI0/XI0_62/d_1_ XI11_4/XI0/XI0_62/d__1_ DECAP_INV_G11
XG6556 XI11_4/XI0/XI0_62/d_0_ XI11_4/XI0/XI0_62/d__0_ DECAP_INV_G11
XG6557 XI11_4/XI0/XI0_61/d__15_ XI11_4/XI0/XI0_61/d_15_ DECAP_INV_G11
XG6558 XI11_4/XI0/XI0_61/d__14_ XI11_4/XI0/XI0_61/d_14_ DECAP_INV_G11
XG6559 XI11_4/XI0/XI0_61/d__13_ XI11_4/XI0/XI0_61/d_13_ DECAP_INV_G11
XG6560 XI11_4/XI0/XI0_61/d__12_ XI11_4/XI0/XI0_61/d_12_ DECAP_INV_G11
XG6561 XI11_4/XI0/XI0_61/d__11_ XI11_4/XI0/XI0_61/d_11_ DECAP_INV_G11
XG6562 XI11_4/XI0/XI0_61/d__10_ XI11_4/XI0/XI0_61/d_10_ DECAP_INV_G11
XG6563 XI11_4/XI0/XI0_61/d__9_ XI11_4/XI0/XI0_61/d_9_ DECAP_INV_G11
XG6564 XI11_4/XI0/XI0_61/d__8_ XI11_4/XI0/XI0_61/d_8_ DECAP_INV_G11
XG6565 XI11_4/XI0/XI0_61/d__7_ XI11_4/XI0/XI0_61/d_7_ DECAP_INV_G11
XG6566 XI11_4/XI0/XI0_61/d__6_ XI11_4/XI0/XI0_61/d_6_ DECAP_INV_G11
XG6567 XI11_4/XI0/XI0_61/d__5_ XI11_4/XI0/XI0_61/d_5_ DECAP_INV_G11
XG6568 XI11_4/XI0/XI0_61/d__4_ XI11_4/XI0/XI0_61/d_4_ DECAP_INV_G11
XG6569 XI11_4/XI0/XI0_61/d__3_ XI11_4/XI0/XI0_61/d_3_ DECAP_INV_G11
XG6570 XI11_4/XI0/XI0_61/d__2_ XI11_4/XI0/XI0_61/d_2_ DECAP_INV_G11
XG6571 XI11_4/XI0/XI0_61/d__1_ XI11_4/XI0/XI0_61/d_1_ DECAP_INV_G11
XG6572 XI11_4/XI0/XI0_61/d__0_ XI11_4/XI0/XI0_61/d_0_ DECAP_INV_G11
XG6573 XI11_4/XI0/XI0_61/d_15_ XI11_4/XI0/XI0_61/d__15_ DECAP_INV_G11
XG6574 XI11_4/XI0/XI0_61/d_14_ XI11_4/XI0/XI0_61/d__14_ DECAP_INV_G11
XG6575 XI11_4/XI0/XI0_61/d_13_ XI11_4/XI0/XI0_61/d__13_ DECAP_INV_G11
XG6576 XI11_4/XI0/XI0_61/d_12_ XI11_4/XI0/XI0_61/d__12_ DECAP_INV_G11
XG6577 XI11_4/XI0/XI0_61/d_11_ XI11_4/XI0/XI0_61/d__11_ DECAP_INV_G11
XG6578 XI11_4/XI0/XI0_61/d_10_ XI11_4/XI0/XI0_61/d__10_ DECAP_INV_G11
XG6579 XI11_4/XI0/XI0_61/d_9_ XI11_4/XI0/XI0_61/d__9_ DECAP_INV_G11
XG6580 XI11_4/XI0/XI0_61/d_8_ XI11_4/XI0/XI0_61/d__8_ DECAP_INV_G11
XG6581 XI11_4/XI0/XI0_61/d_7_ XI11_4/XI0/XI0_61/d__7_ DECAP_INV_G11
XG6582 XI11_4/XI0/XI0_61/d_6_ XI11_4/XI0/XI0_61/d__6_ DECAP_INV_G11
XG6583 XI11_4/XI0/XI0_61/d_5_ XI11_4/XI0/XI0_61/d__5_ DECAP_INV_G11
XG6584 XI11_4/XI0/XI0_61/d_4_ XI11_4/XI0/XI0_61/d__4_ DECAP_INV_G11
XG6585 XI11_4/XI0/XI0_61/d_3_ XI11_4/XI0/XI0_61/d__3_ DECAP_INV_G11
XG6586 XI11_4/XI0/XI0_61/d_2_ XI11_4/XI0/XI0_61/d__2_ DECAP_INV_G11
XG6587 XI11_4/XI0/XI0_61/d_1_ XI11_4/XI0/XI0_61/d__1_ DECAP_INV_G11
XG6588 XI11_4/XI0/XI0_61/d_0_ XI11_4/XI0/XI0_61/d__0_ DECAP_INV_G11
XG6589 XI11_4/XI0/XI0_60/d__15_ XI11_4/XI0/XI0_60/d_15_ DECAP_INV_G11
XG6590 XI11_4/XI0/XI0_60/d__14_ XI11_4/XI0/XI0_60/d_14_ DECAP_INV_G11
XG6591 XI11_4/XI0/XI0_60/d__13_ XI11_4/XI0/XI0_60/d_13_ DECAP_INV_G11
XG6592 XI11_4/XI0/XI0_60/d__12_ XI11_4/XI0/XI0_60/d_12_ DECAP_INV_G11
XG6593 XI11_4/XI0/XI0_60/d__11_ XI11_4/XI0/XI0_60/d_11_ DECAP_INV_G11
XG6594 XI11_4/XI0/XI0_60/d__10_ XI11_4/XI0/XI0_60/d_10_ DECAP_INV_G11
XG6595 XI11_4/XI0/XI0_60/d__9_ XI11_4/XI0/XI0_60/d_9_ DECAP_INV_G11
XG6596 XI11_4/XI0/XI0_60/d__8_ XI11_4/XI0/XI0_60/d_8_ DECAP_INV_G11
XG6597 XI11_4/XI0/XI0_60/d__7_ XI11_4/XI0/XI0_60/d_7_ DECAP_INV_G11
XG6598 XI11_4/XI0/XI0_60/d__6_ XI11_4/XI0/XI0_60/d_6_ DECAP_INV_G11
XG6599 XI11_4/XI0/XI0_60/d__5_ XI11_4/XI0/XI0_60/d_5_ DECAP_INV_G11
XG6600 XI11_4/XI0/XI0_60/d__4_ XI11_4/XI0/XI0_60/d_4_ DECAP_INV_G11
XG6601 XI11_4/XI0/XI0_60/d__3_ XI11_4/XI0/XI0_60/d_3_ DECAP_INV_G11
XG6602 XI11_4/XI0/XI0_60/d__2_ XI11_4/XI0/XI0_60/d_2_ DECAP_INV_G11
XG6603 XI11_4/XI0/XI0_60/d__1_ XI11_4/XI0/XI0_60/d_1_ DECAP_INV_G11
XG6604 XI11_4/XI0/XI0_60/d__0_ XI11_4/XI0/XI0_60/d_0_ DECAP_INV_G11
XG6605 XI11_4/XI0/XI0_60/d_15_ XI11_4/XI0/XI0_60/d__15_ DECAP_INV_G11
XG6606 XI11_4/XI0/XI0_60/d_14_ XI11_4/XI0/XI0_60/d__14_ DECAP_INV_G11
XG6607 XI11_4/XI0/XI0_60/d_13_ XI11_4/XI0/XI0_60/d__13_ DECAP_INV_G11
XG6608 XI11_4/XI0/XI0_60/d_12_ XI11_4/XI0/XI0_60/d__12_ DECAP_INV_G11
XG6609 XI11_4/XI0/XI0_60/d_11_ XI11_4/XI0/XI0_60/d__11_ DECAP_INV_G11
XG6610 XI11_4/XI0/XI0_60/d_10_ XI11_4/XI0/XI0_60/d__10_ DECAP_INV_G11
XG6611 XI11_4/XI0/XI0_60/d_9_ XI11_4/XI0/XI0_60/d__9_ DECAP_INV_G11
XG6612 XI11_4/XI0/XI0_60/d_8_ XI11_4/XI0/XI0_60/d__8_ DECAP_INV_G11
XG6613 XI11_4/XI0/XI0_60/d_7_ XI11_4/XI0/XI0_60/d__7_ DECAP_INV_G11
XG6614 XI11_4/XI0/XI0_60/d_6_ XI11_4/XI0/XI0_60/d__6_ DECAP_INV_G11
XG6615 XI11_4/XI0/XI0_60/d_5_ XI11_4/XI0/XI0_60/d__5_ DECAP_INV_G11
XG6616 XI11_4/XI0/XI0_60/d_4_ XI11_4/XI0/XI0_60/d__4_ DECAP_INV_G11
XG6617 XI11_4/XI0/XI0_60/d_3_ XI11_4/XI0/XI0_60/d__3_ DECAP_INV_G11
XG6618 XI11_4/XI0/XI0_60/d_2_ XI11_4/XI0/XI0_60/d__2_ DECAP_INV_G11
XG6619 XI11_4/XI0/XI0_60/d_1_ XI11_4/XI0/XI0_60/d__1_ DECAP_INV_G11
XG6620 XI11_4/XI0/XI0_60/d_0_ XI11_4/XI0/XI0_60/d__0_ DECAP_INV_G11
XG6621 XI11_4/XI0/XI0_59/d__15_ XI11_4/XI0/XI0_59/d_15_ DECAP_INV_G11
XG6622 XI11_4/XI0/XI0_59/d__14_ XI11_4/XI0/XI0_59/d_14_ DECAP_INV_G11
XG6623 XI11_4/XI0/XI0_59/d__13_ XI11_4/XI0/XI0_59/d_13_ DECAP_INV_G11
XG6624 XI11_4/XI0/XI0_59/d__12_ XI11_4/XI0/XI0_59/d_12_ DECAP_INV_G11
XG6625 XI11_4/XI0/XI0_59/d__11_ XI11_4/XI0/XI0_59/d_11_ DECAP_INV_G11
XG6626 XI11_4/XI0/XI0_59/d__10_ XI11_4/XI0/XI0_59/d_10_ DECAP_INV_G11
XG6627 XI11_4/XI0/XI0_59/d__9_ XI11_4/XI0/XI0_59/d_9_ DECAP_INV_G11
XG6628 XI11_4/XI0/XI0_59/d__8_ XI11_4/XI0/XI0_59/d_8_ DECAP_INV_G11
XG6629 XI11_4/XI0/XI0_59/d__7_ XI11_4/XI0/XI0_59/d_7_ DECAP_INV_G11
XG6630 XI11_4/XI0/XI0_59/d__6_ XI11_4/XI0/XI0_59/d_6_ DECAP_INV_G11
XG6631 XI11_4/XI0/XI0_59/d__5_ XI11_4/XI0/XI0_59/d_5_ DECAP_INV_G11
XG6632 XI11_4/XI0/XI0_59/d__4_ XI11_4/XI0/XI0_59/d_4_ DECAP_INV_G11
XG6633 XI11_4/XI0/XI0_59/d__3_ XI11_4/XI0/XI0_59/d_3_ DECAP_INV_G11
XG6634 XI11_4/XI0/XI0_59/d__2_ XI11_4/XI0/XI0_59/d_2_ DECAP_INV_G11
XG6635 XI11_4/XI0/XI0_59/d__1_ XI11_4/XI0/XI0_59/d_1_ DECAP_INV_G11
XG6636 XI11_4/XI0/XI0_59/d__0_ XI11_4/XI0/XI0_59/d_0_ DECAP_INV_G11
XG6637 XI11_4/XI0/XI0_59/d_15_ XI11_4/XI0/XI0_59/d__15_ DECAP_INV_G11
XG6638 XI11_4/XI0/XI0_59/d_14_ XI11_4/XI0/XI0_59/d__14_ DECAP_INV_G11
XG6639 XI11_4/XI0/XI0_59/d_13_ XI11_4/XI0/XI0_59/d__13_ DECAP_INV_G11
XG6640 XI11_4/XI0/XI0_59/d_12_ XI11_4/XI0/XI0_59/d__12_ DECAP_INV_G11
XG6641 XI11_4/XI0/XI0_59/d_11_ XI11_4/XI0/XI0_59/d__11_ DECAP_INV_G11
XG6642 XI11_4/XI0/XI0_59/d_10_ XI11_4/XI0/XI0_59/d__10_ DECAP_INV_G11
XG6643 XI11_4/XI0/XI0_59/d_9_ XI11_4/XI0/XI0_59/d__9_ DECAP_INV_G11
XG6644 XI11_4/XI0/XI0_59/d_8_ XI11_4/XI0/XI0_59/d__8_ DECAP_INV_G11
XG6645 XI11_4/XI0/XI0_59/d_7_ XI11_4/XI0/XI0_59/d__7_ DECAP_INV_G11
XG6646 XI11_4/XI0/XI0_59/d_6_ XI11_4/XI0/XI0_59/d__6_ DECAP_INV_G11
XG6647 XI11_4/XI0/XI0_59/d_5_ XI11_4/XI0/XI0_59/d__5_ DECAP_INV_G11
XG6648 XI11_4/XI0/XI0_59/d_4_ XI11_4/XI0/XI0_59/d__4_ DECAP_INV_G11
XG6649 XI11_4/XI0/XI0_59/d_3_ XI11_4/XI0/XI0_59/d__3_ DECAP_INV_G11
XG6650 XI11_4/XI0/XI0_59/d_2_ XI11_4/XI0/XI0_59/d__2_ DECAP_INV_G11
XG6651 XI11_4/XI0/XI0_59/d_1_ XI11_4/XI0/XI0_59/d__1_ DECAP_INV_G11
XG6652 XI11_4/XI0/XI0_59/d_0_ XI11_4/XI0/XI0_59/d__0_ DECAP_INV_G11
XG6653 XI11_4/XI0/XI0_58/d__15_ XI11_4/XI0/XI0_58/d_15_ DECAP_INV_G11
XG6654 XI11_4/XI0/XI0_58/d__14_ XI11_4/XI0/XI0_58/d_14_ DECAP_INV_G11
XG6655 XI11_4/XI0/XI0_58/d__13_ XI11_4/XI0/XI0_58/d_13_ DECAP_INV_G11
XG6656 XI11_4/XI0/XI0_58/d__12_ XI11_4/XI0/XI0_58/d_12_ DECAP_INV_G11
XG6657 XI11_4/XI0/XI0_58/d__11_ XI11_4/XI0/XI0_58/d_11_ DECAP_INV_G11
XG6658 XI11_4/XI0/XI0_58/d__10_ XI11_4/XI0/XI0_58/d_10_ DECAP_INV_G11
XG6659 XI11_4/XI0/XI0_58/d__9_ XI11_4/XI0/XI0_58/d_9_ DECAP_INV_G11
XG6660 XI11_4/XI0/XI0_58/d__8_ XI11_4/XI0/XI0_58/d_8_ DECAP_INV_G11
XG6661 XI11_4/XI0/XI0_58/d__7_ XI11_4/XI0/XI0_58/d_7_ DECAP_INV_G11
XG6662 XI11_4/XI0/XI0_58/d__6_ XI11_4/XI0/XI0_58/d_6_ DECAP_INV_G11
XG6663 XI11_4/XI0/XI0_58/d__5_ XI11_4/XI0/XI0_58/d_5_ DECAP_INV_G11
XG6664 XI11_4/XI0/XI0_58/d__4_ XI11_4/XI0/XI0_58/d_4_ DECAP_INV_G11
XG6665 XI11_4/XI0/XI0_58/d__3_ XI11_4/XI0/XI0_58/d_3_ DECAP_INV_G11
XG6666 XI11_4/XI0/XI0_58/d__2_ XI11_4/XI0/XI0_58/d_2_ DECAP_INV_G11
XG6667 XI11_4/XI0/XI0_58/d__1_ XI11_4/XI0/XI0_58/d_1_ DECAP_INV_G11
XG6668 XI11_4/XI0/XI0_58/d__0_ XI11_4/XI0/XI0_58/d_0_ DECAP_INV_G11
XG6669 XI11_4/XI0/XI0_58/d_15_ XI11_4/XI0/XI0_58/d__15_ DECAP_INV_G11
XG6670 XI11_4/XI0/XI0_58/d_14_ XI11_4/XI0/XI0_58/d__14_ DECAP_INV_G11
XG6671 XI11_4/XI0/XI0_58/d_13_ XI11_4/XI0/XI0_58/d__13_ DECAP_INV_G11
XG6672 XI11_4/XI0/XI0_58/d_12_ XI11_4/XI0/XI0_58/d__12_ DECAP_INV_G11
XG6673 XI11_4/XI0/XI0_58/d_11_ XI11_4/XI0/XI0_58/d__11_ DECAP_INV_G11
XG6674 XI11_4/XI0/XI0_58/d_10_ XI11_4/XI0/XI0_58/d__10_ DECAP_INV_G11
XG6675 XI11_4/XI0/XI0_58/d_9_ XI11_4/XI0/XI0_58/d__9_ DECAP_INV_G11
XG6676 XI11_4/XI0/XI0_58/d_8_ XI11_4/XI0/XI0_58/d__8_ DECAP_INV_G11
XG6677 XI11_4/XI0/XI0_58/d_7_ XI11_4/XI0/XI0_58/d__7_ DECAP_INV_G11
XG6678 XI11_4/XI0/XI0_58/d_6_ XI11_4/XI0/XI0_58/d__6_ DECAP_INV_G11
XG6679 XI11_4/XI0/XI0_58/d_5_ XI11_4/XI0/XI0_58/d__5_ DECAP_INV_G11
XG6680 XI11_4/XI0/XI0_58/d_4_ XI11_4/XI0/XI0_58/d__4_ DECAP_INV_G11
XG6681 XI11_4/XI0/XI0_58/d_3_ XI11_4/XI0/XI0_58/d__3_ DECAP_INV_G11
XG6682 XI11_4/XI0/XI0_58/d_2_ XI11_4/XI0/XI0_58/d__2_ DECAP_INV_G11
XG6683 XI11_4/XI0/XI0_58/d_1_ XI11_4/XI0/XI0_58/d__1_ DECAP_INV_G11
XG6684 XI11_4/XI0/XI0_58/d_0_ XI11_4/XI0/XI0_58/d__0_ DECAP_INV_G11
XG6685 XI11_4/XI0/XI0_57/d__15_ XI11_4/XI0/XI0_57/d_15_ DECAP_INV_G11
XG6686 XI11_4/XI0/XI0_57/d__14_ XI11_4/XI0/XI0_57/d_14_ DECAP_INV_G11
XG6687 XI11_4/XI0/XI0_57/d__13_ XI11_4/XI0/XI0_57/d_13_ DECAP_INV_G11
XG6688 XI11_4/XI0/XI0_57/d__12_ XI11_4/XI0/XI0_57/d_12_ DECAP_INV_G11
XG6689 XI11_4/XI0/XI0_57/d__11_ XI11_4/XI0/XI0_57/d_11_ DECAP_INV_G11
XG6690 XI11_4/XI0/XI0_57/d__10_ XI11_4/XI0/XI0_57/d_10_ DECAP_INV_G11
XG6691 XI11_4/XI0/XI0_57/d__9_ XI11_4/XI0/XI0_57/d_9_ DECAP_INV_G11
XG6692 XI11_4/XI0/XI0_57/d__8_ XI11_4/XI0/XI0_57/d_8_ DECAP_INV_G11
XG6693 XI11_4/XI0/XI0_57/d__7_ XI11_4/XI0/XI0_57/d_7_ DECAP_INV_G11
XG6694 XI11_4/XI0/XI0_57/d__6_ XI11_4/XI0/XI0_57/d_6_ DECAP_INV_G11
XG6695 XI11_4/XI0/XI0_57/d__5_ XI11_4/XI0/XI0_57/d_5_ DECAP_INV_G11
XG6696 XI11_4/XI0/XI0_57/d__4_ XI11_4/XI0/XI0_57/d_4_ DECAP_INV_G11
XG6697 XI11_4/XI0/XI0_57/d__3_ XI11_4/XI0/XI0_57/d_3_ DECAP_INV_G11
XG6698 XI11_4/XI0/XI0_57/d__2_ XI11_4/XI0/XI0_57/d_2_ DECAP_INV_G11
XG6699 XI11_4/XI0/XI0_57/d__1_ XI11_4/XI0/XI0_57/d_1_ DECAP_INV_G11
XG6700 XI11_4/XI0/XI0_57/d__0_ XI11_4/XI0/XI0_57/d_0_ DECAP_INV_G11
XG6701 XI11_4/XI0/XI0_57/d_15_ XI11_4/XI0/XI0_57/d__15_ DECAP_INV_G11
XG6702 XI11_4/XI0/XI0_57/d_14_ XI11_4/XI0/XI0_57/d__14_ DECAP_INV_G11
XG6703 XI11_4/XI0/XI0_57/d_13_ XI11_4/XI0/XI0_57/d__13_ DECAP_INV_G11
XG6704 XI11_4/XI0/XI0_57/d_12_ XI11_4/XI0/XI0_57/d__12_ DECAP_INV_G11
XG6705 XI11_4/XI0/XI0_57/d_11_ XI11_4/XI0/XI0_57/d__11_ DECAP_INV_G11
XG6706 XI11_4/XI0/XI0_57/d_10_ XI11_4/XI0/XI0_57/d__10_ DECAP_INV_G11
XG6707 XI11_4/XI0/XI0_57/d_9_ XI11_4/XI0/XI0_57/d__9_ DECAP_INV_G11
XG6708 XI11_4/XI0/XI0_57/d_8_ XI11_4/XI0/XI0_57/d__8_ DECAP_INV_G11
XG6709 XI11_4/XI0/XI0_57/d_7_ XI11_4/XI0/XI0_57/d__7_ DECAP_INV_G11
XG6710 XI11_4/XI0/XI0_57/d_6_ XI11_4/XI0/XI0_57/d__6_ DECAP_INV_G11
XG6711 XI11_4/XI0/XI0_57/d_5_ XI11_4/XI0/XI0_57/d__5_ DECAP_INV_G11
XG6712 XI11_4/XI0/XI0_57/d_4_ XI11_4/XI0/XI0_57/d__4_ DECAP_INV_G11
XG6713 XI11_4/XI0/XI0_57/d_3_ XI11_4/XI0/XI0_57/d__3_ DECAP_INV_G11
XG6714 XI11_4/XI0/XI0_57/d_2_ XI11_4/XI0/XI0_57/d__2_ DECAP_INV_G11
XG6715 XI11_4/XI0/XI0_57/d_1_ XI11_4/XI0/XI0_57/d__1_ DECAP_INV_G11
XG6716 XI11_4/XI0/XI0_57/d_0_ XI11_4/XI0/XI0_57/d__0_ DECAP_INV_G11
XG6717 XI11_4/XI0/XI0_56/d__15_ XI11_4/XI0/XI0_56/d_15_ DECAP_INV_G11
XG6718 XI11_4/XI0/XI0_56/d__14_ XI11_4/XI0/XI0_56/d_14_ DECAP_INV_G11
XG6719 XI11_4/XI0/XI0_56/d__13_ XI11_4/XI0/XI0_56/d_13_ DECAP_INV_G11
XG6720 XI11_4/XI0/XI0_56/d__12_ XI11_4/XI0/XI0_56/d_12_ DECAP_INV_G11
XG6721 XI11_4/XI0/XI0_56/d__11_ XI11_4/XI0/XI0_56/d_11_ DECAP_INV_G11
XG6722 XI11_4/XI0/XI0_56/d__10_ XI11_4/XI0/XI0_56/d_10_ DECAP_INV_G11
XG6723 XI11_4/XI0/XI0_56/d__9_ XI11_4/XI0/XI0_56/d_9_ DECAP_INV_G11
XG6724 XI11_4/XI0/XI0_56/d__8_ XI11_4/XI0/XI0_56/d_8_ DECAP_INV_G11
XG6725 XI11_4/XI0/XI0_56/d__7_ XI11_4/XI0/XI0_56/d_7_ DECAP_INV_G11
XG6726 XI11_4/XI0/XI0_56/d__6_ XI11_4/XI0/XI0_56/d_6_ DECAP_INV_G11
XG6727 XI11_4/XI0/XI0_56/d__5_ XI11_4/XI0/XI0_56/d_5_ DECAP_INV_G11
XG6728 XI11_4/XI0/XI0_56/d__4_ XI11_4/XI0/XI0_56/d_4_ DECAP_INV_G11
XG6729 XI11_4/XI0/XI0_56/d__3_ XI11_4/XI0/XI0_56/d_3_ DECAP_INV_G11
XG6730 XI11_4/XI0/XI0_56/d__2_ XI11_4/XI0/XI0_56/d_2_ DECAP_INV_G11
XG6731 XI11_4/XI0/XI0_56/d__1_ XI11_4/XI0/XI0_56/d_1_ DECAP_INV_G11
XG6732 XI11_4/XI0/XI0_56/d__0_ XI11_4/XI0/XI0_56/d_0_ DECAP_INV_G11
XG6733 XI11_4/XI0/XI0_56/d_15_ XI11_4/XI0/XI0_56/d__15_ DECAP_INV_G11
XG6734 XI11_4/XI0/XI0_56/d_14_ XI11_4/XI0/XI0_56/d__14_ DECAP_INV_G11
XG6735 XI11_4/XI0/XI0_56/d_13_ XI11_4/XI0/XI0_56/d__13_ DECAP_INV_G11
XG6736 XI11_4/XI0/XI0_56/d_12_ XI11_4/XI0/XI0_56/d__12_ DECAP_INV_G11
XG6737 XI11_4/XI0/XI0_56/d_11_ XI11_4/XI0/XI0_56/d__11_ DECAP_INV_G11
XG6738 XI11_4/XI0/XI0_56/d_10_ XI11_4/XI0/XI0_56/d__10_ DECAP_INV_G11
XG6739 XI11_4/XI0/XI0_56/d_9_ XI11_4/XI0/XI0_56/d__9_ DECAP_INV_G11
XG6740 XI11_4/XI0/XI0_56/d_8_ XI11_4/XI0/XI0_56/d__8_ DECAP_INV_G11
XG6741 XI11_4/XI0/XI0_56/d_7_ XI11_4/XI0/XI0_56/d__7_ DECAP_INV_G11
XG6742 XI11_4/XI0/XI0_56/d_6_ XI11_4/XI0/XI0_56/d__6_ DECAP_INV_G11
XG6743 XI11_4/XI0/XI0_56/d_5_ XI11_4/XI0/XI0_56/d__5_ DECAP_INV_G11
XG6744 XI11_4/XI0/XI0_56/d_4_ XI11_4/XI0/XI0_56/d__4_ DECAP_INV_G11
XG6745 XI11_4/XI0/XI0_56/d_3_ XI11_4/XI0/XI0_56/d__3_ DECAP_INV_G11
XG6746 XI11_4/XI0/XI0_56/d_2_ XI11_4/XI0/XI0_56/d__2_ DECAP_INV_G11
XG6747 XI11_4/XI0/XI0_56/d_1_ XI11_4/XI0/XI0_56/d__1_ DECAP_INV_G11
XG6748 XI11_4/XI0/XI0_56/d_0_ XI11_4/XI0/XI0_56/d__0_ DECAP_INV_G11
XG6749 XI11_4/XI0/XI0_55/d__15_ XI11_4/XI0/XI0_55/d_15_ DECAP_INV_G11
XG6750 XI11_4/XI0/XI0_55/d__14_ XI11_4/XI0/XI0_55/d_14_ DECAP_INV_G11
XG6751 XI11_4/XI0/XI0_55/d__13_ XI11_4/XI0/XI0_55/d_13_ DECAP_INV_G11
XG6752 XI11_4/XI0/XI0_55/d__12_ XI11_4/XI0/XI0_55/d_12_ DECAP_INV_G11
XG6753 XI11_4/XI0/XI0_55/d__11_ XI11_4/XI0/XI0_55/d_11_ DECAP_INV_G11
XG6754 XI11_4/XI0/XI0_55/d__10_ XI11_4/XI0/XI0_55/d_10_ DECAP_INV_G11
XG6755 XI11_4/XI0/XI0_55/d__9_ XI11_4/XI0/XI0_55/d_9_ DECAP_INV_G11
XG6756 XI11_4/XI0/XI0_55/d__8_ XI11_4/XI0/XI0_55/d_8_ DECAP_INV_G11
XG6757 XI11_4/XI0/XI0_55/d__7_ XI11_4/XI0/XI0_55/d_7_ DECAP_INV_G11
XG6758 XI11_4/XI0/XI0_55/d__6_ XI11_4/XI0/XI0_55/d_6_ DECAP_INV_G11
XG6759 XI11_4/XI0/XI0_55/d__5_ XI11_4/XI0/XI0_55/d_5_ DECAP_INV_G11
XG6760 XI11_4/XI0/XI0_55/d__4_ XI11_4/XI0/XI0_55/d_4_ DECAP_INV_G11
XG6761 XI11_4/XI0/XI0_55/d__3_ XI11_4/XI0/XI0_55/d_3_ DECAP_INV_G11
XG6762 XI11_4/XI0/XI0_55/d__2_ XI11_4/XI0/XI0_55/d_2_ DECAP_INV_G11
XG6763 XI11_4/XI0/XI0_55/d__1_ XI11_4/XI0/XI0_55/d_1_ DECAP_INV_G11
XG6764 XI11_4/XI0/XI0_55/d__0_ XI11_4/XI0/XI0_55/d_0_ DECAP_INV_G11
XG6765 XI11_4/XI0/XI0_55/d_15_ XI11_4/XI0/XI0_55/d__15_ DECAP_INV_G11
XG6766 XI11_4/XI0/XI0_55/d_14_ XI11_4/XI0/XI0_55/d__14_ DECAP_INV_G11
XG6767 XI11_4/XI0/XI0_55/d_13_ XI11_4/XI0/XI0_55/d__13_ DECAP_INV_G11
XG6768 XI11_4/XI0/XI0_55/d_12_ XI11_4/XI0/XI0_55/d__12_ DECAP_INV_G11
XG6769 XI11_4/XI0/XI0_55/d_11_ XI11_4/XI0/XI0_55/d__11_ DECAP_INV_G11
XG6770 XI11_4/XI0/XI0_55/d_10_ XI11_4/XI0/XI0_55/d__10_ DECAP_INV_G11
XG6771 XI11_4/XI0/XI0_55/d_9_ XI11_4/XI0/XI0_55/d__9_ DECAP_INV_G11
XG6772 XI11_4/XI0/XI0_55/d_8_ XI11_4/XI0/XI0_55/d__8_ DECAP_INV_G11
XG6773 XI11_4/XI0/XI0_55/d_7_ XI11_4/XI0/XI0_55/d__7_ DECAP_INV_G11
XG6774 XI11_4/XI0/XI0_55/d_6_ XI11_4/XI0/XI0_55/d__6_ DECAP_INV_G11
XG6775 XI11_4/XI0/XI0_55/d_5_ XI11_4/XI0/XI0_55/d__5_ DECAP_INV_G11
XG6776 XI11_4/XI0/XI0_55/d_4_ XI11_4/XI0/XI0_55/d__4_ DECAP_INV_G11
XG6777 XI11_4/XI0/XI0_55/d_3_ XI11_4/XI0/XI0_55/d__3_ DECAP_INV_G11
XG6778 XI11_4/XI0/XI0_55/d_2_ XI11_4/XI0/XI0_55/d__2_ DECAP_INV_G11
XG6779 XI11_4/XI0/XI0_55/d_1_ XI11_4/XI0/XI0_55/d__1_ DECAP_INV_G11
XG6780 XI11_4/XI0/XI0_55/d_0_ XI11_4/XI0/XI0_55/d__0_ DECAP_INV_G11
XG6781 XI11_4/XI0/XI0_54/d__15_ XI11_4/XI0/XI0_54/d_15_ DECAP_INV_G11
XG6782 XI11_4/XI0/XI0_54/d__14_ XI11_4/XI0/XI0_54/d_14_ DECAP_INV_G11
XG6783 XI11_4/XI0/XI0_54/d__13_ XI11_4/XI0/XI0_54/d_13_ DECAP_INV_G11
XG6784 XI11_4/XI0/XI0_54/d__12_ XI11_4/XI0/XI0_54/d_12_ DECAP_INV_G11
XG6785 XI11_4/XI0/XI0_54/d__11_ XI11_4/XI0/XI0_54/d_11_ DECAP_INV_G11
XG6786 XI11_4/XI0/XI0_54/d__10_ XI11_4/XI0/XI0_54/d_10_ DECAP_INV_G11
XG6787 XI11_4/XI0/XI0_54/d__9_ XI11_4/XI0/XI0_54/d_9_ DECAP_INV_G11
XG6788 XI11_4/XI0/XI0_54/d__8_ XI11_4/XI0/XI0_54/d_8_ DECAP_INV_G11
XG6789 XI11_4/XI0/XI0_54/d__7_ XI11_4/XI0/XI0_54/d_7_ DECAP_INV_G11
XG6790 XI11_4/XI0/XI0_54/d__6_ XI11_4/XI0/XI0_54/d_6_ DECAP_INV_G11
XG6791 XI11_4/XI0/XI0_54/d__5_ XI11_4/XI0/XI0_54/d_5_ DECAP_INV_G11
XG6792 XI11_4/XI0/XI0_54/d__4_ XI11_4/XI0/XI0_54/d_4_ DECAP_INV_G11
XG6793 XI11_4/XI0/XI0_54/d__3_ XI11_4/XI0/XI0_54/d_3_ DECAP_INV_G11
XG6794 XI11_4/XI0/XI0_54/d__2_ XI11_4/XI0/XI0_54/d_2_ DECAP_INV_G11
XG6795 XI11_4/XI0/XI0_54/d__1_ XI11_4/XI0/XI0_54/d_1_ DECAP_INV_G11
XG6796 XI11_4/XI0/XI0_54/d__0_ XI11_4/XI0/XI0_54/d_0_ DECAP_INV_G11
XG6797 XI11_4/XI0/XI0_54/d_15_ XI11_4/XI0/XI0_54/d__15_ DECAP_INV_G11
XG6798 XI11_4/XI0/XI0_54/d_14_ XI11_4/XI0/XI0_54/d__14_ DECAP_INV_G11
XG6799 XI11_4/XI0/XI0_54/d_13_ XI11_4/XI0/XI0_54/d__13_ DECAP_INV_G11
XG6800 XI11_4/XI0/XI0_54/d_12_ XI11_4/XI0/XI0_54/d__12_ DECAP_INV_G11
XG6801 XI11_4/XI0/XI0_54/d_11_ XI11_4/XI0/XI0_54/d__11_ DECAP_INV_G11
XG6802 XI11_4/XI0/XI0_54/d_10_ XI11_4/XI0/XI0_54/d__10_ DECAP_INV_G11
XG6803 XI11_4/XI0/XI0_54/d_9_ XI11_4/XI0/XI0_54/d__9_ DECAP_INV_G11
XG6804 XI11_4/XI0/XI0_54/d_8_ XI11_4/XI0/XI0_54/d__8_ DECAP_INV_G11
XG6805 XI11_4/XI0/XI0_54/d_7_ XI11_4/XI0/XI0_54/d__7_ DECAP_INV_G11
XG6806 XI11_4/XI0/XI0_54/d_6_ XI11_4/XI0/XI0_54/d__6_ DECAP_INV_G11
XG6807 XI11_4/XI0/XI0_54/d_5_ XI11_4/XI0/XI0_54/d__5_ DECAP_INV_G11
XG6808 XI11_4/XI0/XI0_54/d_4_ XI11_4/XI0/XI0_54/d__4_ DECAP_INV_G11
XG6809 XI11_4/XI0/XI0_54/d_3_ XI11_4/XI0/XI0_54/d__3_ DECAP_INV_G11
XG6810 XI11_4/XI0/XI0_54/d_2_ XI11_4/XI0/XI0_54/d__2_ DECAP_INV_G11
XG6811 XI11_4/XI0/XI0_54/d_1_ XI11_4/XI0/XI0_54/d__1_ DECAP_INV_G11
XG6812 XI11_4/XI0/XI0_54/d_0_ XI11_4/XI0/XI0_54/d__0_ DECAP_INV_G11
XG6813 XI11_4/XI0/XI0_53/d__15_ XI11_4/XI0/XI0_53/d_15_ DECAP_INV_G11
XG6814 XI11_4/XI0/XI0_53/d__14_ XI11_4/XI0/XI0_53/d_14_ DECAP_INV_G11
XG6815 XI11_4/XI0/XI0_53/d__13_ XI11_4/XI0/XI0_53/d_13_ DECAP_INV_G11
XG6816 XI11_4/XI0/XI0_53/d__12_ XI11_4/XI0/XI0_53/d_12_ DECAP_INV_G11
XG6817 XI11_4/XI0/XI0_53/d__11_ XI11_4/XI0/XI0_53/d_11_ DECAP_INV_G11
XG6818 XI11_4/XI0/XI0_53/d__10_ XI11_4/XI0/XI0_53/d_10_ DECAP_INV_G11
XG6819 XI11_4/XI0/XI0_53/d__9_ XI11_4/XI0/XI0_53/d_9_ DECAP_INV_G11
XG6820 XI11_4/XI0/XI0_53/d__8_ XI11_4/XI0/XI0_53/d_8_ DECAP_INV_G11
XG6821 XI11_4/XI0/XI0_53/d__7_ XI11_4/XI0/XI0_53/d_7_ DECAP_INV_G11
XG6822 XI11_4/XI0/XI0_53/d__6_ XI11_4/XI0/XI0_53/d_6_ DECAP_INV_G11
XG6823 XI11_4/XI0/XI0_53/d__5_ XI11_4/XI0/XI0_53/d_5_ DECAP_INV_G11
XG6824 XI11_4/XI0/XI0_53/d__4_ XI11_4/XI0/XI0_53/d_4_ DECAP_INV_G11
XG6825 XI11_4/XI0/XI0_53/d__3_ XI11_4/XI0/XI0_53/d_3_ DECAP_INV_G11
XG6826 XI11_4/XI0/XI0_53/d__2_ XI11_4/XI0/XI0_53/d_2_ DECAP_INV_G11
XG6827 XI11_4/XI0/XI0_53/d__1_ XI11_4/XI0/XI0_53/d_1_ DECAP_INV_G11
XG6828 XI11_4/XI0/XI0_53/d__0_ XI11_4/XI0/XI0_53/d_0_ DECAP_INV_G11
XG6829 XI11_4/XI0/XI0_53/d_15_ XI11_4/XI0/XI0_53/d__15_ DECAP_INV_G11
XG6830 XI11_4/XI0/XI0_53/d_14_ XI11_4/XI0/XI0_53/d__14_ DECAP_INV_G11
XG6831 XI11_4/XI0/XI0_53/d_13_ XI11_4/XI0/XI0_53/d__13_ DECAP_INV_G11
XG6832 XI11_4/XI0/XI0_53/d_12_ XI11_4/XI0/XI0_53/d__12_ DECAP_INV_G11
XG6833 XI11_4/XI0/XI0_53/d_11_ XI11_4/XI0/XI0_53/d__11_ DECAP_INV_G11
XG6834 XI11_4/XI0/XI0_53/d_10_ XI11_4/XI0/XI0_53/d__10_ DECAP_INV_G11
XG6835 XI11_4/XI0/XI0_53/d_9_ XI11_4/XI0/XI0_53/d__9_ DECAP_INV_G11
XG6836 XI11_4/XI0/XI0_53/d_8_ XI11_4/XI0/XI0_53/d__8_ DECAP_INV_G11
XG6837 XI11_4/XI0/XI0_53/d_7_ XI11_4/XI0/XI0_53/d__7_ DECAP_INV_G11
XG6838 XI11_4/XI0/XI0_53/d_6_ XI11_4/XI0/XI0_53/d__6_ DECAP_INV_G11
XG6839 XI11_4/XI0/XI0_53/d_5_ XI11_4/XI0/XI0_53/d__5_ DECAP_INV_G11
XG6840 XI11_4/XI0/XI0_53/d_4_ XI11_4/XI0/XI0_53/d__4_ DECAP_INV_G11
XG6841 XI11_4/XI0/XI0_53/d_3_ XI11_4/XI0/XI0_53/d__3_ DECAP_INV_G11
XG6842 XI11_4/XI0/XI0_53/d_2_ XI11_4/XI0/XI0_53/d__2_ DECAP_INV_G11
XG6843 XI11_4/XI0/XI0_53/d_1_ XI11_4/XI0/XI0_53/d__1_ DECAP_INV_G11
XG6844 XI11_4/XI0/XI0_53/d_0_ XI11_4/XI0/XI0_53/d__0_ DECAP_INV_G11
XG6845 XI11_4/XI0/XI0_52/d__15_ XI11_4/XI0/XI0_52/d_15_ DECAP_INV_G11
XG6846 XI11_4/XI0/XI0_52/d__14_ XI11_4/XI0/XI0_52/d_14_ DECAP_INV_G11
XG6847 XI11_4/XI0/XI0_52/d__13_ XI11_4/XI0/XI0_52/d_13_ DECAP_INV_G11
XG6848 XI11_4/XI0/XI0_52/d__12_ XI11_4/XI0/XI0_52/d_12_ DECAP_INV_G11
XG6849 XI11_4/XI0/XI0_52/d__11_ XI11_4/XI0/XI0_52/d_11_ DECAP_INV_G11
XG6850 XI11_4/XI0/XI0_52/d__10_ XI11_4/XI0/XI0_52/d_10_ DECAP_INV_G11
XG6851 XI11_4/XI0/XI0_52/d__9_ XI11_4/XI0/XI0_52/d_9_ DECAP_INV_G11
XG6852 XI11_4/XI0/XI0_52/d__8_ XI11_4/XI0/XI0_52/d_8_ DECAP_INV_G11
XG6853 XI11_4/XI0/XI0_52/d__7_ XI11_4/XI0/XI0_52/d_7_ DECAP_INV_G11
XG6854 XI11_4/XI0/XI0_52/d__6_ XI11_4/XI0/XI0_52/d_6_ DECAP_INV_G11
XG6855 XI11_4/XI0/XI0_52/d__5_ XI11_4/XI0/XI0_52/d_5_ DECAP_INV_G11
XG6856 XI11_4/XI0/XI0_52/d__4_ XI11_4/XI0/XI0_52/d_4_ DECAP_INV_G11
XG6857 XI11_4/XI0/XI0_52/d__3_ XI11_4/XI0/XI0_52/d_3_ DECAP_INV_G11
XG6858 XI11_4/XI0/XI0_52/d__2_ XI11_4/XI0/XI0_52/d_2_ DECAP_INV_G11
XG6859 XI11_4/XI0/XI0_52/d__1_ XI11_4/XI0/XI0_52/d_1_ DECAP_INV_G11
XG6860 XI11_4/XI0/XI0_52/d__0_ XI11_4/XI0/XI0_52/d_0_ DECAP_INV_G11
XG6861 XI11_4/XI0/XI0_52/d_15_ XI11_4/XI0/XI0_52/d__15_ DECAP_INV_G11
XG6862 XI11_4/XI0/XI0_52/d_14_ XI11_4/XI0/XI0_52/d__14_ DECAP_INV_G11
XG6863 XI11_4/XI0/XI0_52/d_13_ XI11_4/XI0/XI0_52/d__13_ DECAP_INV_G11
XG6864 XI11_4/XI0/XI0_52/d_12_ XI11_4/XI0/XI0_52/d__12_ DECAP_INV_G11
XG6865 XI11_4/XI0/XI0_52/d_11_ XI11_4/XI0/XI0_52/d__11_ DECAP_INV_G11
XG6866 XI11_4/XI0/XI0_52/d_10_ XI11_4/XI0/XI0_52/d__10_ DECAP_INV_G11
XG6867 XI11_4/XI0/XI0_52/d_9_ XI11_4/XI0/XI0_52/d__9_ DECAP_INV_G11
XG6868 XI11_4/XI0/XI0_52/d_8_ XI11_4/XI0/XI0_52/d__8_ DECAP_INV_G11
XG6869 XI11_4/XI0/XI0_52/d_7_ XI11_4/XI0/XI0_52/d__7_ DECAP_INV_G11
XG6870 XI11_4/XI0/XI0_52/d_6_ XI11_4/XI0/XI0_52/d__6_ DECAP_INV_G11
XG6871 XI11_4/XI0/XI0_52/d_5_ XI11_4/XI0/XI0_52/d__5_ DECAP_INV_G11
XG6872 XI11_4/XI0/XI0_52/d_4_ XI11_4/XI0/XI0_52/d__4_ DECAP_INV_G11
XG6873 XI11_4/XI0/XI0_52/d_3_ XI11_4/XI0/XI0_52/d__3_ DECAP_INV_G11
XG6874 XI11_4/XI0/XI0_52/d_2_ XI11_4/XI0/XI0_52/d__2_ DECAP_INV_G11
XG6875 XI11_4/XI0/XI0_52/d_1_ XI11_4/XI0/XI0_52/d__1_ DECAP_INV_G11
XG6876 XI11_4/XI0/XI0_52/d_0_ XI11_4/XI0/XI0_52/d__0_ DECAP_INV_G11
XG6877 XI11_4/XI0/XI0_51/d__15_ XI11_4/XI0/XI0_51/d_15_ DECAP_INV_G11
XG6878 XI11_4/XI0/XI0_51/d__14_ XI11_4/XI0/XI0_51/d_14_ DECAP_INV_G11
XG6879 XI11_4/XI0/XI0_51/d__13_ XI11_4/XI0/XI0_51/d_13_ DECAP_INV_G11
XG6880 XI11_4/XI0/XI0_51/d__12_ XI11_4/XI0/XI0_51/d_12_ DECAP_INV_G11
XG6881 XI11_4/XI0/XI0_51/d__11_ XI11_4/XI0/XI0_51/d_11_ DECAP_INV_G11
XG6882 XI11_4/XI0/XI0_51/d__10_ XI11_4/XI0/XI0_51/d_10_ DECAP_INV_G11
XG6883 XI11_4/XI0/XI0_51/d__9_ XI11_4/XI0/XI0_51/d_9_ DECAP_INV_G11
XG6884 XI11_4/XI0/XI0_51/d__8_ XI11_4/XI0/XI0_51/d_8_ DECAP_INV_G11
XG6885 XI11_4/XI0/XI0_51/d__7_ XI11_4/XI0/XI0_51/d_7_ DECAP_INV_G11
XG6886 XI11_4/XI0/XI0_51/d__6_ XI11_4/XI0/XI0_51/d_6_ DECAP_INV_G11
XG6887 XI11_4/XI0/XI0_51/d__5_ XI11_4/XI0/XI0_51/d_5_ DECAP_INV_G11
XG6888 XI11_4/XI0/XI0_51/d__4_ XI11_4/XI0/XI0_51/d_4_ DECAP_INV_G11
XG6889 XI11_4/XI0/XI0_51/d__3_ XI11_4/XI0/XI0_51/d_3_ DECAP_INV_G11
XG6890 XI11_4/XI0/XI0_51/d__2_ XI11_4/XI0/XI0_51/d_2_ DECAP_INV_G11
XG6891 XI11_4/XI0/XI0_51/d__1_ XI11_4/XI0/XI0_51/d_1_ DECAP_INV_G11
XG6892 XI11_4/XI0/XI0_51/d__0_ XI11_4/XI0/XI0_51/d_0_ DECAP_INV_G11
XG6893 XI11_4/XI0/XI0_51/d_15_ XI11_4/XI0/XI0_51/d__15_ DECAP_INV_G11
XG6894 XI11_4/XI0/XI0_51/d_14_ XI11_4/XI0/XI0_51/d__14_ DECAP_INV_G11
XG6895 XI11_4/XI0/XI0_51/d_13_ XI11_4/XI0/XI0_51/d__13_ DECAP_INV_G11
XG6896 XI11_4/XI0/XI0_51/d_12_ XI11_4/XI0/XI0_51/d__12_ DECAP_INV_G11
XG6897 XI11_4/XI0/XI0_51/d_11_ XI11_4/XI0/XI0_51/d__11_ DECAP_INV_G11
XG6898 XI11_4/XI0/XI0_51/d_10_ XI11_4/XI0/XI0_51/d__10_ DECAP_INV_G11
XG6899 XI11_4/XI0/XI0_51/d_9_ XI11_4/XI0/XI0_51/d__9_ DECAP_INV_G11
XG6900 XI11_4/XI0/XI0_51/d_8_ XI11_4/XI0/XI0_51/d__8_ DECAP_INV_G11
XG6901 XI11_4/XI0/XI0_51/d_7_ XI11_4/XI0/XI0_51/d__7_ DECAP_INV_G11
XG6902 XI11_4/XI0/XI0_51/d_6_ XI11_4/XI0/XI0_51/d__6_ DECAP_INV_G11
XG6903 XI11_4/XI0/XI0_51/d_5_ XI11_4/XI0/XI0_51/d__5_ DECAP_INV_G11
XG6904 XI11_4/XI0/XI0_51/d_4_ XI11_4/XI0/XI0_51/d__4_ DECAP_INV_G11
XG6905 XI11_4/XI0/XI0_51/d_3_ XI11_4/XI0/XI0_51/d__3_ DECAP_INV_G11
XG6906 XI11_4/XI0/XI0_51/d_2_ XI11_4/XI0/XI0_51/d__2_ DECAP_INV_G11
XG6907 XI11_4/XI0/XI0_51/d_1_ XI11_4/XI0/XI0_51/d__1_ DECAP_INV_G11
XG6908 XI11_4/XI0/XI0_51/d_0_ XI11_4/XI0/XI0_51/d__0_ DECAP_INV_G11
XG6909 XI11_4/XI0/XI0_50/d__15_ XI11_4/XI0/XI0_50/d_15_ DECAP_INV_G11
XG6910 XI11_4/XI0/XI0_50/d__14_ XI11_4/XI0/XI0_50/d_14_ DECAP_INV_G11
XG6911 XI11_4/XI0/XI0_50/d__13_ XI11_4/XI0/XI0_50/d_13_ DECAP_INV_G11
XG6912 XI11_4/XI0/XI0_50/d__12_ XI11_4/XI0/XI0_50/d_12_ DECAP_INV_G11
XG6913 XI11_4/XI0/XI0_50/d__11_ XI11_4/XI0/XI0_50/d_11_ DECAP_INV_G11
XG6914 XI11_4/XI0/XI0_50/d__10_ XI11_4/XI0/XI0_50/d_10_ DECAP_INV_G11
XG6915 XI11_4/XI0/XI0_50/d__9_ XI11_4/XI0/XI0_50/d_9_ DECAP_INV_G11
XG6916 XI11_4/XI0/XI0_50/d__8_ XI11_4/XI0/XI0_50/d_8_ DECAP_INV_G11
XG6917 XI11_4/XI0/XI0_50/d__7_ XI11_4/XI0/XI0_50/d_7_ DECAP_INV_G11
XG6918 XI11_4/XI0/XI0_50/d__6_ XI11_4/XI0/XI0_50/d_6_ DECAP_INV_G11
XG6919 XI11_4/XI0/XI0_50/d__5_ XI11_4/XI0/XI0_50/d_5_ DECAP_INV_G11
XG6920 XI11_4/XI0/XI0_50/d__4_ XI11_4/XI0/XI0_50/d_4_ DECAP_INV_G11
XG6921 XI11_4/XI0/XI0_50/d__3_ XI11_4/XI0/XI0_50/d_3_ DECAP_INV_G11
XG6922 XI11_4/XI0/XI0_50/d__2_ XI11_4/XI0/XI0_50/d_2_ DECAP_INV_G11
XG6923 XI11_4/XI0/XI0_50/d__1_ XI11_4/XI0/XI0_50/d_1_ DECAP_INV_G11
XG6924 XI11_4/XI0/XI0_50/d__0_ XI11_4/XI0/XI0_50/d_0_ DECAP_INV_G11
XG6925 XI11_4/XI0/XI0_50/d_15_ XI11_4/XI0/XI0_50/d__15_ DECAP_INV_G11
XG6926 XI11_4/XI0/XI0_50/d_14_ XI11_4/XI0/XI0_50/d__14_ DECAP_INV_G11
XG6927 XI11_4/XI0/XI0_50/d_13_ XI11_4/XI0/XI0_50/d__13_ DECAP_INV_G11
XG6928 XI11_4/XI0/XI0_50/d_12_ XI11_4/XI0/XI0_50/d__12_ DECAP_INV_G11
XG6929 XI11_4/XI0/XI0_50/d_11_ XI11_4/XI0/XI0_50/d__11_ DECAP_INV_G11
XG6930 XI11_4/XI0/XI0_50/d_10_ XI11_4/XI0/XI0_50/d__10_ DECAP_INV_G11
XG6931 XI11_4/XI0/XI0_50/d_9_ XI11_4/XI0/XI0_50/d__9_ DECAP_INV_G11
XG6932 XI11_4/XI0/XI0_50/d_8_ XI11_4/XI0/XI0_50/d__8_ DECAP_INV_G11
XG6933 XI11_4/XI0/XI0_50/d_7_ XI11_4/XI0/XI0_50/d__7_ DECAP_INV_G11
XG6934 XI11_4/XI0/XI0_50/d_6_ XI11_4/XI0/XI0_50/d__6_ DECAP_INV_G11
XG6935 XI11_4/XI0/XI0_50/d_5_ XI11_4/XI0/XI0_50/d__5_ DECAP_INV_G11
XG6936 XI11_4/XI0/XI0_50/d_4_ XI11_4/XI0/XI0_50/d__4_ DECAP_INV_G11
XG6937 XI11_4/XI0/XI0_50/d_3_ XI11_4/XI0/XI0_50/d__3_ DECAP_INV_G11
XG6938 XI11_4/XI0/XI0_50/d_2_ XI11_4/XI0/XI0_50/d__2_ DECAP_INV_G11
XG6939 XI11_4/XI0/XI0_50/d_1_ XI11_4/XI0/XI0_50/d__1_ DECAP_INV_G11
XG6940 XI11_4/XI0/XI0_50/d_0_ XI11_4/XI0/XI0_50/d__0_ DECAP_INV_G11
XG6941 XI11_4/XI0/XI0_49/d__15_ XI11_4/XI0/XI0_49/d_15_ DECAP_INV_G11
XG6942 XI11_4/XI0/XI0_49/d__14_ XI11_4/XI0/XI0_49/d_14_ DECAP_INV_G11
XG6943 XI11_4/XI0/XI0_49/d__13_ XI11_4/XI0/XI0_49/d_13_ DECAP_INV_G11
XG6944 XI11_4/XI0/XI0_49/d__12_ XI11_4/XI0/XI0_49/d_12_ DECAP_INV_G11
XG6945 XI11_4/XI0/XI0_49/d__11_ XI11_4/XI0/XI0_49/d_11_ DECAP_INV_G11
XG6946 XI11_4/XI0/XI0_49/d__10_ XI11_4/XI0/XI0_49/d_10_ DECAP_INV_G11
XG6947 XI11_4/XI0/XI0_49/d__9_ XI11_4/XI0/XI0_49/d_9_ DECAP_INV_G11
XG6948 XI11_4/XI0/XI0_49/d__8_ XI11_4/XI0/XI0_49/d_8_ DECAP_INV_G11
XG6949 XI11_4/XI0/XI0_49/d__7_ XI11_4/XI0/XI0_49/d_7_ DECAP_INV_G11
XG6950 XI11_4/XI0/XI0_49/d__6_ XI11_4/XI0/XI0_49/d_6_ DECAP_INV_G11
XG6951 XI11_4/XI0/XI0_49/d__5_ XI11_4/XI0/XI0_49/d_5_ DECAP_INV_G11
XG6952 XI11_4/XI0/XI0_49/d__4_ XI11_4/XI0/XI0_49/d_4_ DECAP_INV_G11
XG6953 XI11_4/XI0/XI0_49/d__3_ XI11_4/XI0/XI0_49/d_3_ DECAP_INV_G11
XG6954 XI11_4/XI0/XI0_49/d__2_ XI11_4/XI0/XI0_49/d_2_ DECAP_INV_G11
XG6955 XI11_4/XI0/XI0_49/d__1_ XI11_4/XI0/XI0_49/d_1_ DECAP_INV_G11
XG6956 XI11_4/XI0/XI0_49/d__0_ XI11_4/XI0/XI0_49/d_0_ DECAP_INV_G11
XG6957 XI11_4/XI0/XI0_49/d_15_ XI11_4/XI0/XI0_49/d__15_ DECAP_INV_G11
XG6958 XI11_4/XI0/XI0_49/d_14_ XI11_4/XI0/XI0_49/d__14_ DECAP_INV_G11
XG6959 XI11_4/XI0/XI0_49/d_13_ XI11_4/XI0/XI0_49/d__13_ DECAP_INV_G11
XG6960 XI11_4/XI0/XI0_49/d_12_ XI11_4/XI0/XI0_49/d__12_ DECAP_INV_G11
XG6961 XI11_4/XI0/XI0_49/d_11_ XI11_4/XI0/XI0_49/d__11_ DECAP_INV_G11
XG6962 XI11_4/XI0/XI0_49/d_10_ XI11_4/XI0/XI0_49/d__10_ DECAP_INV_G11
XG6963 XI11_4/XI0/XI0_49/d_9_ XI11_4/XI0/XI0_49/d__9_ DECAP_INV_G11
XG6964 XI11_4/XI0/XI0_49/d_8_ XI11_4/XI0/XI0_49/d__8_ DECAP_INV_G11
XG6965 XI11_4/XI0/XI0_49/d_7_ XI11_4/XI0/XI0_49/d__7_ DECAP_INV_G11
XG6966 XI11_4/XI0/XI0_49/d_6_ XI11_4/XI0/XI0_49/d__6_ DECAP_INV_G11
XG6967 XI11_4/XI0/XI0_49/d_5_ XI11_4/XI0/XI0_49/d__5_ DECAP_INV_G11
XG6968 XI11_4/XI0/XI0_49/d_4_ XI11_4/XI0/XI0_49/d__4_ DECAP_INV_G11
XG6969 XI11_4/XI0/XI0_49/d_3_ XI11_4/XI0/XI0_49/d__3_ DECAP_INV_G11
XG6970 XI11_4/XI0/XI0_49/d_2_ XI11_4/XI0/XI0_49/d__2_ DECAP_INV_G11
XG6971 XI11_4/XI0/XI0_49/d_1_ XI11_4/XI0/XI0_49/d__1_ DECAP_INV_G11
XG6972 XI11_4/XI0/XI0_49/d_0_ XI11_4/XI0/XI0_49/d__0_ DECAP_INV_G11
XG6973 XI11_4/XI0/XI0_48/d__15_ XI11_4/XI0/XI0_48/d_15_ DECAP_INV_G11
XG6974 XI11_4/XI0/XI0_48/d__14_ XI11_4/XI0/XI0_48/d_14_ DECAP_INV_G11
XG6975 XI11_4/XI0/XI0_48/d__13_ XI11_4/XI0/XI0_48/d_13_ DECAP_INV_G11
XG6976 XI11_4/XI0/XI0_48/d__12_ XI11_4/XI0/XI0_48/d_12_ DECAP_INV_G11
XG6977 XI11_4/XI0/XI0_48/d__11_ XI11_4/XI0/XI0_48/d_11_ DECAP_INV_G11
XG6978 XI11_4/XI0/XI0_48/d__10_ XI11_4/XI0/XI0_48/d_10_ DECAP_INV_G11
XG6979 XI11_4/XI0/XI0_48/d__9_ XI11_4/XI0/XI0_48/d_9_ DECAP_INV_G11
XG6980 XI11_4/XI0/XI0_48/d__8_ XI11_4/XI0/XI0_48/d_8_ DECAP_INV_G11
XG6981 XI11_4/XI0/XI0_48/d__7_ XI11_4/XI0/XI0_48/d_7_ DECAP_INV_G11
XG6982 XI11_4/XI0/XI0_48/d__6_ XI11_4/XI0/XI0_48/d_6_ DECAP_INV_G11
XG6983 XI11_4/XI0/XI0_48/d__5_ XI11_4/XI0/XI0_48/d_5_ DECAP_INV_G11
XG6984 XI11_4/XI0/XI0_48/d__4_ XI11_4/XI0/XI0_48/d_4_ DECAP_INV_G11
XG6985 XI11_4/XI0/XI0_48/d__3_ XI11_4/XI0/XI0_48/d_3_ DECAP_INV_G11
XG6986 XI11_4/XI0/XI0_48/d__2_ XI11_4/XI0/XI0_48/d_2_ DECAP_INV_G11
XG6987 XI11_4/XI0/XI0_48/d__1_ XI11_4/XI0/XI0_48/d_1_ DECAP_INV_G11
XG6988 XI11_4/XI0/XI0_48/d__0_ XI11_4/XI0/XI0_48/d_0_ DECAP_INV_G11
XG6989 XI11_4/XI0/XI0_48/d_15_ XI11_4/XI0/XI0_48/d__15_ DECAP_INV_G11
XG6990 XI11_4/XI0/XI0_48/d_14_ XI11_4/XI0/XI0_48/d__14_ DECAP_INV_G11
XG6991 XI11_4/XI0/XI0_48/d_13_ XI11_4/XI0/XI0_48/d__13_ DECAP_INV_G11
XG6992 XI11_4/XI0/XI0_48/d_12_ XI11_4/XI0/XI0_48/d__12_ DECAP_INV_G11
XG6993 XI11_4/XI0/XI0_48/d_11_ XI11_4/XI0/XI0_48/d__11_ DECAP_INV_G11
XG6994 XI11_4/XI0/XI0_48/d_10_ XI11_4/XI0/XI0_48/d__10_ DECAP_INV_G11
XG6995 XI11_4/XI0/XI0_48/d_9_ XI11_4/XI0/XI0_48/d__9_ DECAP_INV_G11
XG6996 XI11_4/XI0/XI0_48/d_8_ XI11_4/XI0/XI0_48/d__8_ DECAP_INV_G11
XG6997 XI11_4/XI0/XI0_48/d_7_ XI11_4/XI0/XI0_48/d__7_ DECAP_INV_G11
XG6998 XI11_4/XI0/XI0_48/d_6_ XI11_4/XI0/XI0_48/d__6_ DECAP_INV_G11
XG6999 XI11_4/XI0/XI0_48/d_5_ XI11_4/XI0/XI0_48/d__5_ DECAP_INV_G11
XG7000 XI11_4/XI0/XI0_48/d_4_ XI11_4/XI0/XI0_48/d__4_ DECAP_INV_G11
XG7001 XI11_4/XI0/XI0_48/d_3_ XI11_4/XI0/XI0_48/d__3_ DECAP_INV_G11
XG7002 XI11_4/XI0/XI0_48/d_2_ XI11_4/XI0/XI0_48/d__2_ DECAP_INV_G11
XG7003 XI11_4/XI0/XI0_48/d_1_ XI11_4/XI0/XI0_48/d__1_ DECAP_INV_G11
XG7004 XI11_4/XI0/XI0_48/d_0_ XI11_4/XI0/XI0_48/d__0_ DECAP_INV_G11
XG7005 XI11_4/XI0/XI0_47/d__15_ XI11_4/XI0/XI0_47/d_15_ DECAP_INV_G11
XG7006 XI11_4/XI0/XI0_47/d__14_ XI11_4/XI0/XI0_47/d_14_ DECAP_INV_G11
XG7007 XI11_4/XI0/XI0_47/d__13_ XI11_4/XI0/XI0_47/d_13_ DECAP_INV_G11
XG7008 XI11_4/XI0/XI0_47/d__12_ XI11_4/XI0/XI0_47/d_12_ DECAP_INV_G11
XG7009 XI11_4/XI0/XI0_47/d__11_ XI11_4/XI0/XI0_47/d_11_ DECAP_INV_G11
XG7010 XI11_4/XI0/XI0_47/d__10_ XI11_4/XI0/XI0_47/d_10_ DECAP_INV_G11
XG7011 XI11_4/XI0/XI0_47/d__9_ XI11_4/XI0/XI0_47/d_9_ DECAP_INV_G11
XG7012 XI11_4/XI0/XI0_47/d__8_ XI11_4/XI0/XI0_47/d_8_ DECAP_INV_G11
XG7013 XI11_4/XI0/XI0_47/d__7_ XI11_4/XI0/XI0_47/d_7_ DECAP_INV_G11
XG7014 XI11_4/XI0/XI0_47/d__6_ XI11_4/XI0/XI0_47/d_6_ DECAP_INV_G11
XG7015 XI11_4/XI0/XI0_47/d__5_ XI11_4/XI0/XI0_47/d_5_ DECAP_INV_G11
XG7016 XI11_4/XI0/XI0_47/d__4_ XI11_4/XI0/XI0_47/d_4_ DECAP_INV_G11
XG7017 XI11_4/XI0/XI0_47/d__3_ XI11_4/XI0/XI0_47/d_3_ DECAP_INV_G11
XG7018 XI11_4/XI0/XI0_47/d__2_ XI11_4/XI0/XI0_47/d_2_ DECAP_INV_G11
XG7019 XI11_4/XI0/XI0_47/d__1_ XI11_4/XI0/XI0_47/d_1_ DECAP_INV_G11
XG7020 XI11_4/XI0/XI0_47/d__0_ XI11_4/XI0/XI0_47/d_0_ DECAP_INV_G11
XG7021 XI11_4/XI0/XI0_47/d_15_ XI11_4/XI0/XI0_47/d__15_ DECAP_INV_G11
XG7022 XI11_4/XI0/XI0_47/d_14_ XI11_4/XI0/XI0_47/d__14_ DECAP_INV_G11
XG7023 XI11_4/XI0/XI0_47/d_13_ XI11_4/XI0/XI0_47/d__13_ DECAP_INV_G11
XG7024 XI11_4/XI0/XI0_47/d_12_ XI11_4/XI0/XI0_47/d__12_ DECAP_INV_G11
XG7025 XI11_4/XI0/XI0_47/d_11_ XI11_4/XI0/XI0_47/d__11_ DECAP_INV_G11
XG7026 XI11_4/XI0/XI0_47/d_10_ XI11_4/XI0/XI0_47/d__10_ DECAP_INV_G11
XG7027 XI11_4/XI0/XI0_47/d_9_ XI11_4/XI0/XI0_47/d__9_ DECAP_INV_G11
XG7028 XI11_4/XI0/XI0_47/d_8_ XI11_4/XI0/XI0_47/d__8_ DECAP_INV_G11
XG7029 XI11_4/XI0/XI0_47/d_7_ XI11_4/XI0/XI0_47/d__7_ DECAP_INV_G11
XG7030 XI11_4/XI0/XI0_47/d_6_ XI11_4/XI0/XI0_47/d__6_ DECAP_INV_G11
XG7031 XI11_4/XI0/XI0_47/d_5_ XI11_4/XI0/XI0_47/d__5_ DECAP_INV_G11
XG7032 XI11_4/XI0/XI0_47/d_4_ XI11_4/XI0/XI0_47/d__4_ DECAP_INV_G11
XG7033 XI11_4/XI0/XI0_47/d_3_ XI11_4/XI0/XI0_47/d__3_ DECAP_INV_G11
XG7034 XI11_4/XI0/XI0_47/d_2_ XI11_4/XI0/XI0_47/d__2_ DECAP_INV_G11
XG7035 XI11_4/XI0/XI0_47/d_1_ XI11_4/XI0/XI0_47/d__1_ DECAP_INV_G11
XG7036 XI11_4/XI0/XI0_47/d_0_ XI11_4/XI0/XI0_47/d__0_ DECAP_INV_G11
XG7037 XI11_4/XI0/XI0_46/d__15_ XI11_4/XI0/XI0_46/d_15_ DECAP_INV_G11
XG7038 XI11_4/XI0/XI0_46/d__14_ XI11_4/XI0/XI0_46/d_14_ DECAP_INV_G11
XG7039 XI11_4/XI0/XI0_46/d__13_ XI11_4/XI0/XI0_46/d_13_ DECAP_INV_G11
XG7040 XI11_4/XI0/XI0_46/d__12_ XI11_4/XI0/XI0_46/d_12_ DECAP_INV_G11
XG7041 XI11_4/XI0/XI0_46/d__11_ XI11_4/XI0/XI0_46/d_11_ DECAP_INV_G11
XG7042 XI11_4/XI0/XI0_46/d__10_ XI11_4/XI0/XI0_46/d_10_ DECAP_INV_G11
XG7043 XI11_4/XI0/XI0_46/d__9_ XI11_4/XI0/XI0_46/d_9_ DECAP_INV_G11
XG7044 XI11_4/XI0/XI0_46/d__8_ XI11_4/XI0/XI0_46/d_8_ DECAP_INV_G11
XG7045 XI11_4/XI0/XI0_46/d__7_ XI11_4/XI0/XI0_46/d_7_ DECAP_INV_G11
XG7046 XI11_4/XI0/XI0_46/d__6_ XI11_4/XI0/XI0_46/d_6_ DECAP_INV_G11
XG7047 XI11_4/XI0/XI0_46/d__5_ XI11_4/XI0/XI0_46/d_5_ DECAP_INV_G11
XG7048 XI11_4/XI0/XI0_46/d__4_ XI11_4/XI0/XI0_46/d_4_ DECAP_INV_G11
XG7049 XI11_4/XI0/XI0_46/d__3_ XI11_4/XI0/XI0_46/d_3_ DECAP_INV_G11
XG7050 XI11_4/XI0/XI0_46/d__2_ XI11_4/XI0/XI0_46/d_2_ DECAP_INV_G11
XG7051 XI11_4/XI0/XI0_46/d__1_ XI11_4/XI0/XI0_46/d_1_ DECAP_INV_G11
XG7052 XI11_4/XI0/XI0_46/d__0_ XI11_4/XI0/XI0_46/d_0_ DECAP_INV_G11
XG7053 XI11_4/XI0/XI0_46/d_15_ XI11_4/XI0/XI0_46/d__15_ DECAP_INV_G11
XG7054 XI11_4/XI0/XI0_46/d_14_ XI11_4/XI0/XI0_46/d__14_ DECAP_INV_G11
XG7055 XI11_4/XI0/XI0_46/d_13_ XI11_4/XI0/XI0_46/d__13_ DECAP_INV_G11
XG7056 XI11_4/XI0/XI0_46/d_12_ XI11_4/XI0/XI0_46/d__12_ DECAP_INV_G11
XG7057 XI11_4/XI0/XI0_46/d_11_ XI11_4/XI0/XI0_46/d__11_ DECAP_INV_G11
XG7058 XI11_4/XI0/XI0_46/d_10_ XI11_4/XI0/XI0_46/d__10_ DECAP_INV_G11
XG7059 XI11_4/XI0/XI0_46/d_9_ XI11_4/XI0/XI0_46/d__9_ DECAP_INV_G11
XG7060 XI11_4/XI0/XI0_46/d_8_ XI11_4/XI0/XI0_46/d__8_ DECAP_INV_G11
XG7061 XI11_4/XI0/XI0_46/d_7_ XI11_4/XI0/XI0_46/d__7_ DECAP_INV_G11
XG7062 XI11_4/XI0/XI0_46/d_6_ XI11_4/XI0/XI0_46/d__6_ DECAP_INV_G11
XG7063 XI11_4/XI0/XI0_46/d_5_ XI11_4/XI0/XI0_46/d__5_ DECAP_INV_G11
XG7064 XI11_4/XI0/XI0_46/d_4_ XI11_4/XI0/XI0_46/d__4_ DECAP_INV_G11
XG7065 XI11_4/XI0/XI0_46/d_3_ XI11_4/XI0/XI0_46/d__3_ DECAP_INV_G11
XG7066 XI11_4/XI0/XI0_46/d_2_ XI11_4/XI0/XI0_46/d__2_ DECAP_INV_G11
XG7067 XI11_4/XI0/XI0_46/d_1_ XI11_4/XI0/XI0_46/d__1_ DECAP_INV_G11
XG7068 XI11_4/XI0/XI0_46/d_0_ XI11_4/XI0/XI0_46/d__0_ DECAP_INV_G11
XG7069 XI11_4/XI0/XI0_45/d__15_ XI11_4/XI0/XI0_45/d_15_ DECAP_INV_G11
XG7070 XI11_4/XI0/XI0_45/d__14_ XI11_4/XI0/XI0_45/d_14_ DECAP_INV_G11
XG7071 XI11_4/XI0/XI0_45/d__13_ XI11_4/XI0/XI0_45/d_13_ DECAP_INV_G11
XG7072 XI11_4/XI0/XI0_45/d__12_ XI11_4/XI0/XI0_45/d_12_ DECAP_INV_G11
XG7073 XI11_4/XI0/XI0_45/d__11_ XI11_4/XI0/XI0_45/d_11_ DECAP_INV_G11
XG7074 XI11_4/XI0/XI0_45/d__10_ XI11_4/XI0/XI0_45/d_10_ DECAP_INV_G11
XG7075 XI11_4/XI0/XI0_45/d__9_ XI11_4/XI0/XI0_45/d_9_ DECAP_INV_G11
XG7076 XI11_4/XI0/XI0_45/d__8_ XI11_4/XI0/XI0_45/d_8_ DECAP_INV_G11
XG7077 XI11_4/XI0/XI0_45/d__7_ XI11_4/XI0/XI0_45/d_7_ DECAP_INV_G11
XG7078 XI11_4/XI0/XI0_45/d__6_ XI11_4/XI0/XI0_45/d_6_ DECAP_INV_G11
XG7079 XI11_4/XI0/XI0_45/d__5_ XI11_4/XI0/XI0_45/d_5_ DECAP_INV_G11
XG7080 XI11_4/XI0/XI0_45/d__4_ XI11_4/XI0/XI0_45/d_4_ DECAP_INV_G11
XG7081 XI11_4/XI0/XI0_45/d__3_ XI11_4/XI0/XI0_45/d_3_ DECAP_INV_G11
XG7082 XI11_4/XI0/XI0_45/d__2_ XI11_4/XI0/XI0_45/d_2_ DECAP_INV_G11
XG7083 XI11_4/XI0/XI0_45/d__1_ XI11_4/XI0/XI0_45/d_1_ DECAP_INV_G11
XG7084 XI11_4/XI0/XI0_45/d__0_ XI11_4/XI0/XI0_45/d_0_ DECAP_INV_G11
XG7085 XI11_4/XI0/XI0_45/d_15_ XI11_4/XI0/XI0_45/d__15_ DECAP_INV_G11
XG7086 XI11_4/XI0/XI0_45/d_14_ XI11_4/XI0/XI0_45/d__14_ DECAP_INV_G11
XG7087 XI11_4/XI0/XI0_45/d_13_ XI11_4/XI0/XI0_45/d__13_ DECAP_INV_G11
XG7088 XI11_4/XI0/XI0_45/d_12_ XI11_4/XI0/XI0_45/d__12_ DECAP_INV_G11
XG7089 XI11_4/XI0/XI0_45/d_11_ XI11_4/XI0/XI0_45/d__11_ DECAP_INV_G11
XG7090 XI11_4/XI0/XI0_45/d_10_ XI11_4/XI0/XI0_45/d__10_ DECAP_INV_G11
XG7091 XI11_4/XI0/XI0_45/d_9_ XI11_4/XI0/XI0_45/d__9_ DECAP_INV_G11
XG7092 XI11_4/XI0/XI0_45/d_8_ XI11_4/XI0/XI0_45/d__8_ DECAP_INV_G11
XG7093 XI11_4/XI0/XI0_45/d_7_ XI11_4/XI0/XI0_45/d__7_ DECAP_INV_G11
XG7094 XI11_4/XI0/XI0_45/d_6_ XI11_4/XI0/XI0_45/d__6_ DECAP_INV_G11
XG7095 XI11_4/XI0/XI0_45/d_5_ XI11_4/XI0/XI0_45/d__5_ DECAP_INV_G11
XG7096 XI11_4/XI0/XI0_45/d_4_ XI11_4/XI0/XI0_45/d__4_ DECAP_INV_G11
XG7097 XI11_4/XI0/XI0_45/d_3_ XI11_4/XI0/XI0_45/d__3_ DECAP_INV_G11
XG7098 XI11_4/XI0/XI0_45/d_2_ XI11_4/XI0/XI0_45/d__2_ DECAP_INV_G11
XG7099 XI11_4/XI0/XI0_45/d_1_ XI11_4/XI0/XI0_45/d__1_ DECAP_INV_G11
XG7100 XI11_4/XI0/XI0_45/d_0_ XI11_4/XI0/XI0_45/d__0_ DECAP_INV_G11
XG7101 XI11_4/XI0/XI0_44/d__15_ XI11_4/XI0/XI0_44/d_15_ DECAP_INV_G11
XG7102 XI11_4/XI0/XI0_44/d__14_ XI11_4/XI0/XI0_44/d_14_ DECAP_INV_G11
XG7103 XI11_4/XI0/XI0_44/d__13_ XI11_4/XI0/XI0_44/d_13_ DECAP_INV_G11
XG7104 XI11_4/XI0/XI0_44/d__12_ XI11_4/XI0/XI0_44/d_12_ DECAP_INV_G11
XG7105 XI11_4/XI0/XI0_44/d__11_ XI11_4/XI0/XI0_44/d_11_ DECAP_INV_G11
XG7106 XI11_4/XI0/XI0_44/d__10_ XI11_4/XI0/XI0_44/d_10_ DECAP_INV_G11
XG7107 XI11_4/XI0/XI0_44/d__9_ XI11_4/XI0/XI0_44/d_9_ DECAP_INV_G11
XG7108 XI11_4/XI0/XI0_44/d__8_ XI11_4/XI0/XI0_44/d_8_ DECAP_INV_G11
XG7109 XI11_4/XI0/XI0_44/d__7_ XI11_4/XI0/XI0_44/d_7_ DECAP_INV_G11
XG7110 XI11_4/XI0/XI0_44/d__6_ XI11_4/XI0/XI0_44/d_6_ DECAP_INV_G11
XG7111 XI11_4/XI0/XI0_44/d__5_ XI11_4/XI0/XI0_44/d_5_ DECAP_INV_G11
XG7112 XI11_4/XI0/XI0_44/d__4_ XI11_4/XI0/XI0_44/d_4_ DECAP_INV_G11
XG7113 XI11_4/XI0/XI0_44/d__3_ XI11_4/XI0/XI0_44/d_3_ DECAP_INV_G11
XG7114 XI11_4/XI0/XI0_44/d__2_ XI11_4/XI0/XI0_44/d_2_ DECAP_INV_G11
XG7115 XI11_4/XI0/XI0_44/d__1_ XI11_4/XI0/XI0_44/d_1_ DECAP_INV_G11
XG7116 XI11_4/XI0/XI0_44/d__0_ XI11_4/XI0/XI0_44/d_0_ DECAP_INV_G11
XG7117 XI11_4/XI0/XI0_44/d_15_ XI11_4/XI0/XI0_44/d__15_ DECAP_INV_G11
XG7118 XI11_4/XI0/XI0_44/d_14_ XI11_4/XI0/XI0_44/d__14_ DECAP_INV_G11
XG7119 XI11_4/XI0/XI0_44/d_13_ XI11_4/XI0/XI0_44/d__13_ DECAP_INV_G11
XG7120 XI11_4/XI0/XI0_44/d_12_ XI11_4/XI0/XI0_44/d__12_ DECAP_INV_G11
XG7121 XI11_4/XI0/XI0_44/d_11_ XI11_4/XI0/XI0_44/d__11_ DECAP_INV_G11
XG7122 XI11_4/XI0/XI0_44/d_10_ XI11_4/XI0/XI0_44/d__10_ DECAP_INV_G11
XG7123 XI11_4/XI0/XI0_44/d_9_ XI11_4/XI0/XI0_44/d__9_ DECAP_INV_G11
XG7124 XI11_4/XI0/XI0_44/d_8_ XI11_4/XI0/XI0_44/d__8_ DECAP_INV_G11
XG7125 XI11_4/XI0/XI0_44/d_7_ XI11_4/XI0/XI0_44/d__7_ DECAP_INV_G11
XG7126 XI11_4/XI0/XI0_44/d_6_ XI11_4/XI0/XI0_44/d__6_ DECAP_INV_G11
XG7127 XI11_4/XI0/XI0_44/d_5_ XI11_4/XI0/XI0_44/d__5_ DECAP_INV_G11
XG7128 XI11_4/XI0/XI0_44/d_4_ XI11_4/XI0/XI0_44/d__4_ DECAP_INV_G11
XG7129 XI11_4/XI0/XI0_44/d_3_ XI11_4/XI0/XI0_44/d__3_ DECAP_INV_G11
XG7130 XI11_4/XI0/XI0_44/d_2_ XI11_4/XI0/XI0_44/d__2_ DECAP_INV_G11
XG7131 XI11_4/XI0/XI0_44/d_1_ XI11_4/XI0/XI0_44/d__1_ DECAP_INV_G11
XG7132 XI11_4/XI0/XI0_44/d_0_ XI11_4/XI0/XI0_44/d__0_ DECAP_INV_G11
XG7133 XI11_4/XI0/XI0_43/d__15_ XI11_4/XI0/XI0_43/d_15_ DECAP_INV_G11
XG7134 XI11_4/XI0/XI0_43/d__14_ XI11_4/XI0/XI0_43/d_14_ DECAP_INV_G11
XG7135 XI11_4/XI0/XI0_43/d__13_ XI11_4/XI0/XI0_43/d_13_ DECAP_INV_G11
XG7136 XI11_4/XI0/XI0_43/d__12_ XI11_4/XI0/XI0_43/d_12_ DECAP_INV_G11
XG7137 XI11_4/XI0/XI0_43/d__11_ XI11_4/XI0/XI0_43/d_11_ DECAP_INV_G11
XG7138 XI11_4/XI0/XI0_43/d__10_ XI11_4/XI0/XI0_43/d_10_ DECAP_INV_G11
XG7139 XI11_4/XI0/XI0_43/d__9_ XI11_4/XI0/XI0_43/d_9_ DECAP_INV_G11
XG7140 XI11_4/XI0/XI0_43/d__8_ XI11_4/XI0/XI0_43/d_8_ DECAP_INV_G11
XG7141 XI11_4/XI0/XI0_43/d__7_ XI11_4/XI0/XI0_43/d_7_ DECAP_INV_G11
XG7142 XI11_4/XI0/XI0_43/d__6_ XI11_4/XI0/XI0_43/d_6_ DECAP_INV_G11
XG7143 XI11_4/XI0/XI0_43/d__5_ XI11_4/XI0/XI0_43/d_5_ DECAP_INV_G11
XG7144 XI11_4/XI0/XI0_43/d__4_ XI11_4/XI0/XI0_43/d_4_ DECAP_INV_G11
XG7145 XI11_4/XI0/XI0_43/d__3_ XI11_4/XI0/XI0_43/d_3_ DECAP_INV_G11
XG7146 XI11_4/XI0/XI0_43/d__2_ XI11_4/XI0/XI0_43/d_2_ DECAP_INV_G11
XG7147 XI11_4/XI0/XI0_43/d__1_ XI11_4/XI0/XI0_43/d_1_ DECAP_INV_G11
XG7148 XI11_4/XI0/XI0_43/d__0_ XI11_4/XI0/XI0_43/d_0_ DECAP_INV_G11
XG7149 XI11_4/XI0/XI0_43/d_15_ XI11_4/XI0/XI0_43/d__15_ DECAP_INV_G11
XG7150 XI11_4/XI0/XI0_43/d_14_ XI11_4/XI0/XI0_43/d__14_ DECAP_INV_G11
XG7151 XI11_4/XI0/XI0_43/d_13_ XI11_4/XI0/XI0_43/d__13_ DECAP_INV_G11
XG7152 XI11_4/XI0/XI0_43/d_12_ XI11_4/XI0/XI0_43/d__12_ DECAP_INV_G11
XG7153 XI11_4/XI0/XI0_43/d_11_ XI11_4/XI0/XI0_43/d__11_ DECAP_INV_G11
XG7154 XI11_4/XI0/XI0_43/d_10_ XI11_4/XI0/XI0_43/d__10_ DECAP_INV_G11
XG7155 XI11_4/XI0/XI0_43/d_9_ XI11_4/XI0/XI0_43/d__9_ DECAP_INV_G11
XG7156 XI11_4/XI0/XI0_43/d_8_ XI11_4/XI0/XI0_43/d__8_ DECAP_INV_G11
XG7157 XI11_4/XI0/XI0_43/d_7_ XI11_4/XI0/XI0_43/d__7_ DECAP_INV_G11
XG7158 XI11_4/XI0/XI0_43/d_6_ XI11_4/XI0/XI0_43/d__6_ DECAP_INV_G11
XG7159 XI11_4/XI0/XI0_43/d_5_ XI11_4/XI0/XI0_43/d__5_ DECAP_INV_G11
XG7160 XI11_4/XI0/XI0_43/d_4_ XI11_4/XI0/XI0_43/d__4_ DECAP_INV_G11
XG7161 XI11_4/XI0/XI0_43/d_3_ XI11_4/XI0/XI0_43/d__3_ DECAP_INV_G11
XG7162 XI11_4/XI0/XI0_43/d_2_ XI11_4/XI0/XI0_43/d__2_ DECAP_INV_G11
XG7163 XI11_4/XI0/XI0_43/d_1_ XI11_4/XI0/XI0_43/d__1_ DECAP_INV_G11
XG7164 XI11_4/XI0/XI0_43/d_0_ XI11_4/XI0/XI0_43/d__0_ DECAP_INV_G11
XG7165 XI11_4/XI0/XI0_42/d__15_ XI11_4/XI0/XI0_42/d_15_ DECAP_INV_G11
XG7166 XI11_4/XI0/XI0_42/d__14_ XI11_4/XI0/XI0_42/d_14_ DECAP_INV_G11
XG7167 XI11_4/XI0/XI0_42/d__13_ XI11_4/XI0/XI0_42/d_13_ DECAP_INV_G11
XG7168 XI11_4/XI0/XI0_42/d__12_ XI11_4/XI0/XI0_42/d_12_ DECAP_INV_G11
XG7169 XI11_4/XI0/XI0_42/d__11_ XI11_4/XI0/XI0_42/d_11_ DECAP_INV_G11
XG7170 XI11_4/XI0/XI0_42/d__10_ XI11_4/XI0/XI0_42/d_10_ DECAP_INV_G11
XG7171 XI11_4/XI0/XI0_42/d__9_ XI11_4/XI0/XI0_42/d_9_ DECAP_INV_G11
XG7172 XI11_4/XI0/XI0_42/d__8_ XI11_4/XI0/XI0_42/d_8_ DECAP_INV_G11
XG7173 XI11_4/XI0/XI0_42/d__7_ XI11_4/XI0/XI0_42/d_7_ DECAP_INV_G11
XG7174 XI11_4/XI0/XI0_42/d__6_ XI11_4/XI0/XI0_42/d_6_ DECAP_INV_G11
XG7175 XI11_4/XI0/XI0_42/d__5_ XI11_4/XI0/XI0_42/d_5_ DECAP_INV_G11
XG7176 XI11_4/XI0/XI0_42/d__4_ XI11_4/XI0/XI0_42/d_4_ DECAP_INV_G11
XG7177 XI11_4/XI0/XI0_42/d__3_ XI11_4/XI0/XI0_42/d_3_ DECAP_INV_G11
XG7178 XI11_4/XI0/XI0_42/d__2_ XI11_4/XI0/XI0_42/d_2_ DECAP_INV_G11
XG7179 XI11_4/XI0/XI0_42/d__1_ XI11_4/XI0/XI0_42/d_1_ DECAP_INV_G11
XG7180 XI11_4/XI0/XI0_42/d__0_ XI11_4/XI0/XI0_42/d_0_ DECAP_INV_G11
XG7181 XI11_4/XI0/XI0_42/d_15_ XI11_4/XI0/XI0_42/d__15_ DECAP_INV_G11
XG7182 XI11_4/XI0/XI0_42/d_14_ XI11_4/XI0/XI0_42/d__14_ DECAP_INV_G11
XG7183 XI11_4/XI0/XI0_42/d_13_ XI11_4/XI0/XI0_42/d__13_ DECAP_INV_G11
XG7184 XI11_4/XI0/XI0_42/d_12_ XI11_4/XI0/XI0_42/d__12_ DECAP_INV_G11
XG7185 XI11_4/XI0/XI0_42/d_11_ XI11_4/XI0/XI0_42/d__11_ DECAP_INV_G11
XG7186 XI11_4/XI0/XI0_42/d_10_ XI11_4/XI0/XI0_42/d__10_ DECAP_INV_G11
XG7187 XI11_4/XI0/XI0_42/d_9_ XI11_4/XI0/XI0_42/d__9_ DECAP_INV_G11
XG7188 XI11_4/XI0/XI0_42/d_8_ XI11_4/XI0/XI0_42/d__8_ DECAP_INV_G11
XG7189 XI11_4/XI0/XI0_42/d_7_ XI11_4/XI0/XI0_42/d__7_ DECAP_INV_G11
XG7190 XI11_4/XI0/XI0_42/d_6_ XI11_4/XI0/XI0_42/d__6_ DECAP_INV_G11
XG7191 XI11_4/XI0/XI0_42/d_5_ XI11_4/XI0/XI0_42/d__5_ DECAP_INV_G11
XG7192 XI11_4/XI0/XI0_42/d_4_ XI11_4/XI0/XI0_42/d__4_ DECAP_INV_G11
XG7193 XI11_4/XI0/XI0_42/d_3_ XI11_4/XI0/XI0_42/d__3_ DECAP_INV_G11
XG7194 XI11_4/XI0/XI0_42/d_2_ XI11_4/XI0/XI0_42/d__2_ DECAP_INV_G11
XG7195 XI11_4/XI0/XI0_42/d_1_ XI11_4/XI0/XI0_42/d__1_ DECAP_INV_G11
XG7196 XI11_4/XI0/XI0_42/d_0_ XI11_4/XI0/XI0_42/d__0_ DECAP_INV_G11
XG7197 XI11_4/XI0/XI0_41/d__15_ XI11_4/XI0/XI0_41/d_15_ DECAP_INV_G11
XG7198 XI11_4/XI0/XI0_41/d__14_ XI11_4/XI0/XI0_41/d_14_ DECAP_INV_G11
XG7199 XI11_4/XI0/XI0_41/d__13_ XI11_4/XI0/XI0_41/d_13_ DECAP_INV_G11
XG7200 XI11_4/XI0/XI0_41/d__12_ XI11_4/XI0/XI0_41/d_12_ DECAP_INV_G11
XG7201 XI11_4/XI0/XI0_41/d__11_ XI11_4/XI0/XI0_41/d_11_ DECAP_INV_G11
XG7202 XI11_4/XI0/XI0_41/d__10_ XI11_4/XI0/XI0_41/d_10_ DECAP_INV_G11
XG7203 XI11_4/XI0/XI0_41/d__9_ XI11_4/XI0/XI0_41/d_9_ DECAP_INV_G11
XG7204 XI11_4/XI0/XI0_41/d__8_ XI11_4/XI0/XI0_41/d_8_ DECAP_INV_G11
XG7205 XI11_4/XI0/XI0_41/d__7_ XI11_4/XI0/XI0_41/d_7_ DECAP_INV_G11
XG7206 XI11_4/XI0/XI0_41/d__6_ XI11_4/XI0/XI0_41/d_6_ DECAP_INV_G11
XG7207 XI11_4/XI0/XI0_41/d__5_ XI11_4/XI0/XI0_41/d_5_ DECAP_INV_G11
XG7208 XI11_4/XI0/XI0_41/d__4_ XI11_4/XI0/XI0_41/d_4_ DECAP_INV_G11
XG7209 XI11_4/XI0/XI0_41/d__3_ XI11_4/XI0/XI0_41/d_3_ DECAP_INV_G11
XG7210 XI11_4/XI0/XI0_41/d__2_ XI11_4/XI0/XI0_41/d_2_ DECAP_INV_G11
XG7211 XI11_4/XI0/XI0_41/d__1_ XI11_4/XI0/XI0_41/d_1_ DECAP_INV_G11
XG7212 XI11_4/XI0/XI0_41/d__0_ XI11_4/XI0/XI0_41/d_0_ DECAP_INV_G11
XG7213 XI11_4/XI0/XI0_41/d_15_ XI11_4/XI0/XI0_41/d__15_ DECAP_INV_G11
XG7214 XI11_4/XI0/XI0_41/d_14_ XI11_4/XI0/XI0_41/d__14_ DECAP_INV_G11
XG7215 XI11_4/XI0/XI0_41/d_13_ XI11_4/XI0/XI0_41/d__13_ DECAP_INV_G11
XG7216 XI11_4/XI0/XI0_41/d_12_ XI11_4/XI0/XI0_41/d__12_ DECAP_INV_G11
XG7217 XI11_4/XI0/XI0_41/d_11_ XI11_4/XI0/XI0_41/d__11_ DECAP_INV_G11
XG7218 XI11_4/XI0/XI0_41/d_10_ XI11_4/XI0/XI0_41/d__10_ DECAP_INV_G11
XG7219 XI11_4/XI0/XI0_41/d_9_ XI11_4/XI0/XI0_41/d__9_ DECAP_INV_G11
XG7220 XI11_4/XI0/XI0_41/d_8_ XI11_4/XI0/XI0_41/d__8_ DECAP_INV_G11
XG7221 XI11_4/XI0/XI0_41/d_7_ XI11_4/XI0/XI0_41/d__7_ DECAP_INV_G11
XG7222 XI11_4/XI0/XI0_41/d_6_ XI11_4/XI0/XI0_41/d__6_ DECAP_INV_G11
XG7223 XI11_4/XI0/XI0_41/d_5_ XI11_4/XI0/XI0_41/d__5_ DECAP_INV_G11
XG7224 XI11_4/XI0/XI0_41/d_4_ XI11_4/XI0/XI0_41/d__4_ DECAP_INV_G11
XG7225 XI11_4/XI0/XI0_41/d_3_ XI11_4/XI0/XI0_41/d__3_ DECAP_INV_G11
XG7226 XI11_4/XI0/XI0_41/d_2_ XI11_4/XI0/XI0_41/d__2_ DECAP_INV_G11
XG7227 XI11_4/XI0/XI0_41/d_1_ XI11_4/XI0/XI0_41/d__1_ DECAP_INV_G11
XG7228 XI11_4/XI0/XI0_41/d_0_ XI11_4/XI0/XI0_41/d__0_ DECAP_INV_G11
XG7229 XI11_4/XI0/XI0_40/d__15_ XI11_4/XI0/XI0_40/d_15_ DECAP_INV_G11
XG7230 XI11_4/XI0/XI0_40/d__14_ XI11_4/XI0/XI0_40/d_14_ DECAP_INV_G11
XG7231 XI11_4/XI0/XI0_40/d__13_ XI11_4/XI0/XI0_40/d_13_ DECAP_INV_G11
XG7232 XI11_4/XI0/XI0_40/d__12_ XI11_4/XI0/XI0_40/d_12_ DECAP_INV_G11
XG7233 XI11_4/XI0/XI0_40/d__11_ XI11_4/XI0/XI0_40/d_11_ DECAP_INV_G11
XG7234 XI11_4/XI0/XI0_40/d__10_ XI11_4/XI0/XI0_40/d_10_ DECAP_INV_G11
XG7235 XI11_4/XI0/XI0_40/d__9_ XI11_4/XI0/XI0_40/d_9_ DECAP_INV_G11
XG7236 XI11_4/XI0/XI0_40/d__8_ XI11_4/XI0/XI0_40/d_8_ DECAP_INV_G11
XG7237 XI11_4/XI0/XI0_40/d__7_ XI11_4/XI0/XI0_40/d_7_ DECAP_INV_G11
XG7238 XI11_4/XI0/XI0_40/d__6_ XI11_4/XI0/XI0_40/d_6_ DECAP_INV_G11
XG7239 XI11_4/XI0/XI0_40/d__5_ XI11_4/XI0/XI0_40/d_5_ DECAP_INV_G11
XG7240 XI11_4/XI0/XI0_40/d__4_ XI11_4/XI0/XI0_40/d_4_ DECAP_INV_G11
XG7241 XI11_4/XI0/XI0_40/d__3_ XI11_4/XI0/XI0_40/d_3_ DECAP_INV_G11
XG7242 XI11_4/XI0/XI0_40/d__2_ XI11_4/XI0/XI0_40/d_2_ DECAP_INV_G11
XG7243 XI11_4/XI0/XI0_40/d__1_ XI11_4/XI0/XI0_40/d_1_ DECAP_INV_G11
XG7244 XI11_4/XI0/XI0_40/d__0_ XI11_4/XI0/XI0_40/d_0_ DECAP_INV_G11
XG7245 XI11_4/XI0/XI0_40/d_15_ XI11_4/XI0/XI0_40/d__15_ DECAP_INV_G11
XG7246 XI11_4/XI0/XI0_40/d_14_ XI11_4/XI0/XI0_40/d__14_ DECAP_INV_G11
XG7247 XI11_4/XI0/XI0_40/d_13_ XI11_4/XI0/XI0_40/d__13_ DECAP_INV_G11
XG7248 XI11_4/XI0/XI0_40/d_12_ XI11_4/XI0/XI0_40/d__12_ DECAP_INV_G11
XG7249 XI11_4/XI0/XI0_40/d_11_ XI11_4/XI0/XI0_40/d__11_ DECAP_INV_G11
XG7250 XI11_4/XI0/XI0_40/d_10_ XI11_4/XI0/XI0_40/d__10_ DECAP_INV_G11
XG7251 XI11_4/XI0/XI0_40/d_9_ XI11_4/XI0/XI0_40/d__9_ DECAP_INV_G11
XG7252 XI11_4/XI0/XI0_40/d_8_ XI11_4/XI0/XI0_40/d__8_ DECAP_INV_G11
XG7253 XI11_4/XI0/XI0_40/d_7_ XI11_4/XI0/XI0_40/d__7_ DECAP_INV_G11
XG7254 XI11_4/XI0/XI0_40/d_6_ XI11_4/XI0/XI0_40/d__6_ DECAP_INV_G11
XG7255 XI11_4/XI0/XI0_40/d_5_ XI11_4/XI0/XI0_40/d__5_ DECAP_INV_G11
XG7256 XI11_4/XI0/XI0_40/d_4_ XI11_4/XI0/XI0_40/d__4_ DECAP_INV_G11
XG7257 XI11_4/XI0/XI0_40/d_3_ XI11_4/XI0/XI0_40/d__3_ DECAP_INV_G11
XG7258 XI11_4/XI0/XI0_40/d_2_ XI11_4/XI0/XI0_40/d__2_ DECAP_INV_G11
XG7259 XI11_4/XI0/XI0_40/d_1_ XI11_4/XI0/XI0_40/d__1_ DECAP_INV_G11
XG7260 XI11_4/XI0/XI0_40/d_0_ XI11_4/XI0/XI0_40/d__0_ DECAP_INV_G11
XG7261 XI11_4/XI0/XI0_39/d__15_ XI11_4/XI0/XI0_39/d_15_ DECAP_INV_G11
XG7262 XI11_4/XI0/XI0_39/d__14_ XI11_4/XI0/XI0_39/d_14_ DECAP_INV_G11
XG7263 XI11_4/XI0/XI0_39/d__13_ XI11_4/XI0/XI0_39/d_13_ DECAP_INV_G11
XG7264 XI11_4/XI0/XI0_39/d__12_ XI11_4/XI0/XI0_39/d_12_ DECAP_INV_G11
XG7265 XI11_4/XI0/XI0_39/d__11_ XI11_4/XI0/XI0_39/d_11_ DECAP_INV_G11
XG7266 XI11_4/XI0/XI0_39/d__10_ XI11_4/XI0/XI0_39/d_10_ DECAP_INV_G11
XG7267 XI11_4/XI0/XI0_39/d__9_ XI11_4/XI0/XI0_39/d_9_ DECAP_INV_G11
XG7268 XI11_4/XI0/XI0_39/d__8_ XI11_4/XI0/XI0_39/d_8_ DECAP_INV_G11
XG7269 XI11_4/XI0/XI0_39/d__7_ XI11_4/XI0/XI0_39/d_7_ DECAP_INV_G11
XG7270 XI11_4/XI0/XI0_39/d__6_ XI11_4/XI0/XI0_39/d_6_ DECAP_INV_G11
XG7271 XI11_4/XI0/XI0_39/d__5_ XI11_4/XI0/XI0_39/d_5_ DECAP_INV_G11
XG7272 XI11_4/XI0/XI0_39/d__4_ XI11_4/XI0/XI0_39/d_4_ DECAP_INV_G11
XG7273 XI11_4/XI0/XI0_39/d__3_ XI11_4/XI0/XI0_39/d_3_ DECAP_INV_G11
XG7274 XI11_4/XI0/XI0_39/d__2_ XI11_4/XI0/XI0_39/d_2_ DECAP_INV_G11
XG7275 XI11_4/XI0/XI0_39/d__1_ XI11_4/XI0/XI0_39/d_1_ DECAP_INV_G11
XG7276 XI11_4/XI0/XI0_39/d__0_ XI11_4/XI0/XI0_39/d_0_ DECAP_INV_G11
XG7277 XI11_4/XI0/XI0_39/d_15_ XI11_4/XI0/XI0_39/d__15_ DECAP_INV_G11
XG7278 XI11_4/XI0/XI0_39/d_14_ XI11_4/XI0/XI0_39/d__14_ DECAP_INV_G11
XG7279 XI11_4/XI0/XI0_39/d_13_ XI11_4/XI0/XI0_39/d__13_ DECAP_INV_G11
XG7280 XI11_4/XI0/XI0_39/d_12_ XI11_4/XI0/XI0_39/d__12_ DECAP_INV_G11
XG7281 XI11_4/XI0/XI0_39/d_11_ XI11_4/XI0/XI0_39/d__11_ DECAP_INV_G11
XG7282 XI11_4/XI0/XI0_39/d_10_ XI11_4/XI0/XI0_39/d__10_ DECAP_INV_G11
XG7283 XI11_4/XI0/XI0_39/d_9_ XI11_4/XI0/XI0_39/d__9_ DECAP_INV_G11
XG7284 XI11_4/XI0/XI0_39/d_8_ XI11_4/XI0/XI0_39/d__8_ DECAP_INV_G11
XG7285 XI11_4/XI0/XI0_39/d_7_ XI11_4/XI0/XI0_39/d__7_ DECAP_INV_G11
XG7286 XI11_4/XI0/XI0_39/d_6_ XI11_4/XI0/XI0_39/d__6_ DECAP_INV_G11
XG7287 XI11_4/XI0/XI0_39/d_5_ XI11_4/XI0/XI0_39/d__5_ DECAP_INV_G11
XG7288 XI11_4/XI0/XI0_39/d_4_ XI11_4/XI0/XI0_39/d__4_ DECAP_INV_G11
XG7289 XI11_4/XI0/XI0_39/d_3_ XI11_4/XI0/XI0_39/d__3_ DECAP_INV_G11
XG7290 XI11_4/XI0/XI0_39/d_2_ XI11_4/XI0/XI0_39/d__2_ DECAP_INV_G11
XG7291 XI11_4/XI0/XI0_39/d_1_ XI11_4/XI0/XI0_39/d__1_ DECAP_INV_G11
XG7292 XI11_4/XI0/XI0_39/d_0_ XI11_4/XI0/XI0_39/d__0_ DECAP_INV_G11
XG7293 XI11_4/XI0/XI0_38/d__15_ XI11_4/XI0/XI0_38/d_15_ DECAP_INV_G11
XG7294 XI11_4/XI0/XI0_38/d__14_ XI11_4/XI0/XI0_38/d_14_ DECAP_INV_G11
XG7295 XI11_4/XI0/XI0_38/d__13_ XI11_4/XI0/XI0_38/d_13_ DECAP_INV_G11
XG7296 XI11_4/XI0/XI0_38/d__12_ XI11_4/XI0/XI0_38/d_12_ DECAP_INV_G11
XG7297 XI11_4/XI0/XI0_38/d__11_ XI11_4/XI0/XI0_38/d_11_ DECAP_INV_G11
XG7298 XI11_4/XI0/XI0_38/d__10_ XI11_4/XI0/XI0_38/d_10_ DECAP_INV_G11
XG7299 XI11_4/XI0/XI0_38/d__9_ XI11_4/XI0/XI0_38/d_9_ DECAP_INV_G11
XG7300 XI11_4/XI0/XI0_38/d__8_ XI11_4/XI0/XI0_38/d_8_ DECAP_INV_G11
XG7301 XI11_4/XI0/XI0_38/d__7_ XI11_4/XI0/XI0_38/d_7_ DECAP_INV_G11
XG7302 XI11_4/XI0/XI0_38/d__6_ XI11_4/XI0/XI0_38/d_6_ DECAP_INV_G11
XG7303 XI11_4/XI0/XI0_38/d__5_ XI11_4/XI0/XI0_38/d_5_ DECAP_INV_G11
XG7304 XI11_4/XI0/XI0_38/d__4_ XI11_4/XI0/XI0_38/d_4_ DECAP_INV_G11
XG7305 XI11_4/XI0/XI0_38/d__3_ XI11_4/XI0/XI0_38/d_3_ DECAP_INV_G11
XG7306 XI11_4/XI0/XI0_38/d__2_ XI11_4/XI0/XI0_38/d_2_ DECAP_INV_G11
XG7307 XI11_4/XI0/XI0_38/d__1_ XI11_4/XI0/XI0_38/d_1_ DECAP_INV_G11
XG7308 XI11_4/XI0/XI0_38/d__0_ XI11_4/XI0/XI0_38/d_0_ DECAP_INV_G11
XG7309 XI11_4/XI0/XI0_38/d_15_ XI11_4/XI0/XI0_38/d__15_ DECAP_INV_G11
XG7310 XI11_4/XI0/XI0_38/d_14_ XI11_4/XI0/XI0_38/d__14_ DECAP_INV_G11
XG7311 XI11_4/XI0/XI0_38/d_13_ XI11_4/XI0/XI0_38/d__13_ DECAP_INV_G11
XG7312 XI11_4/XI0/XI0_38/d_12_ XI11_4/XI0/XI0_38/d__12_ DECAP_INV_G11
XG7313 XI11_4/XI0/XI0_38/d_11_ XI11_4/XI0/XI0_38/d__11_ DECAP_INV_G11
XG7314 XI11_4/XI0/XI0_38/d_10_ XI11_4/XI0/XI0_38/d__10_ DECAP_INV_G11
XG7315 XI11_4/XI0/XI0_38/d_9_ XI11_4/XI0/XI0_38/d__9_ DECAP_INV_G11
XG7316 XI11_4/XI0/XI0_38/d_8_ XI11_4/XI0/XI0_38/d__8_ DECAP_INV_G11
XG7317 XI11_4/XI0/XI0_38/d_7_ XI11_4/XI0/XI0_38/d__7_ DECAP_INV_G11
XG7318 XI11_4/XI0/XI0_38/d_6_ XI11_4/XI0/XI0_38/d__6_ DECAP_INV_G11
XG7319 XI11_4/XI0/XI0_38/d_5_ XI11_4/XI0/XI0_38/d__5_ DECAP_INV_G11
XG7320 XI11_4/XI0/XI0_38/d_4_ XI11_4/XI0/XI0_38/d__4_ DECAP_INV_G11
XG7321 XI11_4/XI0/XI0_38/d_3_ XI11_4/XI0/XI0_38/d__3_ DECAP_INV_G11
XG7322 XI11_4/XI0/XI0_38/d_2_ XI11_4/XI0/XI0_38/d__2_ DECAP_INV_G11
XG7323 XI11_4/XI0/XI0_38/d_1_ XI11_4/XI0/XI0_38/d__1_ DECAP_INV_G11
XG7324 XI11_4/XI0/XI0_38/d_0_ XI11_4/XI0/XI0_38/d__0_ DECAP_INV_G11
XG7325 XI11_4/XI0/XI0_37/d__15_ XI11_4/XI0/XI0_37/d_15_ DECAP_INV_G11
XG7326 XI11_4/XI0/XI0_37/d__14_ XI11_4/XI0/XI0_37/d_14_ DECAP_INV_G11
XG7327 XI11_4/XI0/XI0_37/d__13_ XI11_4/XI0/XI0_37/d_13_ DECAP_INV_G11
XG7328 XI11_4/XI0/XI0_37/d__12_ XI11_4/XI0/XI0_37/d_12_ DECAP_INV_G11
XG7329 XI11_4/XI0/XI0_37/d__11_ XI11_4/XI0/XI0_37/d_11_ DECAP_INV_G11
XG7330 XI11_4/XI0/XI0_37/d__10_ XI11_4/XI0/XI0_37/d_10_ DECAP_INV_G11
XG7331 XI11_4/XI0/XI0_37/d__9_ XI11_4/XI0/XI0_37/d_9_ DECAP_INV_G11
XG7332 XI11_4/XI0/XI0_37/d__8_ XI11_4/XI0/XI0_37/d_8_ DECAP_INV_G11
XG7333 XI11_4/XI0/XI0_37/d__7_ XI11_4/XI0/XI0_37/d_7_ DECAP_INV_G11
XG7334 XI11_4/XI0/XI0_37/d__6_ XI11_4/XI0/XI0_37/d_6_ DECAP_INV_G11
XG7335 XI11_4/XI0/XI0_37/d__5_ XI11_4/XI0/XI0_37/d_5_ DECAP_INV_G11
XG7336 XI11_4/XI0/XI0_37/d__4_ XI11_4/XI0/XI0_37/d_4_ DECAP_INV_G11
XG7337 XI11_4/XI0/XI0_37/d__3_ XI11_4/XI0/XI0_37/d_3_ DECAP_INV_G11
XG7338 XI11_4/XI0/XI0_37/d__2_ XI11_4/XI0/XI0_37/d_2_ DECAP_INV_G11
XG7339 XI11_4/XI0/XI0_37/d__1_ XI11_4/XI0/XI0_37/d_1_ DECAP_INV_G11
XG7340 XI11_4/XI0/XI0_37/d__0_ XI11_4/XI0/XI0_37/d_0_ DECAP_INV_G11
XG7341 XI11_4/XI0/XI0_37/d_15_ XI11_4/XI0/XI0_37/d__15_ DECAP_INV_G11
XG7342 XI11_4/XI0/XI0_37/d_14_ XI11_4/XI0/XI0_37/d__14_ DECAP_INV_G11
XG7343 XI11_4/XI0/XI0_37/d_13_ XI11_4/XI0/XI0_37/d__13_ DECAP_INV_G11
XG7344 XI11_4/XI0/XI0_37/d_12_ XI11_4/XI0/XI0_37/d__12_ DECAP_INV_G11
XG7345 XI11_4/XI0/XI0_37/d_11_ XI11_4/XI0/XI0_37/d__11_ DECAP_INV_G11
XG7346 XI11_4/XI0/XI0_37/d_10_ XI11_4/XI0/XI0_37/d__10_ DECAP_INV_G11
XG7347 XI11_4/XI0/XI0_37/d_9_ XI11_4/XI0/XI0_37/d__9_ DECAP_INV_G11
XG7348 XI11_4/XI0/XI0_37/d_8_ XI11_4/XI0/XI0_37/d__8_ DECAP_INV_G11
XG7349 XI11_4/XI0/XI0_37/d_7_ XI11_4/XI0/XI0_37/d__7_ DECAP_INV_G11
XG7350 XI11_4/XI0/XI0_37/d_6_ XI11_4/XI0/XI0_37/d__6_ DECAP_INV_G11
XG7351 XI11_4/XI0/XI0_37/d_5_ XI11_4/XI0/XI0_37/d__5_ DECAP_INV_G11
XG7352 XI11_4/XI0/XI0_37/d_4_ XI11_4/XI0/XI0_37/d__4_ DECAP_INV_G11
XG7353 XI11_4/XI0/XI0_37/d_3_ XI11_4/XI0/XI0_37/d__3_ DECAP_INV_G11
XG7354 XI11_4/XI0/XI0_37/d_2_ XI11_4/XI0/XI0_37/d__2_ DECAP_INV_G11
XG7355 XI11_4/XI0/XI0_37/d_1_ XI11_4/XI0/XI0_37/d__1_ DECAP_INV_G11
XG7356 XI11_4/XI0/XI0_37/d_0_ XI11_4/XI0/XI0_37/d__0_ DECAP_INV_G11
XG7357 XI11_4/XI0/XI0_36/d__15_ XI11_4/XI0/XI0_36/d_15_ DECAP_INV_G11
XG7358 XI11_4/XI0/XI0_36/d__14_ XI11_4/XI0/XI0_36/d_14_ DECAP_INV_G11
XG7359 XI11_4/XI0/XI0_36/d__13_ XI11_4/XI0/XI0_36/d_13_ DECAP_INV_G11
XG7360 XI11_4/XI0/XI0_36/d__12_ XI11_4/XI0/XI0_36/d_12_ DECAP_INV_G11
XG7361 XI11_4/XI0/XI0_36/d__11_ XI11_4/XI0/XI0_36/d_11_ DECAP_INV_G11
XG7362 XI11_4/XI0/XI0_36/d__10_ XI11_4/XI0/XI0_36/d_10_ DECAP_INV_G11
XG7363 XI11_4/XI0/XI0_36/d__9_ XI11_4/XI0/XI0_36/d_9_ DECAP_INV_G11
XG7364 XI11_4/XI0/XI0_36/d__8_ XI11_4/XI0/XI0_36/d_8_ DECAP_INV_G11
XG7365 XI11_4/XI0/XI0_36/d__7_ XI11_4/XI0/XI0_36/d_7_ DECAP_INV_G11
XG7366 XI11_4/XI0/XI0_36/d__6_ XI11_4/XI0/XI0_36/d_6_ DECAP_INV_G11
XG7367 XI11_4/XI0/XI0_36/d__5_ XI11_4/XI0/XI0_36/d_5_ DECAP_INV_G11
XG7368 XI11_4/XI0/XI0_36/d__4_ XI11_4/XI0/XI0_36/d_4_ DECAP_INV_G11
XG7369 XI11_4/XI0/XI0_36/d__3_ XI11_4/XI0/XI0_36/d_3_ DECAP_INV_G11
XG7370 XI11_4/XI0/XI0_36/d__2_ XI11_4/XI0/XI0_36/d_2_ DECAP_INV_G11
XG7371 XI11_4/XI0/XI0_36/d__1_ XI11_4/XI0/XI0_36/d_1_ DECAP_INV_G11
XG7372 XI11_4/XI0/XI0_36/d__0_ XI11_4/XI0/XI0_36/d_0_ DECAP_INV_G11
XG7373 XI11_4/XI0/XI0_36/d_15_ XI11_4/XI0/XI0_36/d__15_ DECAP_INV_G11
XG7374 XI11_4/XI0/XI0_36/d_14_ XI11_4/XI0/XI0_36/d__14_ DECAP_INV_G11
XG7375 XI11_4/XI0/XI0_36/d_13_ XI11_4/XI0/XI0_36/d__13_ DECAP_INV_G11
XG7376 XI11_4/XI0/XI0_36/d_12_ XI11_4/XI0/XI0_36/d__12_ DECAP_INV_G11
XG7377 XI11_4/XI0/XI0_36/d_11_ XI11_4/XI0/XI0_36/d__11_ DECAP_INV_G11
XG7378 XI11_4/XI0/XI0_36/d_10_ XI11_4/XI0/XI0_36/d__10_ DECAP_INV_G11
XG7379 XI11_4/XI0/XI0_36/d_9_ XI11_4/XI0/XI0_36/d__9_ DECAP_INV_G11
XG7380 XI11_4/XI0/XI0_36/d_8_ XI11_4/XI0/XI0_36/d__8_ DECAP_INV_G11
XG7381 XI11_4/XI0/XI0_36/d_7_ XI11_4/XI0/XI0_36/d__7_ DECAP_INV_G11
XG7382 XI11_4/XI0/XI0_36/d_6_ XI11_4/XI0/XI0_36/d__6_ DECAP_INV_G11
XG7383 XI11_4/XI0/XI0_36/d_5_ XI11_4/XI0/XI0_36/d__5_ DECAP_INV_G11
XG7384 XI11_4/XI0/XI0_36/d_4_ XI11_4/XI0/XI0_36/d__4_ DECAP_INV_G11
XG7385 XI11_4/XI0/XI0_36/d_3_ XI11_4/XI0/XI0_36/d__3_ DECAP_INV_G11
XG7386 XI11_4/XI0/XI0_36/d_2_ XI11_4/XI0/XI0_36/d__2_ DECAP_INV_G11
XG7387 XI11_4/XI0/XI0_36/d_1_ XI11_4/XI0/XI0_36/d__1_ DECAP_INV_G11
XG7388 XI11_4/XI0/XI0_36/d_0_ XI11_4/XI0/XI0_36/d__0_ DECAP_INV_G11
XG7389 XI11_4/XI0/XI0_35/d__15_ XI11_4/XI0/XI0_35/d_15_ DECAP_INV_G11
XG7390 XI11_4/XI0/XI0_35/d__14_ XI11_4/XI0/XI0_35/d_14_ DECAP_INV_G11
XG7391 XI11_4/XI0/XI0_35/d__13_ XI11_4/XI0/XI0_35/d_13_ DECAP_INV_G11
XG7392 XI11_4/XI0/XI0_35/d__12_ XI11_4/XI0/XI0_35/d_12_ DECAP_INV_G11
XG7393 XI11_4/XI0/XI0_35/d__11_ XI11_4/XI0/XI0_35/d_11_ DECAP_INV_G11
XG7394 XI11_4/XI0/XI0_35/d__10_ XI11_4/XI0/XI0_35/d_10_ DECAP_INV_G11
XG7395 XI11_4/XI0/XI0_35/d__9_ XI11_4/XI0/XI0_35/d_9_ DECAP_INV_G11
XG7396 XI11_4/XI0/XI0_35/d__8_ XI11_4/XI0/XI0_35/d_8_ DECAP_INV_G11
XG7397 XI11_4/XI0/XI0_35/d__7_ XI11_4/XI0/XI0_35/d_7_ DECAP_INV_G11
XG7398 XI11_4/XI0/XI0_35/d__6_ XI11_4/XI0/XI0_35/d_6_ DECAP_INV_G11
XG7399 XI11_4/XI0/XI0_35/d__5_ XI11_4/XI0/XI0_35/d_5_ DECAP_INV_G11
XG7400 XI11_4/XI0/XI0_35/d__4_ XI11_4/XI0/XI0_35/d_4_ DECAP_INV_G11
XG7401 XI11_4/XI0/XI0_35/d__3_ XI11_4/XI0/XI0_35/d_3_ DECAP_INV_G11
XG7402 XI11_4/XI0/XI0_35/d__2_ XI11_4/XI0/XI0_35/d_2_ DECAP_INV_G11
XG7403 XI11_4/XI0/XI0_35/d__1_ XI11_4/XI0/XI0_35/d_1_ DECAP_INV_G11
XG7404 XI11_4/XI0/XI0_35/d__0_ XI11_4/XI0/XI0_35/d_0_ DECAP_INV_G11
XG7405 XI11_4/XI0/XI0_35/d_15_ XI11_4/XI0/XI0_35/d__15_ DECAP_INV_G11
XG7406 XI11_4/XI0/XI0_35/d_14_ XI11_4/XI0/XI0_35/d__14_ DECAP_INV_G11
XG7407 XI11_4/XI0/XI0_35/d_13_ XI11_4/XI0/XI0_35/d__13_ DECAP_INV_G11
XG7408 XI11_4/XI0/XI0_35/d_12_ XI11_4/XI0/XI0_35/d__12_ DECAP_INV_G11
XG7409 XI11_4/XI0/XI0_35/d_11_ XI11_4/XI0/XI0_35/d__11_ DECAP_INV_G11
XG7410 XI11_4/XI0/XI0_35/d_10_ XI11_4/XI0/XI0_35/d__10_ DECAP_INV_G11
XG7411 XI11_4/XI0/XI0_35/d_9_ XI11_4/XI0/XI0_35/d__9_ DECAP_INV_G11
XG7412 XI11_4/XI0/XI0_35/d_8_ XI11_4/XI0/XI0_35/d__8_ DECAP_INV_G11
XG7413 XI11_4/XI0/XI0_35/d_7_ XI11_4/XI0/XI0_35/d__7_ DECAP_INV_G11
XG7414 XI11_4/XI0/XI0_35/d_6_ XI11_4/XI0/XI0_35/d__6_ DECAP_INV_G11
XG7415 XI11_4/XI0/XI0_35/d_5_ XI11_4/XI0/XI0_35/d__5_ DECAP_INV_G11
XG7416 XI11_4/XI0/XI0_35/d_4_ XI11_4/XI0/XI0_35/d__4_ DECAP_INV_G11
XG7417 XI11_4/XI0/XI0_35/d_3_ XI11_4/XI0/XI0_35/d__3_ DECAP_INV_G11
XG7418 XI11_4/XI0/XI0_35/d_2_ XI11_4/XI0/XI0_35/d__2_ DECAP_INV_G11
XG7419 XI11_4/XI0/XI0_35/d_1_ XI11_4/XI0/XI0_35/d__1_ DECAP_INV_G11
XG7420 XI11_4/XI0/XI0_35/d_0_ XI11_4/XI0/XI0_35/d__0_ DECAP_INV_G11
XG7421 XI11_4/XI0/XI0_34/d__15_ XI11_4/XI0/XI0_34/d_15_ DECAP_INV_G11
XG7422 XI11_4/XI0/XI0_34/d__14_ XI11_4/XI0/XI0_34/d_14_ DECAP_INV_G11
XG7423 XI11_4/XI0/XI0_34/d__13_ XI11_4/XI0/XI0_34/d_13_ DECAP_INV_G11
XG7424 XI11_4/XI0/XI0_34/d__12_ XI11_4/XI0/XI0_34/d_12_ DECAP_INV_G11
XG7425 XI11_4/XI0/XI0_34/d__11_ XI11_4/XI0/XI0_34/d_11_ DECAP_INV_G11
XG7426 XI11_4/XI0/XI0_34/d__10_ XI11_4/XI0/XI0_34/d_10_ DECAP_INV_G11
XG7427 XI11_4/XI0/XI0_34/d__9_ XI11_4/XI0/XI0_34/d_9_ DECAP_INV_G11
XG7428 XI11_4/XI0/XI0_34/d__8_ XI11_4/XI0/XI0_34/d_8_ DECAP_INV_G11
XG7429 XI11_4/XI0/XI0_34/d__7_ XI11_4/XI0/XI0_34/d_7_ DECAP_INV_G11
XG7430 XI11_4/XI0/XI0_34/d__6_ XI11_4/XI0/XI0_34/d_6_ DECAP_INV_G11
XG7431 XI11_4/XI0/XI0_34/d__5_ XI11_4/XI0/XI0_34/d_5_ DECAP_INV_G11
XG7432 XI11_4/XI0/XI0_34/d__4_ XI11_4/XI0/XI0_34/d_4_ DECAP_INV_G11
XG7433 XI11_4/XI0/XI0_34/d__3_ XI11_4/XI0/XI0_34/d_3_ DECAP_INV_G11
XG7434 XI11_4/XI0/XI0_34/d__2_ XI11_4/XI0/XI0_34/d_2_ DECAP_INV_G11
XG7435 XI11_4/XI0/XI0_34/d__1_ XI11_4/XI0/XI0_34/d_1_ DECAP_INV_G11
XG7436 XI11_4/XI0/XI0_34/d__0_ XI11_4/XI0/XI0_34/d_0_ DECAP_INV_G11
XG7437 XI11_4/XI0/XI0_34/d_15_ XI11_4/XI0/XI0_34/d__15_ DECAP_INV_G11
XG7438 XI11_4/XI0/XI0_34/d_14_ XI11_4/XI0/XI0_34/d__14_ DECAP_INV_G11
XG7439 XI11_4/XI0/XI0_34/d_13_ XI11_4/XI0/XI0_34/d__13_ DECAP_INV_G11
XG7440 XI11_4/XI0/XI0_34/d_12_ XI11_4/XI0/XI0_34/d__12_ DECAP_INV_G11
XG7441 XI11_4/XI0/XI0_34/d_11_ XI11_4/XI0/XI0_34/d__11_ DECAP_INV_G11
XG7442 XI11_4/XI0/XI0_34/d_10_ XI11_4/XI0/XI0_34/d__10_ DECAP_INV_G11
XG7443 XI11_4/XI0/XI0_34/d_9_ XI11_4/XI0/XI0_34/d__9_ DECAP_INV_G11
XG7444 XI11_4/XI0/XI0_34/d_8_ XI11_4/XI0/XI0_34/d__8_ DECAP_INV_G11
XG7445 XI11_4/XI0/XI0_34/d_7_ XI11_4/XI0/XI0_34/d__7_ DECAP_INV_G11
XG7446 XI11_4/XI0/XI0_34/d_6_ XI11_4/XI0/XI0_34/d__6_ DECAP_INV_G11
XG7447 XI11_4/XI0/XI0_34/d_5_ XI11_4/XI0/XI0_34/d__5_ DECAP_INV_G11
XG7448 XI11_4/XI0/XI0_34/d_4_ XI11_4/XI0/XI0_34/d__4_ DECAP_INV_G11
XG7449 XI11_4/XI0/XI0_34/d_3_ XI11_4/XI0/XI0_34/d__3_ DECAP_INV_G11
XG7450 XI11_4/XI0/XI0_34/d_2_ XI11_4/XI0/XI0_34/d__2_ DECAP_INV_G11
XG7451 XI11_4/XI0/XI0_34/d_1_ XI11_4/XI0/XI0_34/d__1_ DECAP_INV_G11
XG7452 XI11_4/XI0/XI0_34/d_0_ XI11_4/XI0/XI0_34/d__0_ DECAP_INV_G11
XG7453 XI11_4/XI0/XI0_33/d__15_ XI11_4/XI0/XI0_33/d_15_ DECAP_INV_G11
XG7454 XI11_4/XI0/XI0_33/d__14_ XI11_4/XI0/XI0_33/d_14_ DECAP_INV_G11
XG7455 XI11_4/XI0/XI0_33/d__13_ XI11_4/XI0/XI0_33/d_13_ DECAP_INV_G11
XG7456 XI11_4/XI0/XI0_33/d__12_ XI11_4/XI0/XI0_33/d_12_ DECAP_INV_G11
XG7457 XI11_4/XI0/XI0_33/d__11_ XI11_4/XI0/XI0_33/d_11_ DECAP_INV_G11
XG7458 XI11_4/XI0/XI0_33/d__10_ XI11_4/XI0/XI0_33/d_10_ DECAP_INV_G11
XG7459 XI11_4/XI0/XI0_33/d__9_ XI11_4/XI0/XI0_33/d_9_ DECAP_INV_G11
XG7460 XI11_4/XI0/XI0_33/d__8_ XI11_4/XI0/XI0_33/d_8_ DECAP_INV_G11
XG7461 XI11_4/XI0/XI0_33/d__7_ XI11_4/XI0/XI0_33/d_7_ DECAP_INV_G11
XG7462 XI11_4/XI0/XI0_33/d__6_ XI11_4/XI0/XI0_33/d_6_ DECAP_INV_G11
XG7463 XI11_4/XI0/XI0_33/d__5_ XI11_4/XI0/XI0_33/d_5_ DECAP_INV_G11
XG7464 XI11_4/XI0/XI0_33/d__4_ XI11_4/XI0/XI0_33/d_4_ DECAP_INV_G11
XG7465 XI11_4/XI0/XI0_33/d__3_ XI11_4/XI0/XI0_33/d_3_ DECAP_INV_G11
XG7466 XI11_4/XI0/XI0_33/d__2_ XI11_4/XI0/XI0_33/d_2_ DECAP_INV_G11
XG7467 XI11_4/XI0/XI0_33/d__1_ XI11_4/XI0/XI0_33/d_1_ DECAP_INV_G11
XG7468 XI11_4/XI0/XI0_33/d__0_ XI11_4/XI0/XI0_33/d_0_ DECAP_INV_G11
XG7469 XI11_4/XI0/XI0_33/d_15_ XI11_4/XI0/XI0_33/d__15_ DECAP_INV_G11
XG7470 XI11_4/XI0/XI0_33/d_14_ XI11_4/XI0/XI0_33/d__14_ DECAP_INV_G11
XG7471 XI11_4/XI0/XI0_33/d_13_ XI11_4/XI0/XI0_33/d__13_ DECAP_INV_G11
XG7472 XI11_4/XI0/XI0_33/d_12_ XI11_4/XI0/XI0_33/d__12_ DECAP_INV_G11
XG7473 XI11_4/XI0/XI0_33/d_11_ XI11_4/XI0/XI0_33/d__11_ DECAP_INV_G11
XG7474 XI11_4/XI0/XI0_33/d_10_ XI11_4/XI0/XI0_33/d__10_ DECAP_INV_G11
XG7475 XI11_4/XI0/XI0_33/d_9_ XI11_4/XI0/XI0_33/d__9_ DECAP_INV_G11
XG7476 XI11_4/XI0/XI0_33/d_8_ XI11_4/XI0/XI0_33/d__8_ DECAP_INV_G11
XG7477 XI11_4/XI0/XI0_33/d_7_ XI11_4/XI0/XI0_33/d__7_ DECAP_INV_G11
XG7478 XI11_4/XI0/XI0_33/d_6_ XI11_4/XI0/XI0_33/d__6_ DECAP_INV_G11
XG7479 XI11_4/XI0/XI0_33/d_5_ XI11_4/XI0/XI0_33/d__5_ DECAP_INV_G11
XG7480 XI11_4/XI0/XI0_33/d_4_ XI11_4/XI0/XI0_33/d__4_ DECAP_INV_G11
XG7481 XI11_4/XI0/XI0_33/d_3_ XI11_4/XI0/XI0_33/d__3_ DECAP_INV_G11
XG7482 XI11_4/XI0/XI0_33/d_2_ XI11_4/XI0/XI0_33/d__2_ DECAP_INV_G11
XG7483 XI11_4/XI0/XI0_33/d_1_ XI11_4/XI0/XI0_33/d__1_ DECAP_INV_G11
XG7484 XI11_4/XI0/XI0_33/d_0_ XI11_4/XI0/XI0_33/d__0_ DECAP_INV_G11
XG7485 XI11_4/XI0/XI0_32/d__15_ XI11_4/XI0/XI0_32/d_15_ DECAP_INV_G11
XG7486 XI11_4/XI0/XI0_32/d__14_ XI11_4/XI0/XI0_32/d_14_ DECAP_INV_G11
XG7487 XI11_4/XI0/XI0_32/d__13_ XI11_4/XI0/XI0_32/d_13_ DECAP_INV_G11
XG7488 XI11_4/XI0/XI0_32/d__12_ XI11_4/XI0/XI0_32/d_12_ DECAP_INV_G11
XG7489 XI11_4/XI0/XI0_32/d__11_ XI11_4/XI0/XI0_32/d_11_ DECAP_INV_G11
XG7490 XI11_4/XI0/XI0_32/d__10_ XI11_4/XI0/XI0_32/d_10_ DECAP_INV_G11
XG7491 XI11_4/XI0/XI0_32/d__9_ XI11_4/XI0/XI0_32/d_9_ DECAP_INV_G11
XG7492 XI11_4/XI0/XI0_32/d__8_ XI11_4/XI0/XI0_32/d_8_ DECAP_INV_G11
XG7493 XI11_4/XI0/XI0_32/d__7_ XI11_4/XI0/XI0_32/d_7_ DECAP_INV_G11
XG7494 XI11_4/XI0/XI0_32/d__6_ XI11_4/XI0/XI0_32/d_6_ DECAP_INV_G11
XG7495 XI11_4/XI0/XI0_32/d__5_ XI11_4/XI0/XI0_32/d_5_ DECAP_INV_G11
XG7496 XI11_4/XI0/XI0_32/d__4_ XI11_4/XI0/XI0_32/d_4_ DECAP_INV_G11
XG7497 XI11_4/XI0/XI0_32/d__3_ XI11_4/XI0/XI0_32/d_3_ DECAP_INV_G11
XG7498 XI11_4/XI0/XI0_32/d__2_ XI11_4/XI0/XI0_32/d_2_ DECAP_INV_G11
XG7499 XI11_4/XI0/XI0_32/d__1_ XI11_4/XI0/XI0_32/d_1_ DECAP_INV_G11
XG7500 XI11_4/XI0/XI0_32/d__0_ XI11_4/XI0/XI0_32/d_0_ DECAP_INV_G11
XG7501 XI11_4/XI0/XI0_32/d_15_ XI11_4/XI0/XI0_32/d__15_ DECAP_INV_G11
XG7502 XI11_4/XI0/XI0_32/d_14_ XI11_4/XI0/XI0_32/d__14_ DECAP_INV_G11
XG7503 XI11_4/XI0/XI0_32/d_13_ XI11_4/XI0/XI0_32/d__13_ DECAP_INV_G11
XG7504 XI11_4/XI0/XI0_32/d_12_ XI11_4/XI0/XI0_32/d__12_ DECAP_INV_G11
XG7505 XI11_4/XI0/XI0_32/d_11_ XI11_4/XI0/XI0_32/d__11_ DECAP_INV_G11
XG7506 XI11_4/XI0/XI0_32/d_10_ XI11_4/XI0/XI0_32/d__10_ DECAP_INV_G11
XG7507 XI11_4/XI0/XI0_32/d_9_ XI11_4/XI0/XI0_32/d__9_ DECAP_INV_G11
XG7508 XI11_4/XI0/XI0_32/d_8_ XI11_4/XI0/XI0_32/d__8_ DECAP_INV_G11
XG7509 XI11_4/XI0/XI0_32/d_7_ XI11_4/XI0/XI0_32/d__7_ DECAP_INV_G11
XG7510 XI11_4/XI0/XI0_32/d_6_ XI11_4/XI0/XI0_32/d__6_ DECAP_INV_G11
XG7511 XI11_4/XI0/XI0_32/d_5_ XI11_4/XI0/XI0_32/d__5_ DECAP_INV_G11
XG7512 XI11_4/XI0/XI0_32/d_4_ XI11_4/XI0/XI0_32/d__4_ DECAP_INV_G11
XG7513 XI11_4/XI0/XI0_32/d_3_ XI11_4/XI0/XI0_32/d__3_ DECAP_INV_G11
XG7514 XI11_4/XI0/XI0_32/d_2_ XI11_4/XI0/XI0_32/d__2_ DECAP_INV_G11
XG7515 XI11_4/XI0/XI0_32/d_1_ XI11_4/XI0/XI0_32/d__1_ DECAP_INV_G11
XG7516 XI11_4/XI0/XI0_32/d_0_ XI11_4/XI0/XI0_32/d__0_ DECAP_INV_G11
XG7517 XI11_4/XI0/XI0_31/d__15_ XI11_4/XI0/XI0_31/d_15_ DECAP_INV_G11
XG7518 XI11_4/XI0/XI0_31/d__14_ XI11_4/XI0/XI0_31/d_14_ DECAP_INV_G11
XG7519 XI11_4/XI0/XI0_31/d__13_ XI11_4/XI0/XI0_31/d_13_ DECAP_INV_G11
XG7520 XI11_4/XI0/XI0_31/d__12_ XI11_4/XI0/XI0_31/d_12_ DECAP_INV_G11
XG7521 XI11_4/XI0/XI0_31/d__11_ XI11_4/XI0/XI0_31/d_11_ DECAP_INV_G11
XG7522 XI11_4/XI0/XI0_31/d__10_ XI11_4/XI0/XI0_31/d_10_ DECAP_INV_G11
XG7523 XI11_4/XI0/XI0_31/d__9_ XI11_4/XI0/XI0_31/d_9_ DECAP_INV_G11
XG7524 XI11_4/XI0/XI0_31/d__8_ XI11_4/XI0/XI0_31/d_8_ DECAP_INV_G11
XG7525 XI11_4/XI0/XI0_31/d__7_ XI11_4/XI0/XI0_31/d_7_ DECAP_INV_G11
XG7526 XI11_4/XI0/XI0_31/d__6_ XI11_4/XI0/XI0_31/d_6_ DECAP_INV_G11
XG7527 XI11_4/XI0/XI0_31/d__5_ XI11_4/XI0/XI0_31/d_5_ DECAP_INV_G11
XG7528 XI11_4/XI0/XI0_31/d__4_ XI11_4/XI0/XI0_31/d_4_ DECAP_INV_G11
XG7529 XI11_4/XI0/XI0_31/d__3_ XI11_4/XI0/XI0_31/d_3_ DECAP_INV_G11
XG7530 XI11_4/XI0/XI0_31/d__2_ XI11_4/XI0/XI0_31/d_2_ DECAP_INV_G11
XG7531 XI11_4/XI0/XI0_31/d__1_ XI11_4/XI0/XI0_31/d_1_ DECAP_INV_G11
XG7532 XI11_4/XI0/XI0_31/d__0_ XI11_4/XI0/XI0_31/d_0_ DECAP_INV_G11
XG7533 XI11_4/XI0/XI0_31/d_15_ XI11_4/XI0/XI0_31/d__15_ DECAP_INV_G11
XG7534 XI11_4/XI0/XI0_31/d_14_ XI11_4/XI0/XI0_31/d__14_ DECAP_INV_G11
XG7535 XI11_4/XI0/XI0_31/d_13_ XI11_4/XI0/XI0_31/d__13_ DECAP_INV_G11
XG7536 XI11_4/XI0/XI0_31/d_12_ XI11_4/XI0/XI0_31/d__12_ DECAP_INV_G11
XG7537 XI11_4/XI0/XI0_31/d_11_ XI11_4/XI0/XI0_31/d__11_ DECAP_INV_G11
XG7538 XI11_4/XI0/XI0_31/d_10_ XI11_4/XI0/XI0_31/d__10_ DECAP_INV_G11
XG7539 XI11_4/XI0/XI0_31/d_9_ XI11_4/XI0/XI0_31/d__9_ DECAP_INV_G11
XG7540 XI11_4/XI0/XI0_31/d_8_ XI11_4/XI0/XI0_31/d__8_ DECAP_INV_G11
XG7541 XI11_4/XI0/XI0_31/d_7_ XI11_4/XI0/XI0_31/d__7_ DECAP_INV_G11
XG7542 XI11_4/XI0/XI0_31/d_6_ XI11_4/XI0/XI0_31/d__6_ DECAP_INV_G11
XG7543 XI11_4/XI0/XI0_31/d_5_ XI11_4/XI0/XI0_31/d__5_ DECAP_INV_G11
XG7544 XI11_4/XI0/XI0_31/d_4_ XI11_4/XI0/XI0_31/d__4_ DECAP_INV_G11
XG7545 XI11_4/XI0/XI0_31/d_3_ XI11_4/XI0/XI0_31/d__3_ DECAP_INV_G11
XG7546 XI11_4/XI0/XI0_31/d_2_ XI11_4/XI0/XI0_31/d__2_ DECAP_INV_G11
XG7547 XI11_4/XI0/XI0_31/d_1_ XI11_4/XI0/XI0_31/d__1_ DECAP_INV_G11
XG7548 XI11_4/XI0/XI0_31/d_0_ XI11_4/XI0/XI0_31/d__0_ DECAP_INV_G11
XG7549 XI11_4/XI0/XI0_30/d__15_ XI11_4/XI0/XI0_30/d_15_ DECAP_INV_G11
XG7550 XI11_4/XI0/XI0_30/d__14_ XI11_4/XI0/XI0_30/d_14_ DECAP_INV_G11
XG7551 XI11_4/XI0/XI0_30/d__13_ XI11_4/XI0/XI0_30/d_13_ DECAP_INV_G11
XG7552 XI11_4/XI0/XI0_30/d__12_ XI11_4/XI0/XI0_30/d_12_ DECAP_INV_G11
XG7553 XI11_4/XI0/XI0_30/d__11_ XI11_4/XI0/XI0_30/d_11_ DECAP_INV_G11
XG7554 XI11_4/XI0/XI0_30/d__10_ XI11_4/XI0/XI0_30/d_10_ DECAP_INV_G11
XG7555 XI11_4/XI0/XI0_30/d__9_ XI11_4/XI0/XI0_30/d_9_ DECAP_INV_G11
XG7556 XI11_4/XI0/XI0_30/d__8_ XI11_4/XI0/XI0_30/d_8_ DECAP_INV_G11
XG7557 XI11_4/XI0/XI0_30/d__7_ XI11_4/XI0/XI0_30/d_7_ DECAP_INV_G11
XG7558 XI11_4/XI0/XI0_30/d__6_ XI11_4/XI0/XI0_30/d_6_ DECAP_INV_G11
XG7559 XI11_4/XI0/XI0_30/d__5_ XI11_4/XI0/XI0_30/d_5_ DECAP_INV_G11
XG7560 XI11_4/XI0/XI0_30/d__4_ XI11_4/XI0/XI0_30/d_4_ DECAP_INV_G11
XG7561 XI11_4/XI0/XI0_30/d__3_ XI11_4/XI0/XI0_30/d_3_ DECAP_INV_G11
XG7562 XI11_4/XI0/XI0_30/d__2_ XI11_4/XI0/XI0_30/d_2_ DECAP_INV_G11
XG7563 XI11_4/XI0/XI0_30/d__1_ XI11_4/XI0/XI0_30/d_1_ DECAP_INV_G11
XG7564 XI11_4/XI0/XI0_30/d__0_ XI11_4/XI0/XI0_30/d_0_ DECAP_INV_G11
XG7565 XI11_4/XI0/XI0_30/d_15_ XI11_4/XI0/XI0_30/d__15_ DECAP_INV_G11
XG7566 XI11_4/XI0/XI0_30/d_14_ XI11_4/XI0/XI0_30/d__14_ DECAP_INV_G11
XG7567 XI11_4/XI0/XI0_30/d_13_ XI11_4/XI0/XI0_30/d__13_ DECAP_INV_G11
XG7568 XI11_4/XI0/XI0_30/d_12_ XI11_4/XI0/XI0_30/d__12_ DECAP_INV_G11
XG7569 XI11_4/XI0/XI0_30/d_11_ XI11_4/XI0/XI0_30/d__11_ DECAP_INV_G11
XG7570 XI11_4/XI0/XI0_30/d_10_ XI11_4/XI0/XI0_30/d__10_ DECAP_INV_G11
XG7571 XI11_4/XI0/XI0_30/d_9_ XI11_4/XI0/XI0_30/d__9_ DECAP_INV_G11
XG7572 XI11_4/XI0/XI0_30/d_8_ XI11_4/XI0/XI0_30/d__8_ DECAP_INV_G11
XG7573 XI11_4/XI0/XI0_30/d_7_ XI11_4/XI0/XI0_30/d__7_ DECAP_INV_G11
XG7574 XI11_4/XI0/XI0_30/d_6_ XI11_4/XI0/XI0_30/d__6_ DECAP_INV_G11
XG7575 XI11_4/XI0/XI0_30/d_5_ XI11_4/XI0/XI0_30/d__5_ DECAP_INV_G11
XG7576 XI11_4/XI0/XI0_30/d_4_ XI11_4/XI0/XI0_30/d__4_ DECAP_INV_G11
XG7577 XI11_4/XI0/XI0_30/d_3_ XI11_4/XI0/XI0_30/d__3_ DECAP_INV_G11
XG7578 XI11_4/XI0/XI0_30/d_2_ XI11_4/XI0/XI0_30/d__2_ DECAP_INV_G11
XG7579 XI11_4/XI0/XI0_30/d_1_ XI11_4/XI0/XI0_30/d__1_ DECAP_INV_G11
XG7580 XI11_4/XI0/XI0_30/d_0_ XI11_4/XI0/XI0_30/d__0_ DECAP_INV_G11
XG7581 XI11_4/XI0/XI0_29/d__15_ XI11_4/XI0/XI0_29/d_15_ DECAP_INV_G11
XG7582 XI11_4/XI0/XI0_29/d__14_ XI11_4/XI0/XI0_29/d_14_ DECAP_INV_G11
XG7583 XI11_4/XI0/XI0_29/d__13_ XI11_4/XI0/XI0_29/d_13_ DECAP_INV_G11
XG7584 XI11_4/XI0/XI0_29/d__12_ XI11_4/XI0/XI0_29/d_12_ DECAP_INV_G11
XG7585 XI11_4/XI0/XI0_29/d__11_ XI11_4/XI0/XI0_29/d_11_ DECAP_INV_G11
XG7586 XI11_4/XI0/XI0_29/d__10_ XI11_4/XI0/XI0_29/d_10_ DECAP_INV_G11
XG7587 XI11_4/XI0/XI0_29/d__9_ XI11_4/XI0/XI0_29/d_9_ DECAP_INV_G11
XG7588 XI11_4/XI0/XI0_29/d__8_ XI11_4/XI0/XI0_29/d_8_ DECAP_INV_G11
XG7589 XI11_4/XI0/XI0_29/d__7_ XI11_4/XI0/XI0_29/d_7_ DECAP_INV_G11
XG7590 XI11_4/XI0/XI0_29/d__6_ XI11_4/XI0/XI0_29/d_6_ DECAP_INV_G11
XG7591 XI11_4/XI0/XI0_29/d__5_ XI11_4/XI0/XI0_29/d_5_ DECAP_INV_G11
XG7592 XI11_4/XI0/XI0_29/d__4_ XI11_4/XI0/XI0_29/d_4_ DECAP_INV_G11
XG7593 XI11_4/XI0/XI0_29/d__3_ XI11_4/XI0/XI0_29/d_3_ DECAP_INV_G11
XG7594 XI11_4/XI0/XI0_29/d__2_ XI11_4/XI0/XI0_29/d_2_ DECAP_INV_G11
XG7595 XI11_4/XI0/XI0_29/d__1_ XI11_4/XI0/XI0_29/d_1_ DECAP_INV_G11
XG7596 XI11_4/XI0/XI0_29/d__0_ XI11_4/XI0/XI0_29/d_0_ DECAP_INV_G11
XG7597 XI11_4/XI0/XI0_29/d_15_ XI11_4/XI0/XI0_29/d__15_ DECAP_INV_G11
XG7598 XI11_4/XI0/XI0_29/d_14_ XI11_4/XI0/XI0_29/d__14_ DECAP_INV_G11
XG7599 XI11_4/XI0/XI0_29/d_13_ XI11_4/XI0/XI0_29/d__13_ DECAP_INV_G11
XG7600 XI11_4/XI0/XI0_29/d_12_ XI11_4/XI0/XI0_29/d__12_ DECAP_INV_G11
XG7601 XI11_4/XI0/XI0_29/d_11_ XI11_4/XI0/XI0_29/d__11_ DECAP_INV_G11
XG7602 XI11_4/XI0/XI0_29/d_10_ XI11_4/XI0/XI0_29/d__10_ DECAP_INV_G11
XG7603 XI11_4/XI0/XI0_29/d_9_ XI11_4/XI0/XI0_29/d__9_ DECAP_INV_G11
XG7604 XI11_4/XI0/XI0_29/d_8_ XI11_4/XI0/XI0_29/d__8_ DECAP_INV_G11
XG7605 XI11_4/XI0/XI0_29/d_7_ XI11_4/XI0/XI0_29/d__7_ DECAP_INV_G11
XG7606 XI11_4/XI0/XI0_29/d_6_ XI11_4/XI0/XI0_29/d__6_ DECAP_INV_G11
XG7607 XI11_4/XI0/XI0_29/d_5_ XI11_4/XI0/XI0_29/d__5_ DECAP_INV_G11
XG7608 XI11_4/XI0/XI0_29/d_4_ XI11_4/XI0/XI0_29/d__4_ DECAP_INV_G11
XG7609 XI11_4/XI0/XI0_29/d_3_ XI11_4/XI0/XI0_29/d__3_ DECAP_INV_G11
XG7610 XI11_4/XI0/XI0_29/d_2_ XI11_4/XI0/XI0_29/d__2_ DECAP_INV_G11
XG7611 XI11_4/XI0/XI0_29/d_1_ XI11_4/XI0/XI0_29/d__1_ DECAP_INV_G11
XG7612 XI11_4/XI0/XI0_29/d_0_ XI11_4/XI0/XI0_29/d__0_ DECAP_INV_G11
XG7613 XI11_4/XI0/XI0_28/d__15_ XI11_4/XI0/XI0_28/d_15_ DECAP_INV_G11
XG7614 XI11_4/XI0/XI0_28/d__14_ XI11_4/XI0/XI0_28/d_14_ DECAP_INV_G11
XG7615 XI11_4/XI0/XI0_28/d__13_ XI11_4/XI0/XI0_28/d_13_ DECAP_INV_G11
XG7616 XI11_4/XI0/XI0_28/d__12_ XI11_4/XI0/XI0_28/d_12_ DECAP_INV_G11
XG7617 XI11_4/XI0/XI0_28/d__11_ XI11_4/XI0/XI0_28/d_11_ DECAP_INV_G11
XG7618 XI11_4/XI0/XI0_28/d__10_ XI11_4/XI0/XI0_28/d_10_ DECAP_INV_G11
XG7619 XI11_4/XI0/XI0_28/d__9_ XI11_4/XI0/XI0_28/d_9_ DECAP_INV_G11
XG7620 XI11_4/XI0/XI0_28/d__8_ XI11_4/XI0/XI0_28/d_8_ DECAP_INV_G11
XG7621 XI11_4/XI0/XI0_28/d__7_ XI11_4/XI0/XI0_28/d_7_ DECAP_INV_G11
XG7622 XI11_4/XI0/XI0_28/d__6_ XI11_4/XI0/XI0_28/d_6_ DECAP_INV_G11
XG7623 XI11_4/XI0/XI0_28/d__5_ XI11_4/XI0/XI0_28/d_5_ DECAP_INV_G11
XG7624 XI11_4/XI0/XI0_28/d__4_ XI11_4/XI0/XI0_28/d_4_ DECAP_INV_G11
XG7625 XI11_4/XI0/XI0_28/d__3_ XI11_4/XI0/XI0_28/d_3_ DECAP_INV_G11
XG7626 XI11_4/XI0/XI0_28/d__2_ XI11_4/XI0/XI0_28/d_2_ DECAP_INV_G11
XG7627 XI11_4/XI0/XI0_28/d__1_ XI11_4/XI0/XI0_28/d_1_ DECAP_INV_G11
XG7628 XI11_4/XI0/XI0_28/d__0_ XI11_4/XI0/XI0_28/d_0_ DECAP_INV_G11
XG7629 XI11_4/XI0/XI0_28/d_15_ XI11_4/XI0/XI0_28/d__15_ DECAP_INV_G11
XG7630 XI11_4/XI0/XI0_28/d_14_ XI11_4/XI0/XI0_28/d__14_ DECAP_INV_G11
XG7631 XI11_4/XI0/XI0_28/d_13_ XI11_4/XI0/XI0_28/d__13_ DECAP_INV_G11
XG7632 XI11_4/XI0/XI0_28/d_12_ XI11_4/XI0/XI0_28/d__12_ DECAP_INV_G11
XG7633 XI11_4/XI0/XI0_28/d_11_ XI11_4/XI0/XI0_28/d__11_ DECAP_INV_G11
XG7634 XI11_4/XI0/XI0_28/d_10_ XI11_4/XI0/XI0_28/d__10_ DECAP_INV_G11
XG7635 XI11_4/XI0/XI0_28/d_9_ XI11_4/XI0/XI0_28/d__9_ DECAP_INV_G11
XG7636 XI11_4/XI0/XI0_28/d_8_ XI11_4/XI0/XI0_28/d__8_ DECAP_INV_G11
XG7637 XI11_4/XI0/XI0_28/d_7_ XI11_4/XI0/XI0_28/d__7_ DECAP_INV_G11
XG7638 XI11_4/XI0/XI0_28/d_6_ XI11_4/XI0/XI0_28/d__6_ DECAP_INV_G11
XG7639 XI11_4/XI0/XI0_28/d_5_ XI11_4/XI0/XI0_28/d__5_ DECAP_INV_G11
XG7640 XI11_4/XI0/XI0_28/d_4_ XI11_4/XI0/XI0_28/d__4_ DECAP_INV_G11
XG7641 XI11_4/XI0/XI0_28/d_3_ XI11_4/XI0/XI0_28/d__3_ DECAP_INV_G11
XG7642 XI11_4/XI0/XI0_28/d_2_ XI11_4/XI0/XI0_28/d__2_ DECAP_INV_G11
XG7643 XI11_4/XI0/XI0_28/d_1_ XI11_4/XI0/XI0_28/d__1_ DECAP_INV_G11
XG7644 XI11_4/XI0/XI0_28/d_0_ XI11_4/XI0/XI0_28/d__0_ DECAP_INV_G11
XG7645 XI11_4/XI0/XI0_27/d__15_ XI11_4/XI0/XI0_27/d_15_ DECAP_INV_G11
XG7646 XI11_4/XI0/XI0_27/d__14_ XI11_4/XI0/XI0_27/d_14_ DECAP_INV_G11
XG7647 XI11_4/XI0/XI0_27/d__13_ XI11_4/XI0/XI0_27/d_13_ DECAP_INV_G11
XG7648 XI11_4/XI0/XI0_27/d__12_ XI11_4/XI0/XI0_27/d_12_ DECAP_INV_G11
XG7649 XI11_4/XI0/XI0_27/d__11_ XI11_4/XI0/XI0_27/d_11_ DECAP_INV_G11
XG7650 XI11_4/XI0/XI0_27/d__10_ XI11_4/XI0/XI0_27/d_10_ DECAP_INV_G11
XG7651 XI11_4/XI0/XI0_27/d__9_ XI11_4/XI0/XI0_27/d_9_ DECAP_INV_G11
XG7652 XI11_4/XI0/XI0_27/d__8_ XI11_4/XI0/XI0_27/d_8_ DECAP_INV_G11
XG7653 XI11_4/XI0/XI0_27/d__7_ XI11_4/XI0/XI0_27/d_7_ DECAP_INV_G11
XG7654 XI11_4/XI0/XI0_27/d__6_ XI11_4/XI0/XI0_27/d_6_ DECAP_INV_G11
XG7655 XI11_4/XI0/XI0_27/d__5_ XI11_4/XI0/XI0_27/d_5_ DECAP_INV_G11
XG7656 XI11_4/XI0/XI0_27/d__4_ XI11_4/XI0/XI0_27/d_4_ DECAP_INV_G11
XG7657 XI11_4/XI0/XI0_27/d__3_ XI11_4/XI0/XI0_27/d_3_ DECAP_INV_G11
XG7658 XI11_4/XI0/XI0_27/d__2_ XI11_4/XI0/XI0_27/d_2_ DECAP_INV_G11
XG7659 XI11_4/XI0/XI0_27/d__1_ XI11_4/XI0/XI0_27/d_1_ DECAP_INV_G11
XG7660 XI11_4/XI0/XI0_27/d__0_ XI11_4/XI0/XI0_27/d_0_ DECAP_INV_G11
XG7661 XI11_4/XI0/XI0_27/d_15_ XI11_4/XI0/XI0_27/d__15_ DECAP_INV_G11
XG7662 XI11_4/XI0/XI0_27/d_14_ XI11_4/XI0/XI0_27/d__14_ DECAP_INV_G11
XG7663 XI11_4/XI0/XI0_27/d_13_ XI11_4/XI0/XI0_27/d__13_ DECAP_INV_G11
XG7664 XI11_4/XI0/XI0_27/d_12_ XI11_4/XI0/XI0_27/d__12_ DECAP_INV_G11
XG7665 XI11_4/XI0/XI0_27/d_11_ XI11_4/XI0/XI0_27/d__11_ DECAP_INV_G11
XG7666 XI11_4/XI0/XI0_27/d_10_ XI11_4/XI0/XI0_27/d__10_ DECAP_INV_G11
XG7667 XI11_4/XI0/XI0_27/d_9_ XI11_4/XI0/XI0_27/d__9_ DECAP_INV_G11
XG7668 XI11_4/XI0/XI0_27/d_8_ XI11_4/XI0/XI0_27/d__8_ DECAP_INV_G11
XG7669 XI11_4/XI0/XI0_27/d_7_ XI11_4/XI0/XI0_27/d__7_ DECAP_INV_G11
XG7670 XI11_4/XI0/XI0_27/d_6_ XI11_4/XI0/XI0_27/d__6_ DECAP_INV_G11
XG7671 XI11_4/XI0/XI0_27/d_5_ XI11_4/XI0/XI0_27/d__5_ DECAP_INV_G11
XG7672 XI11_4/XI0/XI0_27/d_4_ XI11_4/XI0/XI0_27/d__4_ DECAP_INV_G11
XG7673 XI11_4/XI0/XI0_27/d_3_ XI11_4/XI0/XI0_27/d__3_ DECAP_INV_G11
XG7674 XI11_4/XI0/XI0_27/d_2_ XI11_4/XI0/XI0_27/d__2_ DECAP_INV_G11
XG7675 XI11_4/XI0/XI0_27/d_1_ XI11_4/XI0/XI0_27/d__1_ DECAP_INV_G11
XG7676 XI11_4/XI0/XI0_27/d_0_ XI11_4/XI0/XI0_27/d__0_ DECAP_INV_G11
XG7677 XI11_4/XI0/XI0_26/d__15_ XI11_4/XI0/XI0_26/d_15_ DECAP_INV_G11
XG7678 XI11_4/XI0/XI0_26/d__14_ XI11_4/XI0/XI0_26/d_14_ DECAP_INV_G11
XG7679 XI11_4/XI0/XI0_26/d__13_ XI11_4/XI0/XI0_26/d_13_ DECAP_INV_G11
XG7680 XI11_4/XI0/XI0_26/d__12_ XI11_4/XI0/XI0_26/d_12_ DECAP_INV_G11
XG7681 XI11_4/XI0/XI0_26/d__11_ XI11_4/XI0/XI0_26/d_11_ DECAP_INV_G11
XG7682 XI11_4/XI0/XI0_26/d__10_ XI11_4/XI0/XI0_26/d_10_ DECAP_INV_G11
XG7683 XI11_4/XI0/XI0_26/d__9_ XI11_4/XI0/XI0_26/d_9_ DECAP_INV_G11
XG7684 XI11_4/XI0/XI0_26/d__8_ XI11_4/XI0/XI0_26/d_8_ DECAP_INV_G11
XG7685 XI11_4/XI0/XI0_26/d__7_ XI11_4/XI0/XI0_26/d_7_ DECAP_INV_G11
XG7686 XI11_4/XI0/XI0_26/d__6_ XI11_4/XI0/XI0_26/d_6_ DECAP_INV_G11
XG7687 XI11_4/XI0/XI0_26/d__5_ XI11_4/XI0/XI0_26/d_5_ DECAP_INV_G11
XG7688 XI11_4/XI0/XI0_26/d__4_ XI11_4/XI0/XI0_26/d_4_ DECAP_INV_G11
XG7689 XI11_4/XI0/XI0_26/d__3_ XI11_4/XI0/XI0_26/d_3_ DECAP_INV_G11
XG7690 XI11_4/XI0/XI0_26/d__2_ XI11_4/XI0/XI0_26/d_2_ DECAP_INV_G11
XG7691 XI11_4/XI0/XI0_26/d__1_ XI11_4/XI0/XI0_26/d_1_ DECAP_INV_G11
XG7692 XI11_4/XI0/XI0_26/d__0_ XI11_4/XI0/XI0_26/d_0_ DECAP_INV_G11
XG7693 XI11_4/XI0/XI0_26/d_15_ XI11_4/XI0/XI0_26/d__15_ DECAP_INV_G11
XG7694 XI11_4/XI0/XI0_26/d_14_ XI11_4/XI0/XI0_26/d__14_ DECAP_INV_G11
XG7695 XI11_4/XI0/XI0_26/d_13_ XI11_4/XI0/XI0_26/d__13_ DECAP_INV_G11
XG7696 XI11_4/XI0/XI0_26/d_12_ XI11_4/XI0/XI0_26/d__12_ DECAP_INV_G11
XG7697 XI11_4/XI0/XI0_26/d_11_ XI11_4/XI0/XI0_26/d__11_ DECAP_INV_G11
XG7698 XI11_4/XI0/XI0_26/d_10_ XI11_4/XI0/XI0_26/d__10_ DECAP_INV_G11
XG7699 XI11_4/XI0/XI0_26/d_9_ XI11_4/XI0/XI0_26/d__9_ DECAP_INV_G11
XG7700 XI11_4/XI0/XI0_26/d_8_ XI11_4/XI0/XI0_26/d__8_ DECAP_INV_G11
XG7701 XI11_4/XI0/XI0_26/d_7_ XI11_4/XI0/XI0_26/d__7_ DECAP_INV_G11
XG7702 XI11_4/XI0/XI0_26/d_6_ XI11_4/XI0/XI0_26/d__6_ DECAP_INV_G11
XG7703 XI11_4/XI0/XI0_26/d_5_ XI11_4/XI0/XI0_26/d__5_ DECAP_INV_G11
XG7704 XI11_4/XI0/XI0_26/d_4_ XI11_4/XI0/XI0_26/d__4_ DECAP_INV_G11
XG7705 XI11_4/XI0/XI0_26/d_3_ XI11_4/XI0/XI0_26/d__3_ DECAP_INV_G11
XG7706 XI11_4/XI0/XI0_26/d_2_ XI11_4/XI0/XI0_26/d__2_ DECAP_INV_G11
XG7707 XI11_4/XI0/XI0_26/d_1_ XI11_4/XI0/XI0_26/d__1_ DECAP_INV_G11
XG7708 XI11_4/XI0/XI0_26/d_0_ XI11_4/XI0/XI0_26/d__0_ DECAP_INV_G11
XG7709 XI11_4/XI0/XI0_25/d__15_ XI11_4/XI0/XI0_25/d_15_ DECAP_INV_G11
XG7710 XI11_4/XI0/XI0_25/d__14_ XI11_4/XI0/XI0_25/d_14_ DECAP_INV_G11
XG7711 XI11_4/XI0/XI0_25/d__13_ XI11_4/XI0/XI0_25/d_13_ DECAP_INV_G11
XG7712 XI11_4/XI0/XI0_25/d__12_ XI11_4/XI0/XI0_25/d_12_ DECAP_INV_G11
XG7713 XI11_4/XI0/XI0_25/d__11_ XI11_4/XI0/XI0_25/d_11_ DECAP_INV_G11
XG7714 XI11_4/XI0/XI0_25/d__10_ XI11_4/XI0/XI0_25/d_10_ DECAP_INV_G11
XG7715 XI11_4/XI0/XI0_25/d__9_ XI11_4/XI0/XI0_25/d_9_ DECAP_INV_G11
XG7716 XI11_4/XI0/XI0_25/d__8_ XI11_4/XI0/XI0_25/d_8_ DECAP_INV_G11
XG7717 XI11_4/XI0/XI0_25/d__7_ XI11_4/XI0/XI0_25/d_7_ DECAP_INV_G11
XG7718 XI11_4/XI0/XI0_25/d__6_ XI11_4/XI0/XI0_25/d_6_ DECAP_INV_G11
XG7719 XI11_4/XI0/XI0_25/d__5_ XI11_4/XI0/XI0_25/d_5_ DECAP_INV_G11
XG7720 XI11_4/XI0/XI0_25/d__4_ XI11_4/XI0/XI0_25/d_4_ DECAP_INV_G11
XG7721 XI11_4/XI0/XI0_25/d__3_ XI11_4/XI0/XI0_25/d_3_ DECAP_INV_G11
XG7722 XI11_4/XI0/XI0_25/d__2_ XI11_4/XI0/XI0_25/d_2_ DECAP_INV_G11
XG7723 XI11_4/XI0/XI0_25/d__1_ XI11_4/XI0/XI0_25/d_1_ DECAP_INV_G11
XG7724 XI11_4/XI0/XI0_25/d__0_ XI11_4/XI0/XI0_25/d_0_ DECAP_INV_G11
XG7725 XI11_4/XI0/XI0_25/d_15_ XI11_4/XI0/XI0_25/d__15_ DECAP_INV_G11
XG7726 XI11_4/XI0/XI0_25/d_14_ XI11_4/XI0/XI0_25/d__14_ DECAP_INV_G11
XG7727 XI11_4/XI0/XI0_25/d_13_ XI11_4/XI0/XI0_25/d__13_ DECAP_INV_G11
XG7728 XI11_4/XI0/XI0_25/d_12_ XI11_4/XI0/XI0_25/d__12_ DECAP_INV_G11
XG7729 XI11_4/XI0/XI0_25/d_11_ XI11_4/XI0/XI0_25/d__11_ DECAP_INV_G11
XG7730 XI11_4/XI0/XI0_25/d_10_ XI11_4/XI0/XI0_25/d__10_ DECAP_INV_G11
XG7731 XI11_4/XI0/XI0_25/d_9_ XI11_4/XI0/XI0_25/d__9_ DECAP_INV_G11
XG7732 XI11_4/XI0/XI0_25/d_8_ XI11_4/XI0/XI0_25/d__8_ DECAP_INV_G11
XG7733 XI11_4/XI0/XI0_25/d_7_ XI11_4/XI0/XI0_25/d__7_ DECAP_INV_G11
XG7734 XI11_4/XI0/XI0_25/d_6_ XI11_4/XI0/XI0_25/d__6_ DECAP_INV_G11
XG7735 XI11_4/XI0/XI0_25/d_5_ XI11_4/XI0/XI0_25/d__5_ DECAP_INV_G11
XG7736 XI11_4/XI0/XI0_25/d_4_ XI11_4/XI0/XI0_25/d__4_ DECAP_INV_G11
XG7737 XI11_4/XI0/XI0_25/d_3_ XI11_4/XI0/XI0_25/d__3_ DECAP_INV_G11
XG7738 XI11_4/XI0/XI0_25/d_2_ XI11_4/XI0/XI0_25/d__2_ DECAP_INV_G11
XG7739 XI11_4/XI0/XI0_25/d_1_ XI11_4/XI0/XI0_25/d__1_ DECAP_INV_G11
XG7740 XI11_4/XI0/XI0_25/d_0_ XI11_4/XI0/XI0_25/d__0_ DECAP_INV_G11
XG7741 XI11_4/XI0/XI0_24/d__15_ XI11_4/XI0/XI0_24/d_15_ DECAP_INV_G11
XG7742 XI11_4/XI0/XI0_24/d__14_ XI11_4/XI0/XI0_24/d_14_ DECAP_INV_G11
XG7743 XI11_4/XI0/XI0_24/d__13_ XI11_4/XI0/XI0_24/d_13_ DECAP_INV_G11
XG7744 XI11_4/XI0/XI0_24/d__12_ XI11_4/XI0/XI0_24/d_12_ DECAP_INV_G11
XG7745 XI11_4/XI0/XI0_24/d__11_ XI11_4/XI0/XI0_24/d_11_ DECAP_INV_G11
XG7746 XI11_4/XI0/XI0_24/d__10_ XI11_4/XI0/XI0_24/d_10_ DECAP_INV_G11
XG7747 XI11_4/XI0/XI0_24/d__9_ XI11_4/XI0/XI0_24/d_9_ DECAP_INV_G11
XG7748 XI11_4/XI0/XI0_24/d__8_ XI11_4/XI0/XI0_24/d_8_ DECAP_INV_G11
XG7749 XI11_4/XI0/XI0_24/d__7_ XI11_4/XI0/XI0_24/d_7_ DECAP_INV_G11
XG7750 XI11_4/XI0/XI0_24/d__6_ XI11_4/XI0/XI0_24/d_6_ DECAP_INV_G11
XG7751 XI11_4/XI0/XI0_24/d__5_ XI11_4/XI0/XI0_24/d_5_ DECAP_INV_G11
XG7752 XI11_4/XI0/XI0_24/d__4_ XI11_4/XI0/XI0_24/d_4_ DECAP_INV_G11
XG7753 XI11_4/XI0/XI0_24/d__3_ XI11_4/XI0/XI0_24/d_3_ DECAP_INV_G11
XG7754 XI11_4/XI0/XI0_24/d__2_ XI11_4/XI0/XI0_24/d_2_ DECAP_INV_G11
XG7755 XI11_4/XI0/XI0_24/d__1_ XI11_4/XI0/XI0_24/d_1_ DECAP_INV_G11
XG7756 XI11_4/XI0/XI0_24/d__0_ XI11_4/XI0/XI0_24/d_0_ DECAP_INV_G11
XG7757 XI11_4/XI0/XI0_24/d_15_ XI11_4/XI0/XI0_24/d__15_ DECAP_INV_G11
XG7758 XI11_4/XI0/XI0_24/d_14_ XI11_4/XI0/XI0_24/d__14_ DECAP_INV_G11
XG7759 XI11_4/XI0/XI0_24/d_13_ XI11_4/XI0/XI0_24/d__13_ DECAP_INV_G11
XG7760 XI11_4/XI0/XI0_24/d_12_ XI11_4/XI0/XI0_24/d__12_ DECAP_INV_G11
XG7761 XI11_4/XI0/XI0_24/d_11_ XI11_4/XI0/XI0_24/d__11_ DECAP_INV_G11
XG7762 XI11_4/XI0/XI0_24/d_10_ XI11_4/XI0/XI0_24/d__10_ DECAP_INV_G11
XG7763 XI11_4/XI0/XI0_24/d_9_ XI11_4/XI0/XI0_24/d__9_ DECAP_INV_G11
XG7764 XI11_4/XI0/XI0_24/d_8_ XI11_4/XI0/XI0_24/d__8_ DECAP_INV_G11
XG7765 XI11_4/XI0/XI0_24/d_7_ XI11_4/XI0/XI0_24/d__7_ DECAP_INV_G11
XG7766 XI11_4/XI0/XI0_24/d_6_ XI11_4/XI0/XI0_24/d__6_ DECAP_INV_G11
XG7767 XI11_4/XI0/XI0_24/d_5_ XI11_4/XI0/XI0_24/d__5_ DECAP_INV_G11
XG7768 XI11_4/XI0/XI0_24/d_4_ XI11_4/XI0/XI0_24/d__4_ DECAP_INV_G11
XG7769 XI11_4/XI0/XI0_24/d_3_ XI11_4/XI0/XI0_24/d__3_ DECAP_INV_G11
XG7770 XI11_4/XI0/XI0_24/d_2_ XI11_4/XI0/XI0_24/d__2_ DECAP_INV_G11
XG7771 XI11_4/XI0/XI0_24/d_1_ XI11_4/XI0/XI0_24/d__1_ DECAP_INV_G11
XG7772 XI11_4/XI0/XI0_24/d_0_ XI11_4/XI0/XI0_24/d__0_ DECAP_INV_G11
XG7773 XI11_4/XI0/XI0_23/d__15_ XI11_4/XI0/XI0_23/d_15_ DECAP_INV_G11
XG7774 XI11_4/XI0/XI0_23/d__14_ XI11_4/XI0/XI0_23/d_14_ DECAP_INV_G11
XG7775 XI11_4/XI0/XI0_23/d__13_ XI11_4/XI0/XI0_23/d_13_ DECAP_INV_G11
XG7776 XI11_4/XI0/XI0_23/d__12_ XI11_4/XI0/XI0_23/d_12_ DECAP_INV_G11
XG7777 XI11_4/XI0/XI0_23/d__11_ XI11_4/XI0/XI0_23/d_11_ DECAP_INV_G11
XG7778 XI11_4/XI0/XI0_23/d__10_ XI11_4/XI0/XI0_23/d_10_ DECAP_INV_G11
XG7779 XI11_4/XI0/XI0_23/d__9_ XI11_4/XI0/XI0_23/d_9_ DECAP_INV_G11
XG7780 XI11_4/XI0/XI0_23/d__8_ XI11_4/XI0/XI0_23/d_8_ DECAP_INV_G11
XG7781 XI11_4/XI0/XI0_23/d__7_ XI11_4/XI0/XI0_23/d_7_ DECAP_INV_G11
XG7782 XI11_4/XI0/XI0_23/d__6_ XI11_4/XI0/XI0_23/d_6_ DECAP_INV_G11
XG7783 XI11_4/XI0/XI0_23/d__5_ XI11_4/XI0/XI0_23/d_5_ DECAP_INV_G11
XG7784 XI11_4/XI0/XI0_23/d__4_ XI11_4/XI0/XI0_23/d_4_ DECAP_INV_G11
XG7785 XI11_4/XI0/XI0_23/d__3_ XI11_4/XI0/XI0_23/d_3_ DECAP_INV_G11
XG7786 XI11_4/XI0/XI0_23/d__2_ XI11_4/XI0/XI0_23/d_2_ DECAP_INV_G11
XG7787 XI11_4/XI0/XI0_23/d__1_ XI11_4/XI0/XI0_23/d_1_ DECAP_INV_G11
XG7788 XI11_4/XI0/XI0_23/d__0_ XI11_4/XI0/XI0_23/d_0_ DECAP_INV_G11
XG7789 XI11_4/XI0/XI0_23/d_15_ XI11_4/XI0/XI0_23/d__15_ DECAP_INV_G11
XG7790 XI11_4/XI0/XI0_23/d_14_ XI11_4/XI0/XI0_23/d__14_ DECAP_INV_G11
XG7791 XI11_4/XI0/XI0_23/d_13_ XI11_4/XI0/XI0_23/d__13_ DECAP_INV_G11
XG7792 XI11_4/XI0/XI0_23/d_12_ XI11_4/XI0/XI0_23/d__12_ DECAP_INV_G11
XG7793 XI11_4/XI0/XI0_23/d_11_ XI11_4/XI0/XI0_23/d__11_ DECAP_INV_G11
XG7794 XI11_4/XI0/XI0_23/d_10_ XI11_4/XI0/XI0_23/d__10_ DECAP_INV_G11
XG7795 XI11_4/XI0/XI0_23/d_9_ XI11_4/XI0/XI0_23/d__9_ DECAP_INV_G11
XG7796 XI11_4/XI0/XI0_23/d_8_ XI11_4/XI0/XI0_23/d__8_ DECAP_INV_G11
XG7797 XI11_4/XI0/XI0_23/d_7_ XI11_4/XI0/XI0_23/d__7_ DECAP_INV_G11
XG7798 XI11_4/XI0/XI0_23/d_6_ XI11_4/XI0/XI0_23/d__6_ DECAP_INV_G11
XG7799 XI11_4/XI0/XI0_23/d_5_ XI11_4/XI0/XI0_23/d__5_ DECAP_INV_G11
XG7800 XI11_4/XI0/XI0_23/d_4_ XI11_4/XI0/XI0_23/d__4_ DECAP_INV_G11
XG7801 XI11_4/XI0/XI0_23/d_3_ XI11_4/XI0/XI0_23/d__3_ DECAP_INV_G11
XG7802 XI11_4/XI0/XI0_23/d_2_ XI11_4/XI0/XI0_23/d__2_ DECAP_INV_G11
XG7803 XI11_4/XI0/XI0_23/d_1_ XI11_4/XI0/XI0_23/d__1_ DECAP_INV_G11
XG7804 XI11_4/XI0/XI0_23/d_0_ XI11_4/XI0/XI0_23/d__0_ DECAP_INV_G11
XG7805 XI11_4/XI0/XI0_22/d__15_ XI11_4/XI0/XI0_22/d_15_ DECAP_INV_G11
XG7806 XI11_4/XI0/XI0_22/d__14_ XI11_4/XI0/XI0_22/d_14_ DECAP_INV_G11
XG7807 XI11_4/XI0/XI0_22/d__13_ XI11_4/XI0/XI0_22/d_13_ DECAP_INV_G11
XG7808 XI11_4/XI0/XI0_22/d__12_ XI11_4/XI0/XI0_22/d_12_ DECAP_INV_G11
XG7809 XI11_4/XI0/XI0_22/d__11_ XI11_4/XI0/XI0_22/d_11_ DECAP_INV_G11
XG7810 XI11_4/XI0/XI0_22/d__10_ XI11_4/XI0/XI0_22/d_10_ DECAP_INV_G11
XG7811 XI11_4/XI0/XI0_22/d__9_ XI11_4/XI0/XI0_22/d_9_ DECAP_INV_G11
XG7812 XI11_4/XI0/XI0_22/d__8_ XI11_4/XI0/XI0_22/d_8_ DECAP_INV_G11
XG7813 XI11_4/XI0/XI0_22/d__7_ XI11_4/XI0/XI0_22/d_7_ DECAP_INV_G11
XG7814 XI11_4/XI0/XI0_22/d__6_ XI11_4/XI0/XI0_22/d_6_ DECAP_INV_G11
XG7815 XI11_4/XI0/XI0_22/d__5_ XI11_4/XI0/XI0_22/d_5_ DECAP_INV_G11
XG7816 XI11_4/XI0/XI0_22/d__4_ XI11_4/XI0/XI0_22/d_4_ DECAP_INV_G11
XG7817 XI11_4/XI0/XI0_22/d__3_ XI11_4/XI0/XI0_22/d_3_ DECAP_INV_G11
XG7818 XI11_4/XI0/XI0_22/d__2_ XI11_4/XI0/XI0_22/d_2_ DECAP_INV_G11
XG7819 XI11_4/XI0/XI0_22/d__1_ XI11_4/XI0/XI0_22/d_1_ DECAP_INV_G11
XG7820 XI11_4/XI0/XI0_22/d__0_ XI11_4/XI0/XI0_22/d_0_ DECAP_INV_G11
XG7821 XI11_4/XI0/XI0_22/d_15_ XI11_4/XI0/XI0_22/d__15_ DECAP_INV_G11
XG7822 XI11_4/XI0/XI0_22/d_14_ XI11_4/XI0/XI0_22/d__14_ DECAP_INV_G11
XG7823 XI11_4/XI0/XI0_22/d_13_ XI11_4/XI0/XI0_22/d__13_ DECAP_INV_G11
XG7824 XI11_4/XI0/XI0_22/d_12_ XI11_4/XI0/XI0_22/d__12_ DECAP_INV_G11
XG7825 XI11_4/XI0/XI0_22/d_11_ XI11_4/XI0/XI0_22/d__11_ DECAP_INV_G11
XG7826 XI11_4/XI0/XI0_22/d_10_ XI11_4/XI0/XI0_22/d__10_ DECAP_INV_G11
XG7827 XI11_4/XI0/XI0_22/d_9_ XI11_4/XI0/XI0_22/d__9_ DECAP_INV_G11
XG7828 XI11_4/XI0/XI0_22/d_8_ XI11_4/XI0/XI0_22/d__8_ DECAP_INV_G11
XG7829 XI11_4/XI0/XI0_22/d_7_ XI11_4/XI0/XI0_22/d__7_ DECAP_INV_G11
XG7830 XI11_4/XI0/XI0_22/d_6_ XI11_4/XI0/XI0_22/d__6_ DECAP_INV_G11
XG7831 XI11_4/XI0/XI0_22/d_5_ XI11_4/XI0/XI0_22/d__5_ DECAP_INV_G11
XG7832 XI11_4/XI0/XI0_22/d_4_ XI11_4/XI0/XI0_22/d__4_ DECAP_INV_G11
XG7833 XI11_4/XI0/XI0_22/d_3_ XI11_4/XI0/XI0_22/d__3_ DECAP_INV_G11
XG7834 XI11_4/XI0/XI0_22/d_2_ XI11_4/XI0/XI0_22/d__2_ DECAP_INV_G11
XG7835 XI11_4/XI0/XI0_22/d_1_ XI11_4/XI0/XI0_22/d__1_ DECAP_INV_G11
XG7836 XI11_4/XI0/XI0_22/d_0_ XI11_4/XI0/XI0_22/d__0_ DECAP_INV_G11
XG7837 XI11_4/XI0/XI0_21/d__15_ XI11_4/XI0/XI0_21/d_15_ DECAP_INV_G11
XG7838 XI11_4/XI0/XI0_21/d__14_ XI11_4/XI0/XI0_21/d_14_ DECAP_INV_G11
XG7839 XI11_4/XI0/XI0_21/d__13_ XI11_4/XI0/XI0_21/d_13_ DECAP_INV_G11
XG7840 XI11_4/XI0/XI0_21/d__12_ XI11_4/XI0/XI0_21/d_12_ DECAP_INV_G11
XG7841 XI11_4/XI0/XI0_21/d__11_ XI11_4/XI0/XI0_21/d_11_ DECAP_INV_G11
XG7842 XI11_4/XI0/XI0_21/d__10_ XI11_4/XI0/XI0_21/d_10_ DECAP_INV_G11
XG7843 XI11_4/XI0/XI0_21/d__9_ XI11_4/XI0/XI0_21/d_9_ DECAP_INV_G11
XG7844 XI11_4/XI0/XI0_21/d__8_ XI11_4/XI0/XI0_21/d_8_ DECAP_INV_G11
XG7845 XI11_4/XI0/XI0_21/d__7_ XI11_4/XI0/XI0_21/d_7_ DECAP_INV_G11
XG7846 XI11_4/XI0/XI0_21/d__6_ XI11_4/XI0/XI0_21/d_6_ DECAP_INV_G11
XG7847 XI11_4/XI0/XI0_21/d__5_ XI11_4/XI0/XI0_21/d_5_ DECAP_INV_G11
XG7848 XI11_4/XI0/XI0_21/d__4_ XI11_4/XI0/XI0_21/d_4_ DECAP_INV_G11
XG7849 XI11_4/XI0/XI0_21/d__3_ XI11_4/XI0/XI0_21/d_3_ DECAP_INV_G11
XG7850 XI11_4/XI0/XI0_21/d__2_ XI11_4/XI0/XI0_21/d_2_ DECAP_INV_G11
XG7851 XI11_4/XI0/XI0_21/d__1_ XI11_4/XI0/XI0_21/d_1_ DECAP_INV_G11
XG7852 XI11_4/XI0/XI0_21/d__0_ XI11_4/XI0/XI0_21/d_0_ DECAP_INV_G11
XG7853 XI11_4/XI0/XI0_21/d_15_ XI11_4/XI0/XI0_21/d__15_ DECAP_INV_G11
XG7854 XI11_4/XI0/XI0_21/d_14_ XI11_4/XI0/XI0_21/d__14_ DECAP_INV_G11
XG7855 XI11_4/XI0/XI0_21/d_13_ XI11_4/XI0/XI0_21/d__13_ DECAP_INV_G11
XG7856 XI11_4/XI0/XI0_21/d_12_ XI11_4/XI0/XI0_21/d__12_ DECAP_INV_G11
XG7857 XI11_4/XI0/XI0_21/d_11_ XI11_4/XI0/XI0_21/d__11_ DECAP_INV_G11
XG7858 XI11_4/XI0/XI0_21/d_10_ XI11_4/XI0/XI0_21/d__10_ DECAP_INV_G11
XG7859 XI11_4/XI0/XI0_21/d_9_ XI11_4/XI0/XI0_21/d__9_ DECAP_INV_G11
XG7860 XI11_4/XI0/XI0_21/d_8_ XI11_4/XI0/XI0_21/d__8_ DECAP_INV_G11
XG7861 XI11_4/XI0/XI0_21/d_7_ XI11_4/XI0/XI0_21/d__7_ DECAP_INV_G11
XG7862 XI11_4/XI0/XI0_21/d_6_ XI11_4/XI0/XI0_21/d__6_ DECAP_INV_G11
XG7863 XI11_4/XI0/XI0_21/d_5_ XI11_4/XI0/XI0_21/d__5_ DECAP_INV_G11
XG7864 XI11_4/XI0/XI0_21/d_4_ XI11_4/XI0/XI0_21/d__4_ DECAP_INV_G11
XG7865 XI11_4/XI0/XI0_21/d_3_ XI11_4/XI0/XI0_21/d__3_ DECAP_INV_G11
XG7866 XI11_4/XI0/XI0_21/d_2_ XI11_4/XI0/XI0_21/d__2_ DECAP_INV_G11
XG7867 XI11_4/XI0/XI0_21/d_1_ XI11_4/XI0/XI0_21/d__1_ DECAP_INV_G11
XG7868 XI11_4/XI0/XI0_21/d_0_ XI11_4/XI0/XI0_21/d__0_ DECAP_INV_G11
XG7869 XI11_4/XI0/XI0_20/d__15_ XI11_4/XI0/XI0_20/d_15_ DECAP_INV_G11
XG7870 XI11_4/XI0/XI0_20/d__14_ XI11_4/XI0/XI0_20/d_14_ DECAP_INV_G11
XG7871 XI11_4/XI0/XI0_20/d__13_ XI11_4/XI0/XI0_20/d_13_ DECAP_INV_G11
XG7872 XI11_4/XI0/XI0_20/d__12_ XI11_4/XI0/XI0_20/d_12_ DECAP_INV_G11
XG7873 XI11_4/XI0/XI0_20/d__11_ XI11_4/XI0/XI0_20/d_11_ DECAP_INV_G11
XG7874 XI11_4/XI0/XI0_20/d__10_ XI11_4/XI0/XI0_20/d_10_ DECAP_INV_G11
XG7875 XI11_4/XI0/XI0_20/d__9_ XI11_4/XI0/XI0_20/d_9_ DECAP_INV_G11
XG7876 XI11_4/XI0/XI0_20/d__8_ XI11_4/XI0/XI0_20/d_8_ DECAP_INV_G11
XG7877 XI11_4/XI0/XI0_20/d__7_ XI11_4/XI0/XI0_20/d_7_ DECAP_INV_G11
XG7878 XI11_4/XI0/XI0_20/d__6_ XI11_4/XI0/XI0_20/d_6_ DECAP_INV_G11
XG7879 XI11_4/XI0/XI0_20/d__5_ XI11_4/XI0/XI0_20/d_5_ DECAP_INV_G11
XG7880 XI11_4/XI0/XI0_20/d__4_ XI11_4/XI0/XI0_20/d_4_ DECAP_INV_G11
XG7881 XI11_4/XI0/XI0_20/d__3_ XI11_4/XI0/XI0_20/d_3_ DECAP_INV_G11
XG7882 XI11_4/XI0/XI0_20/d__2_ XI11_4/XI0/XI0_20/d_2_ DECAP_INV_G11
XG7883 XI11_4/XI0/XI0_20/d__1_ XI11_4/XI0/XI0_20/d_1_ DECAP_INV_G11
XG7884 XI11_4/XI0/XI0_20/d__0_ XI11_4/XI0/XI0_20/d_0_ DECAP_INV_G11
XG7885 XI11_4/XI0/XI0_20/d_15_ XI11_4/XI0/XI0_20/d__15_ DECAP_INV_G11
XG7886 XI11_4/XI0/XI0_20/d_14_ XI11_4/XI0/XI0_20/d__14_ DECAP_INV_G11
XG7887 XI11_4/XI0/XI0_20/d_13_ XI11_4/XI0/XI0_20/d__13_ DECAP_INV_G11
XG7888 XI11_4/XI0/XI0_20/d_12_ XI11_4/XI0/XI0_20/d__12_ DECAP_INV_G11
XG7889 XI11_4/XI0/XI0_20/d_11_ XI11_4/XI0/XI0_20/d__11_ DECAP_INV_G11
XG7890 XI11_4/XI0/XI0_20/d_10_ XI11_4/XI0/XI0_20/d__10_ DECAP_INV_G11
XG7891 XI11_4/XI0/XI0_20/d_9_ XI11_4/XI0/XI0_20/d__9_ DECAP_INV_G11
XG7892 XI11_4/XI0/XI0_20/d_8_ XI11_4/XI0/XI0_20/d__8_ DECAP_INV_G11
XG7893 XI11_4/XI0/XI0_20/d_7_ XI11_4/XI0/XI0_20/d__7_ DECAP_INV_G11
XG7894 XI11_4/XI0/XI0_20/d_6_ XI11_4/XI0/XI0_20/d__6_ DECAP_INV_G11
XG7895 XI11_4/XI0/XI0_20/d_5_ XI11_4/XI0/XI0_20/d__5_ DECAP_INV_G11
XG7896 XI11_4/XI0/XI0_20/d_4_ XI11_4/XI0/XI0_20/d__4_ DECAP_INV_G11
XG7897 XI11_4/XI0/XI0_20/d_3_ XI11_4/XI0/XI0_20/d__3_ DECAP_INV_G11
XG7898 XI11_4/XI0/XI0_20/d_2_ XI11_4/XI0/XI0_20/d__2_ DECAP_INV_G11
XG7899 XI11_4/XI0/XI0_20/d_1_ XI11_4/XI0/XI0_20/d__1_ DECAP_INV_G11
XG7900 XI11_4/XI0/XI0_20/d_0_ XI11_4/XI0/XI0_20/d__0_ DECAP_INV_G11
XG7901 XI11_4/XI0/XI0_19/d__15_ XI11_4/XI0/XI0_19/d_15_ DECAP_INV_G11
XG7902 XI11_4/XI0/XI0_19/d__14_ XI11_4/XI0/XI0_19/d_14_ DECAP_INV_G11
XG7903 XI11_4/XI0/XI0_19/d__13_ XI11_4/XI0/XI0_19/d_13_ DECAP_INV_G11
XG7904 XI11_4/XI0/XI0_19/d__12_ XI11_4/XI0/XI0_19/d_12_ DECAP_INV_G11
XG7905 XI11_4/XI0/XI0_19/d__11_ XI11_4/XI0/XI0_19/d_11_ DECAP_INV_G11
XG7906 XI11_4/XI0/XI0_19/d__10_ XI11_4/XI0/XI0_19/d_10_ DECAP_INV_G11
XG7907 XI11_4/XI0/XI0_19/d__9_ XI11_4/XI0/XI0_19/d_9_ DECAP_INV_G11
XG7908 XI11_4/XI0/XI0_19/d__8_ XI11_4/XI0/XI0_19/d_8_ DECAP_INV_G11
XG7909 XI11_4/XI0/XI0_19/d__7_ XI11_4/XI0/XI0_19/d_7_ DECAP_INV_G11
XG7910 XI11_4/XI0/XI0_19/d__6_ XI11_4/XI0/XI0_19/d_6_ DECAP_INV_G11
XG7911 XI11_4/XI0/XI0_19/d__5_ XI11_4/XI0/XI0_19/d_5_ DECAP_INV_G11
XG7912 XI11_4/XI0/XI0_19/d__4_ XI11_4/XI0/XI0_19/d_4_ DECAP_INV_G11
XG7913 XI11_4/XI0/XI0_19/d__3_ XI11_4/XI0/XI0_19/d_3_ DECAP_INV_G11
XG7914 XI11_4/XI0/XI0_19/d__2_ XI11_4/XI0/XI0_19/d_2_ DECAP_INV_G11
XG7915 XI11_4/XI0/XI0_19/d__1_ XI11_4/XI0/XI0_19/d_1_ DECAP_INV_G11
XG7916 XI11_4/XI0/XI0_19/d__0_ XI11_4/XI0/XI0_19/d_0_ DECAP_INV_G11
XG7917 XI11_4/XI0/XI0_19/d_15_ XI11_4/XI0/XI0_19/d__15_ DECAP_INV_G11
XG7918 XI11_4/XI0/XI0_19/d_14_ XI11_4/XI0/XI0_19/d__14_ DECAP_INV_G11
XG7919 XI11_4/XI0/XI0_19/d_13_ XI11_4/XI0/XI0_19/d__13_ DECAP_INV_G11
XG7920 XI11_4/XI0/XI0_19/d_12_ XI11_4/XI0/XI0_19/d__12_ DECAP_INV_G11
XG7921 XI11_4/XI0/XI0_19/d_11_ XI11_4/XI0/XI0_19/d__11_ DECAP_INV_G11
XG7922 XI11_4/XI0/XI0_19/d_10_ XI11_4/XI0/XI0_19/d__10_ DECAP_INV_G11
XG7923 XI11_4/XI0/XI0_19/d_9_ XI11_4/XI0/XI0_19/d__9_ DECAP_INV_G11
XG7924 XI11_4/XI0/XI0_19/d_8_ XI11_4/XI0/XI0_19/d__8_ DECAP_INV_G11
XG7925 XI11_4/XI0/XI0_19/d_7_ XI11_4/XI0/XI0_19/d__7_ DECAP_INV_G11
XG7926 XI11_4/XI0/XI0_19/d_6_ XI11_4/XI0/XI0_19/d__6_ DECAP_INV_G11
XG7927 XI11_4/XI0/XI0_19/d_5_ XI11_4/XI0/XI0_19/d__5_ DECAP_INV_G11
XG7928 XI11_4/XI0/XI0_19/d_4_ XI11_4/XI0/XI0_19/d__4_ DECAP_INV_G11
XG7929 XI11_4/XI0/XI0_19/d_3_ XI11_4/XI0/XI0_19/d__3_ DECAP_INV_G11
XG7930 XI11_4/XI0/XI0_19/d_2_ XI11_4/XI0/XI0_19/d__2_ DECAP_INV_G11
XG7931 XI11_4/XI0/XI0_19/d_1_ XI11_4/XI0/XI0_19/d__1_ DECAP_INV_G11
XG7932 XI11_4/XI0/XI0_19/d_0_ XI11_4/XI0/XI0_19/d__0_ DECAP_INV_G11
XG7933 XI11_4/XI0/XI0_18/d__15_ XI11_4/XI0/XI0_18/d_15_ DECAP_INV_G11
XG7934 XI11_4/XI0/XI0_18/d__14_ XI11_4/XI0/XI0_18/d_14_ DECAP_INV_G11
XG7935 XI11_4/XI0/XI0_18/d__13_ XI11_4/XI0/XI0_18/d_13_ DECAP_INV_G11
XG7936 XI11_4/XI0/XI0_18/d__12_ XI11_4/XI0/XI0_18/d_12_ DECAP_INV_G11
XG7937 XI11_4/XI0/XI0_18/d__11_ XI11_4/XI0/XI0_18/d_11_ DECAP_INV_G11
XG7938 XI11_4/XI0/XI0_18/d__10_ XI11_4/XI0/XI0_18/d_10_ DECAP_INV_G11
XG7939 XI11_4/XI0/XI0_18/d__9_ XI11_4/XI0/XI0_18/d_9_ DECAP_INV_G11
XG7940 XI11_4/XI0/XI0_18/d__8_ XI11_4/XI0/XI0_18/d_8_ DECAP_INV_G11
XG7941 XI11_4/XI0/XI0_18/d__7_ XI11_4/XI0/XI0_18/d_7_ DECAP_INV_G11
XG7942 XI11_4/XI0/XI0_18/d__6_ XI11_4/XI0/XI0_18/d_6_ DECAP_INV_G11
XG7943 XI11_4/XI0/XI0_18/d__5_ XI11_4/XI0/XI0_18/d_5_ DECAP_INV_G11
XG7944 XI11_4/XI0/XI0_18/d__4_ XI11_4/XI0/XI0_18/d_4_ DECAP_INV_G11
XG7945 XI11_4/XI0/XI0_18/d__3_ XI11_4/XI0/XI0_18/d_3_ DECAP_INV_G11
XG7946 XI11_4/XI0/XI0_18/d__2_ XI11_4/XI0/XI0_18/d_2_ DECAP_INV_G11
XG7947 XI11_4/XI0/XI0_18/d__1_ XI11_4/XI0/XI0_18/d_1_ DECAP_INV_G11
XG7948 XI11_4/XI0/XI0_18/d__0_ XI11_4/XI0/XI0_18/d_0_ DECAP_INV_G11
XG7949 XI11_4/XI0/XI0_18/d_15_ XI11_4/XI0/XI0_18/d__15_ DECAP_INV_G11
XG7950 XI11_4/XI0/XI0_18/d_14_ XI11_4/XI0/XI0_18/d__14_ DECAP_INV_G11
XG7951 XI11_4/XI0/XI0_18/d_13_ XI11_4/XI0/XI0_18/d__13_ DECAP_INV_G11
XG7952 XI11_4/XI0/XI0_18/d_12_ XI11_4/XI0/XI0_18/d__12_ DECAP_INV_G11
XG7953 XI11_4/XI0/XI0_18/d_11_ XI11_4/XI0/XI0_18/d__11_ DECAP_INV_G11
XG7954 XI11_4/XI0/XI0_18/d_10_ XI11_4/XI0/XI0_18/d__10_ DECAP_INV_G11
XG7955 XI11_4/XI0/XI0_18/d_9_ XI11_4/XI0/XI0_18/d__9_ DECAP_INV_G11
XG7956 XI11_4/XI0/XI0_18/d_8_ XI11_4/XI0/XI0_18/d__8_ DECAP_INV_G11
XG7957 XI11_4/XI0/XI0_18/d_7_ XI11_4/XI0/XI0_18/d__7_ DECAP_INV_G11
XG7958 XI11_4/XI0/XI0_18/d_6_ XI11_4/XI0/XI0_18/d__6_ DECAP_INV_G11
XG7959 XI11_4/XI0/XI0_18/d_5_ XI11_4/XI0/XI0_18/d__5_ DECAP_INV_G11
XG7960 XI11_4/XI0/XI0_18/d_4_ XI11_4/XI0/XI0_18/d__4_ DECAP_INV_G11
XG7961 XI11_4/XI0/XI0_18/d_3_ XI11_4/XI0/XI0_18/d__3_ DECAP_INV_G11
XG7962 XI11_4/XI0/XI0_18/d_2_ XI11_4/XI0/XI0_18/d__2_ DECAP_INV_G11
XG7963 XI11_4/XI0/XI0_18/d_1_ XI11_4/XI0/XI0_18/d__1_ DECAP_INV_G11
XG7964 XI11_4/XI0/XI0_18/d_0_ XI11_4/XI0/XI0_18/d__0_ DECAP_INV_G11
XG7965 XI11_4/XI0/XI0_17/d__15_ XI11_4/XI0/XI0_17/d_15_ DECAP_INV_G11
XG7966 XI11_4/XI0/XI0_17/d__14_ XI11_4/XI0/XI0_17/d_14_ DECAP_INV_G11
XG7967 XI11_4/XI0/XI0_17/d__13_ XI11_4/XI0/XI0_17/d_13_ DECAP_INV_G11
XG7968 XI11_4/XI0/XI0_17/d__12_ XI11_4/XI0/XI0_17/d_12_ DECAP_INV_G11
XG7969 XI11_4/XI0/XI0_17/d__11_ XI11_4/XI0/XI0_17/d_11_ DECAP_INV_G11
XG7970 XI11_4/XI0/XI0_17/d__10_ XI11_4/XI0/XI0_17/d_10_ DECAP_INV_G11
XG7971 XI11_4/XI0/XI0_17/d__9_ XI11_4/XI0/XI0_17/d_9_ DECAP_INV_G11
XG7972 XI11_4/XI0/XI0_17/d__8_ XI11_4/XI0/XI0_17/d_8_ DECAP_INV_G11
XG7973 XI11_4/XI0/XI0_17/d__7_ XI11_4/XI0/XI0_17/d_7_ DECAP_INV_G11
XG7974 XI11_4/XI0/XI0_17/d__6_ XI11_4/XI0/XI0_17/d_6_ DECAP_INV_G11
XG7975 XI11_4/XI0/XI0_17/d__5_ XI11_4/XI0/XI0_17/d_5_ DECAP_INV_G11
XG7976 XI11_4/XI0/XI0_17/d__4_ XI11_4/XI0/XI0_17/d_4_ DECAP_INV_G11
XG7977 XI11_4/XI0/XI0_17/d__3_ XI11_4/XI0/XI0_17/d_3_ DECAP_INV_G11
XG7978 XI11_4/XI0/XI0_17/d__2_ XI11_4/XI0/XI0_17/d_2_ DECAP_INV_G11
XG7979 XI11_4/XI0/XI0_17/d__1_ XI11_4/XI0/XI0_17/d_1_ DECAP_INV_G11
XG7980 XI11_4/XI0/XI0_17/d__0_ XI11_4/XI0/XI0_17/d_0_ DECAP_INV_G11
XG7981 XI11_4/XI0/XI0_17/d_15_ XI11_4/XI0/XI0_17/d__15_ DECAP_INV_G11
XG7982 XI11_4/XI0/XI0_17/d_14_ XI11_4/XI0/XI0_17/d__14_ DECAP_INV_G11
XG7983 XI11_4/XI0/XI0_17/d_13_ XI11_4/XI0/XI0_17/d__13_ DECAP_INV_G11
XG7984 XI11_4/XI0/XI0_17/d_12_ XI11_4/XI0/XI0_17/d__12_ DECAP_INV_G11
XG7985 XI11_4/XI0/XI0_17/d_11_ XI11_4/XI0/XI0_17/d__11_ DECAP_INV_G11
XG7986 XI11_4/XI0/XI0_17/d_10_ XI11_4/XI0/XI0_17/d__10_ DECAP_INV_G11
XG7987 XI11_4/XI0/XI0_17/d_9_ XI11_4/XI0/XI0_17/d__9_ DECAP_INV_G11
XG7988 XI11_4/XI0/XI0_17/d_8_ XI11_4/XI0/XI0_17/d__8_ DECAP_INV_G11
XG7989 XI11_4/XI0/XI0_17/d_7_ XI11_4/XI0/XI0_17/d__7_ DECAP_INV_G11
XG7990 XI11_4/XI0/XI0_17/d_6_ XI11_4/XI0/XI0_17/d__6_ DECAP_INV_G11
XG7991 XI11_4/XI0/XI0_17/d_5_ XI11_4/XI0/XI0_17/d__5_ DECAP_INV_G11
XG7992 XI11_4/XI0/XI0_17/d_4_ XI11_4/XI0/XI0_17/d__4_ DECAP_INV_G11
XG7993 XI11_4/XI0/XI0_17/d_3_ XI11_4/XI0/XI0_17/d__3_ DECAP_INV_G11
XG7994 XI11_4/XI0/XI0_17/d_2_ XI11_4/XI0/XI0_17/d__2_ DECAP_INV_G11
XG7995 XI11_4/XI0/XI0_17/d_1_ XI11_4/XI0/XI0_17/d__1_ DECAP_INV_G11
XG7996 XI11_4/XI0/XI0_17/d_0_ XI11_4/XI0/XI0_17/d__0_ DECAP_INV_G11
XG7997 XI11_4/XI0/XI0_16/d__15_ XI11_4/XI0/XI0_16/d_15_ DECAP_INV_G11
XG7998 XI11_4/XI0/XI0_16/d__14_ XI11_4/XI0/XI0_16/d_14_ DECAP_INV_G11
XG7999 XI11_4/XI0/XI0_16/d__13_ XI11_4/XI0/XI0_16/d_13_ DECAP_INV_G11
XG8000 XI11_4/XI0/XI0_16/d__12_ XI11_4/XI0/XI0_16/d_12_ DECAP_INV_G11
XG8001 XI11_4/XI0/XI0_16/d__11_ XI11_4/XI0/XI0_16/d_11_ DECAP_INV_G11
XG8002 XI11_4/XI0/XI0_16/d__10_ XI11_4/XI0/XI0_16/d_10_ DECAP_INV_G11
XG8003 XI11_4/XI0/XI0_16/d__9_ XI11_4/XI0/XI0_16/d_9_ DECAP_INV_G11
XG8004 XI11_4/XI0/XI0_16/d__8_ XI11_4/XI0/XI0_16/d_8_ DECAP_INV_G11
XG8005 XI11_4/XI0/XI0_16/d__7_ XI11_4/XI0/XI0_16/d_7_ DECAP_INV_G11
XG8006 XI11_4/XI0/XI0_16/d__6_ XI11_4/XI0/XI0_16/d_6_ DECAP_INV_G11
XG8007 XI11_4/XI0/XI0_16/d__5_ XI11_4/XI0/XI0_16/d_5_ DECAP_INV_G11
XG8008 XI11_4/XI0/XI0_16/d__4_ XI11_4/XI0/XI0_16/d_4_ DECAP_INV_G11
XG8009 XI11_4/XI0/XI0_16/d__3_ XI11_4/XI0/XI0_16/d_3_ DECAP_INV_G11
XG8010 XI11_4/XI0/XI0_16/d__2_ XI11_4/XI0/XI0_16/d_2_ DECAP_INV_G11
XG8011 XI11_4/XI0/XI0_16/d__1_ XI11_4/XI0/XI0_16/d_1_ DECAP_INV_G11
XG8012 XI11_4/XI0/XI0_16/d__0_ XI11_4/XI0/XI0_16/d_0_ DECAP_INV_G11
XG8013 XI11_4/XI0/XI0_16/d_15_ XI11_4/XI0/XI0_16/d__15_ DECAP_INV_G11
XG8014 XI11_4/XI0/XI0_16/d_14_ XI11_4/XI0/XI0_16/d__14_ DECAP_INV_G11
XG8015 XI11_4/XI0/XI0_16/d_13_ XI11_4/XI0/XI0_16/d__13_ DECAP_INV_G11
XG8016 XI11_4/XI0/XI0_16/d_12_ XI11_4/XI0/XI0_16/d__12_ DECAP_INV_G11
XG8017 XI11_4/XI0/XI0_16/d_11_ XI11_4/XI0/XI0_16/d__11_ DECAP_INV_G11
XG8018 XI11_4/XI0/XI0_16/d_10_ XI11_4/XI0/XI0_16/d__10_ DECAP_INV_G11
XG8019 XI11_4/XI0/XI0_16/d_9_ XI11_4/XI0/XI0_16/d__9_ DECAP_INV_G11
XG8020 XI11_4/XI0/XI0_16/d_8_ XI11_4/XI0/XI0_16/d__8_ DECAP_INV_G11
XG8021 XI11_4/XI0/XI0_16/d_7_ XI11_4/XI0/XI0_16/d__7_ DECAP_INV_G11
XG8022 XI11_4/XI0/XI0_16/d_6_ XI11_4/XI0/XI0_16/d__6_ DECAP_INV_G11
XG8023 XI11_4/XI0/XI0_16/d_5_ XI11_4/XI0/XI0_16/d__5_ DECAP_INV_G11
XG8024 XI11_4/XI0/XI0_16/d_4_ XI11_4/XI0/XI0_16/d__4_ DECAP_INV_G11
XG8025 XI11_4/XI0/XI0_16/d_3_ XI11_4/XI0/XI0_16/d__3_ DECAP_INV_G11
XG8026 XI11_4/XI0/XI0_16/d_2_ XI11_4/XI0/XI0_16/d__2_ DECAP_INV_G11
XG8027 XI11_4/XI0/XI0_16/d_1_ XI11_4/XI0/XI0_16/d__1_ DECAP_INV_G11
XG8028 XI11_4/XI0/XI0_16/d_0_ XI11_4/XI0/XI0_16/d__0_ DECAP_INV_G11
XG8029 XI11_4/XI0/XI0_15/d__15_ XI11_4/XI0/XI0_15/d_15_ DECAP_INV_G11
XG8030 XI11_4/XI0/XI0_15/d__14_ XI11_4/XI0/XI0_15/d_14_ DECAP_INV_G11
XG8031 XI11_4/XI0/XI0_15/d__13_ XI11_4/XI0/XI0_15/d_13_ DECAP_INV_G11
XG8032 XI11_4/XI0/XI0_15/d__12_ XI11_4/XI0/XI0_15/d_12_ DECAP_INV_G11
XG8033 XI11_4/XI0/XI0_15/d__11_ XI11_4/XI0/XI0_15/d_11_ DECAP_INV_G11
XG8034 XI11_4/XI0/XI0_15/d__10_ XI11_4/XI0/XI0_15/d_10_ DECAP_INV_G11
XG8035 XI11_4/XI0/XI0_15/d__9_ XI11_4/XI0/XI0_15/d_9_ DECAP_INV_G11
XG8036 XI11_4/XI0/XI0_15/d__8_ XI11_4/XI0/XI0_15/d_8_ DECAP_INV_G11
XG8037 XI11_4/XI0/XI0_15/d__7_ XI11_4/XI0/XI0_15/d_7_ DECAP_INV_G11
XG8038 XI11_4/XI0/XI0_15/d__6_ XI11_4/XI0/XI0_15/d_6_ DECAP_INV_G11
XG8039 XI11_4/XI0/XI0_15/d__5_ XI11_4/XI0/XI0_15/d_5_ DECAP_INV_G11
XG8040 XI11_4/XI0/XI0_15/d__4_ XI11_4/XI0/XI0_15/d_4_ DECAP_INV_G11
XG8041 XI11_4/XI0/XI0_15/d__3_ XI11_4/XI0/XI0_15/d_3_ DECAP_INV_G11
XG8042 XI11_4/XI0/XI0_15/d__2_ XI11_4/XI0/XI0_15/d_2_ DECAP_INV_G11
XG8043 XI11_4/XI0/XI0_15/d__1_ XI11_4/XI0/XI0_15/d_1_ DECAP_INV_G11
XG8044 XI11_4/XI0/XI0_15/d__0_ XI11_4/XI0/XI0_15/d_0_ DECAP_INV_G11
XG8045 XI11_4/XI0/XI0_15/d_15_ XI11_4/XI0/XI0_15/d__15_ DECAP_INV_G11
XG8046 XI11_4/XI0/XI0_15/d_14_ XI11_4/XI0/XI0_15/d__14_ DECAP_INV_G11
XG8047 XI11_4/XI0/XI0_15/d_13_ XI11_4/XI0/XI0_15/d__13_ DECAP_INV_G11
XG8048 XI11_4/XI0/XI0_15/d_12_ XI11_4/XI0/XI0_15/d__12_ DECAP_INV_G11
XG8049 XI11_4/XI0/XI0_15/d_11_ XI11_4/XI0/XI0_15/d__11_ DECAP_INV_G11
XG8050 XI11_4/XI0/XI0_15/d_10_ XI11_4/XI0/XI0_15/d__10_ DECAP_INV_G11
XG8051 XI11_4/XI0/XI0_15/d_9_ XI11_4/XI0/XI0_15/d__9_ DECAP_INV_G11
XG8052 XI11_4/XI0/XI0_15/d_8_ XI11_4/XI0/XI0_15/d__8_ DECAP_INV_G11
XG8053 XI11_4/XI0/XI0_15/d_7_ XI11_4/XI0/XI0_15/d__7_ DECAP_INV_G11
XG8054 XI11_4/XI0/XI0_15/d_6_ XI11_4/XI0/XI0_15/d__6_ DECAP_INV_G11
XG8055 XI11_4/XI0/XI0_15/d_5_ XI11_4/XI0/XI0_15/d__5_ DECAP_INV_G11
XG8056 XI11_4/XI0/XI0_15/d_4_ XI11_4/XI0/XI0_15/d__4_ DECAP_INV_G11
XG8057 XI11_4/XI0/XI0_15/d_3_ XI11_4/XI0/XI0_15/d__3_ DECAP_INV_G11
XG8058 XI11_4/XI0/XI0_15/d_2_ XI11_4/XI0/XI0_15/d__2_ DECAP_INV_G11
XG8059 XI11_4/XI0/XI0_15/d_1_ XI11_4/XI0/XI0_15/d__1_ DECAP_INV_G11
XG8060 XI11_4/XI0/XI0_15/d_0_ XI11_4/XI0/XI0_15/d__0_ DECAP_INV_G11
XG8061 XI11_4/XI0/XI0_14/d__15_ XI11_4/XI0/XI0_14/d_15_ DECAP_INV_G11
XG8062 XI11_4/XI0/XI0_14/d__14_ XI11_4/XI0/XI0_14/d_14_ DECAP_INV_G11
XG8063 XI11_4/XI0/XI0_14/d__13_ XI11_4/XI0/XI0_14/d_13_ DECAP_INV_G11
XG8064 XI11_4/XI0/XI0_14/d__12_ XI11_4/XI0/XI0_14/d_12_ DECAP_INV_G11
XG8065 XI11_4/XI0/XI0_14/d__11_ XI11_4/XI0/XI0_14/d_11_ DECAP_INV_G11
XG8066 XI11_4/XI0/XI0_14/d__10_ XI11_4/XI0/XI0_14/d_10_ DECAP_INV_G11
XG8067 XI11_4/XI0/XI0_14/d__9_ XI11_4/XI0/XI0_14/d_9_ DECAP_INV_G11
XG8068 XI11_4/XI0/XI0_14/d__8_ XI11_4/XI0/XI0_14/d_8_ DECAP_INV_G11
XG8069 XI11_4/XI0/XI0_14/d__7_ XI11_4/XI0/XI0_14/d_7_ DECAP_INV_G11
XG8070 XI11_4/XI0/XI0_14/d__6_ XI11_4/XI0/XI0_14/d_6_ DECAP_INV_G11
XG8071 XI11_4/XI0/XI0_14/d__5_ XI11_4/XI0/XI0_14/d_5_ DECAP_INV_G11
XG8072 XI11_4/XI0/XI0_14/d__4_ XI11_4/XI0/XI0_14/d_4_ DECAP_INV_G11
XG8073 XI11_4/XI0/XI0_14/d__3_ XI11_4/XI0/XI0_14/d_3_ DECAP_INV_G11
XG8074 XI11_4/XI0/XI0_14/d__2_ XI11_4/XI0/XI0_14/d_2_ DECAP_INV_G11
XG8075 XI11_4/XI0/XI0_14/d__1_ XI11_4/XI0/XI0_14/d_1_ DECAP_INV_G11
XG8076 XI11_4/XI0/XI0_14/d__0_ XI11_4/XI0/XI0_14/d_0_ DECAP_INV_G11
XG8077 XI11_4/XI0/XI0_14/d_15_ XI11_4/XI0/XI0_14/d__15_ DECAP_INV_G11
XG8078 XI11_4/XI0/XI0_14/d_14_ XI11_4/XI0/XI0_14/d__14_ DECAP_INV_G11
XG8079 XI11_4/XI0/XI0_14/d_13_ XI11_4/XI0/XI0_14/d__13_ DECAP_INV_G11
XG8080 XI11_4/XI0/XI0_14/d_12_ XI11_4/XI0/XI0_14/d__12_ DECAP_INV_G11
XG8081 XI11_4/XI0/XI0_14/d_11_ XI11_4/XI0/XI0_14/d__11_ DECAP_INV_G11
XG8082 XI11_4/XI0/XI0_14/d_10_ XI11_4/XI0/XI0_14/d__10_ DECAP_INV_G11
XG8083 XI11_4/XI0/XI0_14/d_9_ XI11_4/XI0/XI0_14/d__9_ DECAP_INV_G11
XG8084 XI11_4/XI0/XI0_14/d_8_ XI11_4/XI0/XI0_14/d__8_ DECAP_INV_G11
XG8085 XI11_4/XI0/XI0_14/d_7_ XI11_4/XI0/XI0_14/d__7_ DECAP_INV_G11
XG8086 XI11_4/XI0/XI0_14/d_6_ XI11_4/XI0/XI0_14/d__6_ DECAP_INV_G11
XG8087 XI11_4/XI0/XI0_14/d_5_ XI11_4/XI0/XI0_14/d__5_ DECAP_INV_G11
XG8088 XI11_4/XI0/XI0_14/d_4_ XI11_4/XI0/XI0_14/d__4_ DECAP_INV_G11
XG8089 XI11_4/XI0/XI0_14/d_3_ XI11_4/XI0/XI0_14/d__3_ DECAP_INV_G11
XG8090 XI11_4/XI0/XI0_14/d_2_ XI11_4/XI0/XI0_14/d__2_ DECAP_INV_G11
XG8091 XI11_4/XI0/XI0_14/d_1_ XI11_4/XI0/XI0_14/d__1_ DECAP_INV_G11
XG8092 XI11_4/XI0/XI0_14/d_0_ XI11_4/XI0/XI0_14/d__0_ DECAP_INV_G11
XG8093 XI11_4/XI0/XI0_13/d__15_ XI11_4/XI0/XI0_13/d_15_ DECAP_INV_G11
XG8094 XI11_4/XI0/XI0_13/d__14_ XI11_4/XI0/XI0_13/d_14_ DECAP_INV_G11
XG8095 XI11_4/XI0/XI0_13/d__13_ XI11_4/XI0/XI0_13/d_13_ DECAP_INV_G11
XG8096 XI11_4/XI0/XI0_13/d__12_ XI11_4/XI0/XI0_13/d_12_ DECAP_INV_G11
XG8097 XI11_4/XI0/XI0_13/d__11_ XI11_4/XI0/XI0_13/d_11_ DECAP_INV_G11
XG8098 XI11_4/XI0/XI0_13/d__10_ XI11_4/XI0/XI0_13/d_10_ DECAP_INV_G11
XG8099 XI11_4/XI0/XI0_13/d__9_ XI11_4/XI0/XI0_13/d_9_ DECAP_INV_G11
XG8100 XI11_4/XI0/XI0_13/d__8_ XI11_4/XI0/XI0_13/d_8_ DECAP_INV_G11
XG8101 XI11_4/XI0/XI0_13/d__7_ XI11_4/XI0/XI0_13/d_7_ DECAP_INV_G11
XG8102 XI11_4/XI0/XI0_13/d__6_ XI11_4/XI0/XI0_13/d_6_ DECAP_INV_G11
XG8103 XI11_4/XI0/XI0_13/d__5_ XI11_4/XI0/XI0_13/d_5_ DECAP_INV_G11
XG8104 XI11_4/XI0/XI0_13/d__4_ XI11_4/XI0/XI0_13/d_4_ DECAP_INV_G11
XG8105 XI11_4/XI0/XI0_13/d__3_ XI11_4/XI0/XI0_13/d_3_ DECAP_INV_G11
XG8106 XI11_4/XI0/XI0_13/d__2_ XI11_4/XI0/XI0_13/d_2_ DECAP_INV_G11
XG8107 XI11_4/XI0/XI0_13/d__1_ XI11_4/XI0/XI0_13/d_1_ DECAP_INV_G11
XG8108 XI11_4/XI0/XI0_13/d__0_ XI11_4/XI0/XI0_13/d_0_ DECAP_INV_G11
XG8109 XI11_4/XI0/XI0_13/d_15_ XI11_4/XI0/XI0_13/d__15_ DECAP_INV_G11
XG8110 XI11_4/XI0/XI0_13/d_14_ XI11_4/XI0/XI0_13/d__14_ DECAP_INV_G11
XG8111 XI11_4/XI0/XI0_13/d_13_ XI11_4/XI0/XI0_13/d__13_ DECAP_INV_G11
XG8112 XI11_4/XI0/XI0_13/d_12_ XI11_4/XI0/XI0_13/d__12_ DECAP_INV_G11
XG8113 XI11_4/XI0/XI0_13/d_11_ XI11_4/XI0/XI0_13/d__11_ DECAP_INV_G11
XG8114 XI11_4/XI0/XI0_13/d_10_ XI11_4/XI0/XI0_13/d__10_ DECAP_INV_G11
XG8115 XI11_4/XI0/XI0_13/d_9_ XI11_4/XI0/XI0_13/d__9_ DECAP_INV_G11
XG8116 XI11_4/XI0/XI0_13/d_8_ XI11_4/XI0/XI0_13/d__8_ DECAP_INV_G11
XG8117 XI11_4/XI0/XI0_13/d_7_ XI11_4/XI0/XI0_13/d__7_ DECAP_INV_G11
XG8118 XI11_4/XI0/XI0_13/d_6_ XI11_4/XI0/XI0_13/d__6_ DECAP_INV_G11
XG8119 XI11_4/XI0/XI0_13/d_5_ XI11_4/XI0/XI0_13/d__5_ DECAP_INV_G11
XG8120 XI11_4/XI0/XI0_13/d_4_ XI11_4/XI0/XI0_13/d__4_ DECAP_INV_G11
XG8121 XI11_4/XI0/XI0_13/d_3_ XI11_4/XI0/XI0_13/d__3_ DECAP_INV_G11
XG8122 XI11_4/XI0/XI0_13/d_2_ XI11_4/XI0/XI0_13/d__2_ DECAP_INV_G11
XG8123 XI11_4/XI0/XI0_13/d_1_ XI11_4/XI0/XI0_13/d__1_ DECAP_INV_G11
XG8124 XI11_4/XI0/XI0_13/d_0_ XI11_4/XI0/XI0_13/d__0_ DECAP_INV_G11
XG8125 XI11_4/XI0/XI0_12/d__15_ XI11_4/XI0/XI0_12/d_15_ DECAP_INV_G11
XG8126 XI11_4/XI0/XI0_12/d__14_ XI11_4/XI0/XI0_12/d_14_ DECAP_INV_G11
XG8127 XI11_4/XI0/XI0_12/d__13_ XI11_4/XI0/XI0_12/d_13_ DECAP_INV_G11
XG8128 XI11_4/XI0/XI0_12/d__12_ XI11_4/XI0/XI0_12/d_12_ DECAP_INV_G11
XG8129 XI11_4/XI0/XI0_12/d__11_ XI11_4/XI0/XI0_12/d_11_ DECAP_INV_G11
XG8130 XI11_4/XI0/XI0_12/d__10_ XI11_4/XI0/XI0_12/d_10_ DECAP_INV_G11
XG8131 XI11_4/XI0/XI0_12/d__9_ XI11_4/XI0/XI0_12/d_9_ DECAP_INV_G11
XG8132 XI11_4/XI0/XI0_12/d__8_ XI11_4/XI0/XI0_12/d_8_ DECAP_INV_G11
XG8133 XI11_4/XI0/XI0_12/d__7_ XI11_4/XI0/XI0_12/d_7_ DECAP_INV_G11
XG8134 XI11_4/XI0/XI0_12/d__6_ XI11_4/XI0/XI0_12/d_6_ DECAP_INV_G11
XG8135 XI11_4/XI0/XI0_12/d__5_ XI11_4/XI0/XI0_12/d_5_ DECAP_INV_G11
XG8136 XI11_4/XI0/XI0_12/d__4_ XI11_4/XI0/XI0_12/d_4_ DECAP_INV_G11
XG8137 XI11_4/XI0/XI0_12/d__3_ XI11_4/XI0/XI0_12/d_3_ DECAP_INV_G11
XG8138 XI11_4/XI0/XI0_12/d__2_ XI11_4/XI0/XI0_12/d_2_ DECAP_INV_G11
XG8139 XI11_4/XI0/XI0_12/d__1_ XI11_4/XI0/XI0_12/d_1_ DECAP_INV_G11
XG8140 XI11_4/XI0/XI0_12/d__0_ XI11_4/XI0/XI0_12/d_0_ DECAP_INV_G11
XG8141 XI11_4/XI0/XI0_12/d_15_ XI11_4/XI0/XI0_12/d__15_ DECAP_INV_G11
XG8142 XI11_4/XI0/XI0_12/d_14_ XI11_4/XI0/XI0_12/d__14_ DECAP_INV_G11
XG8143 XI11_4/XI0/XI0_12/d_13_ XI11_4/XI0/XI0_12/d__13_ DECAP_INV_G11
XG8144 XI11_4/XI0/XI0_12/d_12_ XI11_4/XI0/XI0_12/d__12_ DECAP_INV_G11
XG8145 XI11_4/XI0/XI0_12/d_11_ XI11_4/XI0/XI0_12/d__11_ DECAP_INV_G11
XG8146 XI11_4/XI0/XI0_12/d_10_ XI11_4/XI0/XI0_12/d__10_ DECAP_INV_G11
XG8147 XI11_4/XI0/XI0_12/d_9_ XI11_4/XI0/XI0_12/d__9_ DECAP_INV_G11
XG8148 XI11_4/XI0/XI0_12/d_8_ XI11_4/XI0/XI0_12/d__8_ DECAP_INV_G11
XG8149 XI11_4/XI0/XI0_12/d_7_ XI11_4/XI0/XI0_12/d__7_ DECAP_INV_G11
XG8150 XI11_4/XI0/XI0_12/d_6_ XI11_4/XI0/XI0_12/d__6_ DECAP_INV_G11
XG8151 XI11_4/XI0/XI0_12/d_5_ XI11_4/XI0/XI0_12/d__5_ DECAP_INV_G11
XG8152 XI11_4/XI0/XI0_12/d_4_ XI11_4/XI0/XI0_12/d__4_ DECAP_INV_G11
XG8153 XI11_4/XI0/XI0_12/d_3_ XI11_4/XI0/XI0_12/d__3_ DECAP_INV_G11
XG8154 XI11_4/XI0/XI0_12/d_2_ XI11_4/XI0/XI0_12/d__2_ DECAP_INV_G11
XG8155 XI11_4/XI0/XI0_12/d_1_ XI11_4/XI0/XI0_12/d__1_ DECAP_INV_G11
XG8156 XI11_4/XI0/XI0_12/d_0_ XI11_4/XI0/XI0_12/d__0_ DECAP_INV_G11
XG8157 XI11_4/XI0/XI0_11/d__15_ XI11_4/XI0/XI0_11/d_15_ DECAP_INV_G11
XG8158 XI11_4/XI0/XI0_11/d__14_ XI11_4/XI0/XI0_11/d_14_ DECAP_INV_G11
XG8159 XI11_4/XI0/XI0_11/d__13_ XI11_4/XI0/XI0_11/d_13_ DECAP_INV_G11
XG8160 XI11_4/XI0/XI0_11/d__12_ XI11_4/XI0/XI0_11/d_12_ DECAP_INV_G11
XG8161 XI11_4/XI0/XI0_11/d__11_ XI11_4/XI0/XI0_11/d_11_ DECAP_INV_G11
XG8162 XI11_4/XI0/XI0_11/d__10_ XI11_4/XI0/XI0_11/d_10_ DECAP_INV_G11
XG8163 XI11_4/XI0/XI0_11/d__9_ XI11_4/XI0/XI0_11/d_9_ DECAP_INV_G11
XG8164 XI11_4/XI0/XI0_11/d__8_ XI11_4/XI0/XI0_11/d_8_ DECAP_INV_G11
XG8165 XI11_4/XI0/XI0_11/d__7_ XI11_4/XI0/XI0_11/d_7_ DECAP_INV_G11
XG8166 XI11_4/XI0/XI0_11/d__6_ XI11_4/XI0/XI0_11/d_6_ DECAP_INV_G11
XG8167 XI11_4/XI0/XI0_11/d__5_ XI11_4/XI0/XI0_11/d_5_ DECAP_INV_G11
XG8168 XI11_4/XI0/XI0_11/d__4_ XI11_4/XI0/XI0_11/d_4_ DECAP_INV_G11
XG8169 XI11_4/XI0/XI0_11/d__3_ XI11_4/XI0/XI0_11/d_3_ DECAP_INV_G11
XG8170 XI11_4/XI0/XI0_11/d__2_ XI11_4/XI0/XI0_11/d_2_ DECAP_INV_G11
XG8171 XI11_4/XI0/XI0_11/d__1_ XI11_4/XI0/XI0_11/d_1_ DECAP_INV_G11
XG8172 XI11_4/XI0/XI0_11/d__0_ XI11_4/XI0/XI0_11/d_0_ DECAP_INV_G11
XG8173 XI11_4/XI0/XI0_11/d_15_ XI11_4/XI0/XI0_11/d__15_ DECAP_INV_G11
XG8174 XI11_4/XI0/XI0_11/d_14_ XI11_4/XI0/XI0_11/d__14_ DECAP_INV_G11
XG8175 XI11_4/XI0/XI0_11/d_13_ XI11_4/XI0/XI0_11/d__13_ DECAP_INV_G11
XG8176 XI11_4/XI0/XI0_11/d_12_ XI11_4/XI0/XI0_11/d__12_ DECAP_INV_G11
XG8177 XI11_4/XI0/XI0_11/d_11_ XI11_4/XI0/XI0_11/d__11_ DECAP_INV_G11
XG8178 XI11_4/XI0/XI0_11/d_10_ XI11_4/XI0/XI0_11/d__10_ DECAP_INV_G11
XG8179 XI11_4/XI0/XI0_11/d_9_ XI11_4/XI0/XI0_11/d__9_ DECAP_INV_G11
XG8180 XI11_4/XI0/XI0_11/d_8_ XI11_4/XI0/XI0_11/d__8_ DECAP_INV_G11
XG8181 XI11_4/XI0/XI0_11/d_7_ XI11_4/XI0/XI0_11/d__7_ DECAP_INV_G11
XG8182 XI11_4/XI0/XI0_11/d_6_ XI11_4/XI0/XI0_11/d__6_ DECAP_INV_G11
XG8183 XI11_4/XI0/XI0_11/d_5_ XI11_4/XI0/XI0_11/d__5_ DECAP_INV_G11
XG8184 XI11_4/XI0/XI0_11/d_4_ XI11_4/XI0/XI0_11/d__4_ DECAP_INV_G11
XG8185 XI11_4/XI0/XI0_11/d_3_ XI11_4/XI0/XI0_11/d__3_ DECAP_INV_G11
XG8186 XI11_4/XI0/XI0_11/d_2_ XI11_4/XI0/XI0_11/d__2_ DECAP_INV_G11
XG8187 XI11_4/XI0/XI0_11/d_1_ XI11_4/XI0/XI0_11/d__1_ DECAP_INV_G11
XG8188 XI11_4/XI0/XI0_11/d_0_ XI11_4/XI0/XI0_11/d__0_ DECAP_INV_G11
XG8189 XI11_4/XI0/XI0_10/d__15_ XI11_4/XI0/XI0_10/d_15_ DECAP_INV_G11
XG8190 XI11_4/XI0/XI0_10/d__14_ XI11_4/XI0/XI0_10/d_14_ DECAP_INV_G11
XG8191 XI11_4/XI0/XI0_10/d__13_ XI11_4/XI0/XI0_10/d_13_ DECAP_INV_G11
XG8192 XI11_4/XI0/XI0_10/d__12_ XI11_4/XI0/XI0_10/d_12_ DECAP_INV_G11
XG8193 XI11_4/XI0/XI0_10/d__11_ XI11_4/XI0/XI0_10/d_11_ DECAP_INV_G11
XG8194 XI11_4/XI0/XI0_10/d__10_ XI11_4/XI0/XI0_10/d_10_ DECAP_INV_G11
XG8195 XI11_4/XI0/XI0_10/d__9_ XI11_4/XI0/XI0_10/d_9_ DECAP_INV_G11
XG8196 XI11_4/XI0/XI0_10/d__8_ XI11_4/XI0/XI0_10/d_8_ DECAP_INV_G11
XG8197 XI11_4/XI0/XI0_10/d__7_ XI11_4/XI0/XI0_10/d_7_ DECAP_INV_G11
XG8198 XI11_4/XI0/XI0_10/d__6_ XI11_4/XI0/XI0_10/d_6_ DECAP_INV_G11
XG8199 XI11_4/XI0/XI0_10/d__5_ XI11_4/XI0/XI0_10/d_5_ DECAP_INV_G11
XG8200 XI11_4/XI0/XI0_10/d__4_ XI11_4/XI0/XI0_10/d_4_ DECAP_INV_G11
XG8201 XI11_4/XI0/XI0_10/d__3_ XI11_4/XI0/XI0_10/d_3_ DECAP_INV_G11
XG8202 XI11_4/XI0/XI0_10/d__2_ XI11_4/XI0/XI0_10/d_2_ DECAP_INV_G11
XG8203 XI11_4/XI0/XI0_10/d__1_ XI11_4/XI0/XI0_10/d_1_ DECAP_INV_G11
XG8204 XI11_4/XI0/XI0_10/d__0_ XI11_4/XI0/XI0_10/d_0_ DECAP_INV_G11
XG8205 XI11_4/XI0/XI0_10/d_15_ XI11_4/XI0/XI0_10/d__15_ DECAP_INV_G11
XG8206 XI11_4/XI0/XI0_10/d_14_ XI11_4/XI0/XI0_10/d__14_ DECAP_INV_G11
XG8207 XI11_4/XI0/XI0_10/d_13_ XI11_4/XI0/XI0_10/d__13_ DECAP_INV_G11
XG8208 XI11_4/XI0/XI0_10/d_12_ XI11_4/XI0/XI0_10/d__12_ DECAP_INV_G11
XG8209 XI11_4/XI0/XI0_10/d_11_ XI11_4/XI0/XI0_10/d__11_ DECAP_INV_G11
XG8210 XI11_4/XI0/XI0_10/d_10_ XI11_4/XI0/XI0_10/d__10_ DECAP_INV_G11
XG8211 XI11_4/XI0/XI0_10/d_9_ XI11_4/XI0/XI0_10/d__9_ DECAP_INV_G11
XG8212 XI11_4/XI0/XI0_10/d_8_ XI11_4/XI0/XI0_10/d__8_ DECAP_INV_G11
XG8213 XI11_4/XI0/XI0_10/d_7_ XI11_4/XI0/XI0_10/d__7_ DECAP_INV_G11
XG8214 XI11_4/XI0/XI0_10/d_6_ XI11_4/XI0/XI0_10/d__6_ DECAP_INV_G11
XG8215 XI11_4/XI0/XI0_10/d_5_ XI11_4/XI0/XI0_10/d__5_ DECAP_INV_G11
XG8216 XI11_4/XI0/XI0_10/d_4_ XI11_4/XI0/XI0_10/d__4_ DECAP_INV_G11
XG8217 XI11_4/XI0/XI0_10/d_3_ XI11_4/XI0/XI0_10/d__3_ DECAP_INV_G11
XG8218 XI11_4/XI0/XI0_10/d_2_ XI11_4/XI0/XI0_10/d__2_ DECAP_INV_G11
XG8219 XI11_4/XI0/XI0_10/d_1_ XI11_4/XI0/XI0_10/d__1_ DECAP_INV_G11
XG8220 XI11_4/XI0/XI0_10/d_0_ XI11_4/XI0/XI0_10/d__0_ DECAP_INV_G11
XG8221 XI11_4/XI0/XI0_9/d__15_ XI11_4/XI0/XI0_9/d_15_ DECAP_INV_G11
XG8222 XI11_4/XI0/XI0_9/d__14_ XI11_4/XI0/XI0_9/d_14_ DECAP_INV_G11
XG8223 XI11_4/XI0/XI0_9/d__13_ XI11_4/XI0/XI0_9/d_13_ DECAP_INV_G11
XG8224 XI11_4/XI0/XI0_9/d__12_ XI11_4/XI0/XI0_9/d_12_ DECAP_INV_G11
XG8225 XI11_4/XI0/XI0_9/d__11_ XI11_4/XI0/XI0_9/d_11_ DECAP_INV_G11
XG8226 XI11_4/XI0/XI0_9/d__10_ XI11_4/XI0/XI0_9/d_10_ DECAP_INV_G11
XG8227 XI11_4/XI0/XI0_9/d__9_ XI11_4/XI0/XI0_9/d_9_ DECAP_INV_G11
XG8228 XI11_4/XI0/XI0_9/d__8_ XI11_4/XI0/XI0_9/d_8_ DECAP_INV_G11
XG8229 XI11_4/XI0/XI0_9/d__7_ XI11_4/XI0/XI0_9/d_7_ DECAP_INV_G11
XG8230 XI11_4/XI0/XI0_9/d__6_ XI11_4/XI0/XI0_9/d_6_ DECAP_INV_G11
XG8231 XI11_4/XI0/XI0_9/d__5_ XI11_4/XI0/XI0_9/d_5_ DECAP_INV_G11
XG8232 XI11_4/XI0/XI0_9/d__4_ XI11_4/XI0/XI0_9/d_4_ DECAP_INV_G11
XG8233 XI11_4/XI0/XI0_9/d__3_ XI11_4/XI0/XI0_9/d_3_ DECAP_INV_G11
XG8234 XI11_4/XI0/XI0_9/d__2_ XI11_4/XI0/XI0_9/d_2_ DECAP_INV_G11
XG8235 XI11_4/XI0/XI0_9/d__1_ XI11_4/XI0/XI0_9/d_1_ DECAP_INV_G11
XG8236 XI11_4/XI0/XI0_9/d__0_ XI11_4/XI0/XI0_9/d_0_ DECAP_INV_G11
XG8237 XI11_4/XI0/XI0_9/d_15_ XI11_4/XI0/XI0_9/d__15_ DECAP_INV_G11
XG8238 XI11_4/XI0/XI0_9/d_14_ XI11_4/XI0/XI0_9/d__14_ DECAP_INV_G11
XG8239 XI11_4/XI0/XI0_9/d_13_ XI11_4/XI0/XI0_9/d__13_ DECAP_INV_G11
XG8240 XI11_4/XI0/XI0_9/d_12_ XI11_4/XI0/XI0_9/d__12_ DECAP_INV_G11
XG8241 XI11_4/XI0/XI0_9/d_11_ XI11_4/XI0/XI0_9/d__11_ DECAP_INV_G11
XG8242 XI11_4/XI0/XI0_9/d_10_ XI11_4/XI0/XI0_9/d__10_ DECAP_INV_G11
XG8243 XI11_4/XI0/XI0_9/d_9_ XI11_4/XI0/XI0_9/d__9_ DECAP_INV_G11
XG8244 XI11_4/XI0/XI0_9/d_8_ XI11_4/XI0/XI0_9/d__8_ DECAP_INV_G11
XG8245 XI11_4/XI0/XI0_9/d_7_ XI11_4/XI0/XI0_9/d__7_ DECAP_INV_G11
XG8246 XI11_4/XI0/XI0_9/d_6_ XI11_4/XI0/XI0_9/d__6_ DECAP_INV_G11
XG8247 XI11_4/XI0/XI0_9/d_5_ XI11_4/XI0/XI0_9/d__5_ DECAP_INV_G11
XG8248 XI11_4/XI0/XI0_9/d_4_ XI11_4/XI0/XI0_9/d__4_ DECAP_INV_G11
XG8249 XI11_4/XI0/XI0_9/d_3_ XI11_4/XI0/XI0_9/d__3_ DECAP_INV_G11
XG8250 XI11_4/XI0/XI0_9/d_2_ XI11_4/XI0/XI0_9/d__2_ DECAP_INV_G11
XG8251 XI11_4/XI0/XI0_9/d_1_ XI11_4/XI0/XI0_9/d__1_ DECAP_INV_G11
XG8252 XI11_4/XI0/XI0_9/d_0_ XI11_4/XI0/XI0_9/d__0_ DECAP_INV_G11
XG8253 XI11_4/XI0/XI0_8/d__15_ XI11_4/XI0/XI0_8/d_15_ DECAP_INV_G11
XG8254 XI11_4/XI0/XI0_8/d__14_ XI11_4/XI0/XI0_8/d_14_ DECAP_INV_G11
XG8255 XI11_4/XI0/XI0_8/d__13_ XI11_4/XI0/XI0_8/d_13_ DECAP_INV_G11
XG8256 XI11_4/XI0/XI0_8/d__12_ XI11_4/XI0/XI0_8/d_12_ DECAP_INV_G11
XG8257 XI11_4/XI0/XI0_8/d__11_ XI11_4/XI0/XI0_8/d_11_ DECAP_INV_G11
XG8258 XI11_4/XI0/XI0_8/d__10_ XI11_4/XI0/XI0_8/d_10_ DECAP_INV_G11
XG8259 XI11_4/XI0/XI0_8/d__9_ XI11_4/XI0/XI0_8/d_9_ DECAP_INV_G11
XG8260 XI11_4/XI0/XI0_8/d__8_ XI11_4/XI0/XI0_8/d_8_ DECAP_INV_G11
XG8261 XI11_4/XI0/XI0_8/d__7_ XI11_4/XI0/XI0_8/d_7_ DECAP_INV_G11
XG8262 XI11_4/XI0/XI0_8/d__6_ XI11_4/XI0/XI0_8/d_6_ DECAP_INV_G11
XG8263 XI11_4/XI0/XI0_8/d__5_ XI11_4/XI0/XI0_8/d_5_ DECAP_INV_G11
XG8264 XI11_4/XI0/XI0_8/d__4_ XI11_4/XI0/XI0_8/d_4_ DECAP_INV_G11
XG8265 XI11_4/XI0/XI0_8/d__3_ XI11_4/XI0/XI0_8/d_3_ DECAP_INV_G11
XG8266 XI11_4/XI0/XI0_8/d__2_ XI11_4/XI0/XI0_8/d_2_ DECAP_INV_G11
XG8267 XI11_4/XI0/XI0_8/d__1_ XI11_4/XI0/XI0_8/d_1_ DECAP_INV_G11
XG8268 XI11_4/XI0/XI0_8/d__0_ XI11_4/XI0/XI0_8/d_0_ DECAP_INV_G11
XG8269 XI11_4/XI0/XI0_8/d_15_ XI11_4/XI0/XI0_8/d__15_ DECAP_INV_G11
XG8270 XI11_4/XI0/XI0_8/d_14_ XI11_4/XI0/XI0_8/d__14_ DECAP_INV_G11
XG8271 XI11_4/XI0/XI0_8/d_13_ XI11_4/XI0/XI0_8/d__13_ DECAP_INV_G11
XG8272 XI11_4/XI0/XI0_8/d_12_ XI11_4/XI0/XI0_8/d__12_ DECAP_INV_G11
XG8273 XI11_4/XI0/XI0_8/d_11_ XI11_4/XI0/XI0_8/d__11_ DECAP_INV_G11
XG8274 XI11_4/XI0/XI0_8/d_10_ XI11_4/XI0/XI0_8/d__10_ DECAP_INV_G11
XG8275 XI11_4/XI0/XI0_8/d_9_ XI11_4/XI0/XI0_8/d__9_ DECAP_INV_G11
XG8276 XI11_4/XI0/XI0_8/d_8_ XI11_4/XI0/XI0_8/d__8_ DECAP_INV_G11
XG8277 XI11_4/XI0/XI0_8/d_7_ XI11_4/XI0/XI0_8/d__7_ DECAP_INV_G11
XG8278 XI11_4/XI0/XI0_8/d_6_ XI11_4/XI0/XI0_8/d__6_ DECAP_INV_G11
XG8279 XI11_4/XI0/XI0_8/d_5_ XI11_4/XI0/XI0_8/d__5_ DECAP_INV_G11
XG8280 XI11_4/XI0/XI0_8/d_4_ XI11_4/XI0/XI0_8/d__4_ DECAP_INV_G11
XG8281 XI11_4/XI0/XI0_8/d_3_ XI11_4/XI0/XI0_8/d__3_ DECAP_INV_G11
XG8282 XI11_4/XI0/XI0_8/d_2_ XI11_4/XI0/XI0_8/d__2_ DECAP_INV_G11
XG8283 XI11_4/XI0/XI0_8/d_1_ XI11_4/XI0/XI0_8/d__1_ DECAP_INV_G11
XG8284 XI11_4/XI0/XI0_8/d_0_ XI11_4/XI0/XI0_8/d__0_ DECAP_INV_G11
XG8285 XI11_4/XI0/XI0_7/d__15_ XI11_4/XI0/XI0_7/d_15_ DECAP_INV_G11
XG8286 XI11_4/XI0/XI0_7/d__14_ XI11_4/XI0/XI0_7/d_14_ DECAP_INV_G11
XG8287 XI11_4/XI0/XI0_7/d__13_ XI11_4/XI0/XI0_7/d_13_ DECAP_INV_G11
XG8288 XI11_4/XI0/XI0_7/d__12_ XI11_4/XI0/XI0_7/d_12_ DECAP_INV_G11
XG8289 XI11_4/XI0/XI0_7/d__11_ XI11_4/XI0/XI0_7/d_11_ DECAP_INV_G11
XG8290 XI11_4/XI0/XI0_7/d__10_ XI11_4/XI0/XI0_7/d_10_ DECAP_INV_G11
XG8291 XI11_4/XI0/XI0_7/d__9_ XI11_4/XI0/XI0_7/d_9_ DECAP_INV_G11
XG8292 XI11_4/XI0/XI0_7/d__8_ XI11_4/XI0/XI0_7/d_8_ DECAP_INV_G11
XG8293 XI11_4/XI0/XI0_7/d__7_ XI11_4/XI0/XI0_7/d_7_ DECAP_INV_G11
XG8294 XI11_4/XI0/XI0_7/d__6_ XI11_4/XI0/XI0_7/d_6_ DECAP_INV_G11
XG8295 XI11_4/XI0/XI0_7/d__5_ XI11_4/XI0/XI0_7/d_5_ DECAP_INV_G11
XG8296 XI11_4/XI0/XI0_7/d__4_ XI11_4/XI0/XI0_7/d_4_ DECAP_INV_G11
XG8297 XI11_4/XI0/XI0_7/d__3_ XI11_4/XI0/XI0_7/d_3_ DECAP_INV_G11
XG8298 XI11_4/XI0/XI0_7/d__2_ XI11_4/XI0/XI0_7/d_2_ DECAP_INV_G11
XG8299 XI11_4/XI0/XI0_7/d__1_ XI11_4/XI0/XI0_7/d_1_ DECAP_INV_G11
XG8300 XI11_4/XI0/XI0_7/d__0_ XI11_4/XI0/XI0_7/d_0_ DECAP_INV_G11
XG8301 XI11_4/XI0/XI0_7/d_15_ XI11_4/XI0/XI0_7/d__15_ DECAP_INV_G11
XG8302 XI11_4/XI0/XI0_7/d_14_ XI11_4/XI0/XI0_7/d__14_ DECAP_INV_G11
XG8303 XI11_4/XI0/XI0_7/d_13_ XI11_4/XI0/XI0_7/d__13_ DECAP_INV_G11
XG8304 XI11_4/XI0/XI0_7/d_12_ XI11_4/XI0/XI0_7/d__12_ DECAP_INV_G11
XG8305 XI11_4/XI0/XI0_7/d_11_ XI11_4/XI0/XI0_7/d__11_ DECAP_INV_G11
XG8306 XI11_4/XI0/XI0_7/d_10_ XI11_4/XI0/XI0_7/d__10_ DECAP_INV_G11
XG8307 XI11_4/XI0/XI0_7/d_9_ XI11_4/XI0/XI0_7/d__9_ DECAP_INV_G11
XG8308 XI11_4/XI0/XI0_7/d_8_ XI11_4/XI0/XI0_7/d__8_ DECAP_INV_G11
XG8309 XI11_4/XI0/XI0_7/d_7_ XI11_4/XI0/XI0_7/d__7_ DECAP_INV_G11
XG8310 XI11_4/XI0/XI0_7/d_6_ XI11_4/XI0/XI0_7/d__6_ DECAP_INV_G11
XG8311 XI11_4/XI0/XI0_7/d_5_ XI11_4/XI0/XI0_7/d__5_ DECAP_INV_G11
XG8312 XI11_4/XI0/XI0_7/d_4_ XI11_4/XI0/XI0_7/d__4_ DECAP_INV_G11
XG8313 XI11_4/XI0/XI0_7/d_3_ XI11_4/XI0/XI0_7/d__3_ DECAP_INV_G11
XG8314 XI11_4/XI0/XI0_7/d_2_ XI11_4/XI0/XI0_7/d__2_ DECAP_INV_G11
XG8315 XI11_4/XI0/XI0_7/d_1_ XI11_4/XI0/XI0_7/d__1_ DECAP_INV_G11
XG8316 XI11_4/XI0/XI0_7/d_0_ XI11_4/XI0/XI0_7/d__0_ DECAP_INV_G11
XG8317 XI11_4/XI0/XI0_6/d__15_ XI11_4/XI0/XI0_6/d_15_ DECAP_INV_G11
XG8318 XI11_4/XI0/XI0_6/d__14_ XI11_4/XI0/XI0_6/d_14_ DECAP_INV_G11
XG8319 XI11_4/XI0/XI0_6/d__13_ XI11_4/XI0/XI0_6/d_13_ DECAP_INV_G11
XG8320 XI11_4/XI0/XI0_6/d__12_ XI11_4/XI0/XI0_6/d_12_ DECAP_INV_G11
XG8321 XI11_4/XI0/XI0_6/d__11_ XI11_4/XI0/XI0_6/d_11_ DECAP_INV_G11
XG8322 XI11_4/XI0/XI0_6/d__10_ XI11_4/XI0/XI0_6/d_10_ DECAP_INV_G11
XG8323 XI11_4/XI0/XI0_6/d__9_ XI11_4/XI0/XI0_6/d_9_ DECAP_INV_G11
XG8324 XI11_4/XI0/XI0_6/d__8_ XI11_4/XI0/XI0_6/d_8_ DECAP_INV_G11
XG8325 XI11_4/XI0/XI0_6/d__7_ XI11_4/XI0/XI0_6/d_7_ DECAP_INV_G11
XG8326 XI11_4/XI0/XI0_6/d__6_ XI11_4/XI0/XI0_6/d_6_ DECAP_INV_G11
XG8327 XI11_4/XI0/XI0_6/d__5_ XI11_4/XI0/XI0_6/d_5_ DECAP_INV_G11
XG8328 XI11_4/XI0/XI0_6/d__4_ XI11_4/XI0/XI0_6/d_4_ DECAP_INV_G11
XG8329 XI11_4/XI0/XI0_6/d__3_ XI11_4/XI0/XI0_6/d_3_ DECAP_INV_G11
XG8330 XI11_4/XI0/XI0_6/d__2_ XI11_4/XI0/XI0_6/d_2_ DECAP_INV_G11
XG8331 XI11_4/XI0/XI0_6/d__1_ XI11_4/XI0/XI0_6/d_1_ DECAP_INV_G11
XG8332 XI11_4/XI0/XI0_6/d__0_ XI11_4/XI0/XI0_6/d_0_ DECAP_INV_G11
XG8333 XI11_4/XI0/XI0_6/d_15_ XI11_4/XI0/XI0_6/d__15_ DECAP_INV_G11
XG8334 XI11_4/XI0/XI0_6/d_14_ XI11_4/XI0/XI0_6/d__14_ DECAP_INV_G11
XG8335 XI11_4/XI0/XI0_6/d_13_ XI11_4/XI0/XI0_6/d__13_ DECAP_INV_G11
XG8336 XI11_4/XI0/XI0_6/d_12_ XI11_4/XI0/XI0_6/d__12_ DECAP_INV_G11
XG8337 XI11_4/XI0/XI0_6/d_11_ XI11_4/XI0/XI0_6/d__11_ DECAP_INV_G11
XG8338 XI11_4/XI0/XI0_6/d_10_ XI11_4/XI0/XI0_6/d__10_ DECAP_INV_G11
XG8339 XI11_4/XI0/XI0_6/d_9_ XI11_4/XI0/XI0_6/d__9_ DECAP_INV_G11
XG8340 XI11_4/XI0/XI0_6/d_8_ XI11_4/XI0/XI0_6/d__8_ DECAP_INV_G11
XG8341 XI11_4/XI0/XI0_6/d_7_ XI11_4/XI0/XI0_6/d__7_ DECAP_INV_G11
XG8342 XI11_4/XI0/XI0_6/d_6_ XI11_4/XI0/XI0_6/d__6_ DECAP_INV_G11
XG8343 XI11_4/XI0/XI0_6/d_5_ XI11_4/XI0/XI0_6/d__5_ DECAP_INV_G11
XG8344 XI11_4/XI0/XI0_6/d_4_ XI11_4/XI0/XI0_6/d__4_ DECAP_INV_G11
XG8345 XI11_4/XI0/XI0_6/d_3_ XI11_4/XI0/XI0_6/d__3_ DECAP_INV_G11
XG8346 XI11_4/XI0/XI0_6/d_2_ XI11_4/XI0/XI0_6/d__2_ DECAP_INV_G11
XG8347 XI11_4/XI0/XI0_6/d_1_ XI11_4/XI0/XI0_6/d__1_ DECAP_INV_G11
XG8348 XI11_4/XI0/XI0_6/d_0_ XI11_4/XI0/XI0_6/d__0_ DECAP_INV_G11
XG8349 XI11_4/XI0/XI0_5/d__15_ XI11_4/XI0/XI0_5/d_15_ DECAP_INV_G11
XG8350 XI11_4/XI0/XI0_5/d__14_ XI11_4/XI0/XI0_5/d_14_ DECAP_INV_G11
XG8351 XI11_4/XI0/XI0_5/d__13_ XI11_4/XI0/XI0_5/d_13_ DECAP_INV_G11
XG8352 XI11_4/XI0/XI0_5/d__12_ XI11_4/XI0/XI0_5/d_12_ DECAP_INV_G11
XG8353 XI11_4/XI0/XI0_5/d__11_ XI11_4/XI0/XI0_5/d_11_ DECAP_INV_G11
XG8354 XI11_4/XI0/XI0_5/d__10_ XI11_4/XI0/XI0_5/d_10_ DECAP_INV_G11
XG8355 XI11_4/XI0/XI0_5/d__9_ XI11_4/XI0/XI0_5/d_9_ DECAP_INV_G11
XG8356 XI11_4/XI0/XI0_5/d__8_ XI11_4/XI0/XI0_5/d_8_ DECAP_INV_G11
XG8357 XI11_4/XI0/XI0_5/d__7_ XI11_4/XI0/XI0_5/d_7_ DECAP_INV_G11
XG8358 XI11_4/XI0/XI0_5/d__6_ XI11_4/XI0/XI0_5/d_6_ DECAP_INV_G11
XG8359 XI11_4/XI0/XI0_5/d__5_ XI11_4/XI0/XI0_5/d_5_ DECAP_INV_G11
XG8360 XI11_4/XI0/XI0_5/d__4_ XI11_4/XI0/XI0_5/d_4_ DECAP_INV_G11
XG8361 XI11_4/XI0/XI0_5/d__3_ XI11_4/XI0/XI0_5/d_3_ DECAP_INV_G11
XG8362 XI11_4/XI0/XI0_5/d__2_ XI11_4/XI0/XI0_5/d_2_ DECAP_INV_G11
XG8363 XI11_4/XI0/XI0_5/d__1_ XI11_4/XI0/XI0_5/d_1_ DECAP_INV_G11
XG8364 XI11_4/XI0/XI0_5/d__0_ XI11_4/XI0/XI0_5/d_0_ DECAP_INV_G11
XG8365 XI11_4/XI0/XI0_5/d_15_ XI11_4/XI0/XI0_5/d__15_ DECAP_INV_G11
XG8366 XI11_4/XI0/XI0_5/d_14_ XI11_4/XI0/XI0_5/d__14_ DECAP_INV_G11
XG8367 XI11_4/XI0/XI0_5/d_13_ XI11_4/XI0/XI0_5/d__13_ DECAP_INV_G11
XG8368 XI11_4/XI0/XI0_5/d_12_ XI11_4/XI0/XI0_5/d__12_ DECAP_INV_G11
XG8369 XI11_4/XI0/XI0_5/d_11_ XI11_4/XI0/XI0_5/d__11_ DECAP_INV_G11
XG8370 XI11_4/XI0/XI0_5/d_10_ XI11_4/XI0/XI0_5/d__10_ DECAP_INV_G11
XG8371 XI11_4/XI0/XI0_5/d_9_ XI11_4/XI0/XI0_5/d__9_ DECAP_INV_G11
XG8372 XI11_4/XI0/XI0_5/d_8_ XI11_4/XI0/XI0_5/d__8_ DECAP_INV_G11
XG8373 XI11_4/XI0/XI0_5/d_7_ XI11_4/XI0/XI0_5/d__7_ DECAP_INV_G11
XG8374 XI11_4/XI0/XI0_5/d_6_ XI11_4/XI0/XI0_5/d__6_ DECAP_INV_G11
XG8375 XI11_4/XI0/XI0_5/d_5_ XI11_4/XI0/XI0_5/d__5_ DECAP_INV_G11
XG8376 XI11_4/XI0/XI0_5/d_4_ XI11_4/XI0/XI0_5/d__4_ DECAP_INV_G11
XG8377 XI11_4/XI0/XI0_5/d_3_ XI11_4/XI0/XI0_5/d__3_ DECAP_INV_G11
XG8378 XI11_4/XI0/XI0_5/d_2_ XI11_4/XI0/XI0_5/d__2_ DECAP_INV_G11
XG8379 XI11_4/XI0/XI0_5/d_1_ XI11_4/XI0/XI0_5/d__1_ DECAP_INV_G11
XG8380 XI11_4/XI0/XI0_5/d_0_ XI11_4/XI0/XI0_5/d__0_ DECAP_INV_G11
XG8381 XI11_4/XI0/XI0_4/d__15_ XI11_4/XI0/XI0_4/d_15_ DECAP_INV_G11
XG8382 XI11_4/XI0/XI0_4/d__14_ XI11_4/XI0/XI0_4/d_14_ DECAP_INV_G11
XG8383 XI11_4/XI0/XI0_4/d__13_ XI11_4/XI0/XI0_4/d_13_ DECAP_INV_G11
XG8384 XI11_4/XI0/XI0_4/d__12_ XI11_4/XI0/XI0_4/d_12_ DECAP_INV_G11
XG8385 XI11_4/XI0/XI0_4/d__11_ XI11_4/XI0/XI0_4/d_11_ DECAP_INV_G11
XG8386 XI11_4/XI0/XI0_4/d__10_ XI11_4/XI0/XI0_4/d_10_ DECAP_INV_G11
XG8387 XI11_4/XI0/XI0_4/d__9_ XI11_4/XI0/XI0_4/d_9_ DECAP_INV_G11
XG8388 XI11_4/XI0/XI0_4/d__8_ XI11_4/XI0/XI0_4/d_8_ DECAP_INV_G11
XG8389 XI11_4/XI0/XI0_4/d__7_ XI11_4/XI0/XI0_4/d_7_ DECAP_INV_G11
XG8390 XI11_4/XI0/XI0_4/d__6_ XI11_4/XI0/XI0_4/d_6_ DECAP_INV_G11
XG8391 XI11_4/XI0/XI0_4/d__5_ XI11_4/XI0/XI0_4/d_5_ DECAP_INV_G11
XG8392 XI11_4/XI0/XI0_4/d__4_ XI11_4/XI0/XI0_4/d_4_ DECAP_INV_G11
XG8393 XI11_4/XI0/XI0_4/d__3_ XI11_4/XI0/XI0_4/d_3_ DECAP_INV_G11
XG8394 XI11_4/XI0/XI0_4/d__2_ XI11_4/XI0/XI0_4/d_2_ DECAP_INV_G11
XG8395 XI11_4/XI0/XI0_4/d__1_ XI11_4/XI0/XI0_4/d_1_ DECAP_INV_G11
XG8396 XI11_4/XI0/XI0_4/d__0_ XI11_4/XI0/XI0_4/d_0_ DECAP_INV_G11
XG8397 XI11_4/XI0/XI0_4/d_15_ XI11_4/XI0/XI0_4/d__15_ DECAP_INV_G11
XG8398 XI11_4/XI0/XI0_4/d_14_ XI11_4/XI0/XI0_4/d__14_ DECAP_INV_G11
XG8399 XI11_4/XI0/XI0_4/d_13_ XI11_4/XI0/XI0_4/d__13_ DECAP_INV_G11
XG8400 XI11_4/XI0/XI0_4/d_12_ XI11_4/XI0/XI0_4/d__12_ DECAP_INV_G11
XG8401 XI11_4/XI0/XI0_4/d_11_ XI11_4/XI0/XI0_4/d__11_ DECAP_INV_G11
XG8402 XI11_4/XI0/XI0_4/d_10_ XI11_4/XI0/XI0_4/d__10_ DECAP_INV_G11
XG8403 XI11_4/XI0/XI0_4/d_9_ XI11_4/XI0/XI0_4/d__9_ DECAP_INV_G11
XG8404 XI11_4/XI0/XI0_4/d_8_ XI11_4/XI0/XI0_4/d__8_ DECAP_INV_G11
XG8405 XI11_4/XI0/XI0_4/d_7_ XI11_4/XI0/XI0_4/d__7_ DECAP_INV_G11
XG8406 XI11_4/XI0/XI0_4/d_6_ XI11_4/XI0/XI0_4/d__6_ DECAP_INV_G11
XG8407 XI11_4/XI0/XI0_4/d_5_ XI11_4/XI0/XI0_4/d__5_ DECAP_INV_G11
XG8408 XI11_4/XI0/XI0_4/d_4_ XI11_4/XI0/XI0_4/d__4_ DECAP_INV_G11
XG8409 XI11_4/XI0/XI0_4/d_3_ XI11_4/XI0/XI0_4/d__3_ DECAP_INV_G11
XG8410 XI11_4/XI0/XI0_4/d_2_ XI11_4/XI0/XI0_4/d__2_ DECAP_INV_G11
XG8411 XI11_4/XI0/XI0_4/d_1_ XI11_4/XI0/XI0_4/d__1_ DECAP_INV_G11
XG8412 XI11_4/XI0/XI0_4/d_0_ XI11_4/XI0/XI0_4/d__0_ DECAP_INV_G11
XG8413 XI11_4/XI0/XI0_3/d__15_ XI11_4/XI0/XI0_3/d_15_ DECAP_INV_G11
XG8414 XI11_4/XI0/XI0_3/d__14_ XI11_4/XI0/XI0_3/d_14_ DECAP_INV_G11
XG8415 XI11_4/XI0/XI0_3/d__13_ XI11_4/XI0/XI0_3/d_13_ DECAP_INV_G11
XG8416 XI11_4/XI0/XI0_3/d__12_ XI11_4/XI0/XI0_3/d_12_ DECAP_INV_G11
XG8417 XI11_4/XI0/XI0_3/d__11_ XI11_4/XI0/XI0_3/d_11_ DECAP_INV_G11
XG8418 XI11_4/XI0/XI0_3/d__10_ XI11_4/XI0/XI0_3/d_10_ DECAP_INV_G11
XG8419 XI11_4/XI0/XI0_3/d__9_ XI11_4/XI0/XI0_3/d_9_ DECAP_INV_G11
XG8420 XI11_4/XI0/XI0_3/d__8_ XI11_4/XI0/XI0_3/d_8_ DECAP_INV_G11
XG8421 XI11_4/XI0/XI0_3/d__7_ XI11_4/XI0/XI0_3/d_7_ DECAP_INV_G11
XG8422 XI11_4/XI0/XI0_3/d__6_ XI11_4/XI0/XI0_3/d_6_ DECAP_INV_G11
XG8423 XI11_4/XI0/XI0_3/d__5_ XI11_4/XI0/XI0_3/d_5_ DECAP_INV_G11
XG8424 XI11_4/XI0/XI0_3/d__4_ XI11_4/XI0/XI0_3/d_4_ DECAP_INV_G11
XG8425 XI11_4/XI0/XI0_3/d__3_ XI11_4/XI0/XI0_3/d_3_ DECAP_INV_G11
XG8426 XI11_4/XI0/XI0_3/d__2_ XI11_4/XI0/XI0_3/d_2_ DECAP_INV_G11
XG8427 XI11_4/XI0/XI0_3/d__1_ XI11_4/XI0/XI0_3/d_1_ DECAP_INV_G11
XG8428 XI11_4/XI0/XI0_3/d__0_ XI11_4/XI0/XI0_3/d_0_ DECAP_INV_G11
XG8429 XI11_4/XI0/XI0_3/d_15_ XI11_4/XI0/XI0_3/d__15_ DECAP_INV_G11
XG8430 XI11_4/XI0/XI0_3/d_14_ XI11_4/XI0/XI0_3/d__14_ DECAP_INV_G11
XG8431 XI11_4/XI0/XI0_3/d_13_ XI11_4/XI0/XI0_3/d__13_ DECAP_INV_G11
XG8432 XI11_4/XI0/XI0_3/d_12_ XI11_4/XI0/XI0_3/d__12_ DECAP_INV_G11
XG8433 XI11_4/XI0/XI0_3/d_11_ XI11_4/XI0/XI0_3/d__11_ DECAP_INV_G11
XG8434 XI11_4/XI0/XI0_3/d_10_ XI11_4/XI0/XI0_3/d__10_ DECAP_INV_G11
XG8435 XI11_4/XI0/XI0_3/d_9_ XI11_4/XI0/XI0_3/d__9_ DECAP_INV_G11
XG8436 XI11_4/XI0/XI0_3/d_8_ XI11_4/XI0/XI0_3/d__8_ DECAP_INV_G11
XG8437 XI11_4/XI0/XI0_3/d_7_ XI11_4/XI0/XI0_3/d__7_ DECAP_INV_G11
XG8438 XI11_4/XI0/XI0_3/d_6_ XI11_4/XI0/XI0_3/d__6_ DECAP_INV_G11
XG8439 XI11_4/XI0/XI0_3/d_5_ XI11_4/XI0/XI0_3/d__5_ DECAP_INV_G11
XG8440 XI11_4/XI0/XI0_3/d_4_ XI11_4/XI0/XI0_3/d__4_ DECAP_INV_G11
XG8441 XI11_4/XI0/XI0_3/d_3_ XI11_4/XI0/XI0_3/d__3_ DECAP_INV_G11
XG8442 XI11_4/XI0/XI0_3/d_2_ XI11_4/XI0/XI0_3/d__2_ DECAP_INV_G11
XG8443 XI11_4/XI0/XI0_3/d_1_ XI11_4/XI0/XI0_3/d__1_ DECAP_INV_G11
XG8444 XI11_4/XI0/XI0_3/d_0_ XI11_4/XI0/XI0_3/d__0_ DECAP_INV_G11
XG8445 XI11_4/XI0/XI0_2/d__15_ XI11_4/XI0/XI0_2/d_15_ DECAP_INV_G11
XG8446 XI11_4/XI0/XI0_2/d__14_ XI11_4/XI0/XI0_2/d_14_ DECAP_INV_G11
XG8447 XI11_4/XI0/XI0_2/d__13_ XI11_4/XI0/XI0_2/d_13_ DECAP_INV_G11
XG8448 XI11_4/XI0/XI0_2/d__12_ XI11_4/XI0/XI0_2/d_12_ DECAP_INV_G11
XG8449 XI11_4/XI0/XI0_2/d__11_ XI11_4/XI0/XI0_2/d_11_ DECAP_INV_G11
XG8450 XI11_4/XI0/XI0_2/d__10_ XI11_4/XI0/XI0_2/d_10_ DECAP_INV_G11
XG8451 XI11_4/XI0/XI0_2/d__9_ XI11_4/XI0/XI0_2/d_9_ DECAP_INV_G11
XG8452 XI11_4/XI0/XI0_2/d__8_ XI11_4/XI0/XI0_2/d_8_ DECAP_INV_G11
XG8453 XI11_4/XI0/XI0_2/d__7_ XI11_4/XI0/XI0_2/d_7_ DECAP_INV_G11
XG8454 XI11_4/XI0/XI0_2/d__6_ XI11_4/XI0/XI0_2/d_6_ DECAP_INV_G11
XG8455 XI11_4/XI0/XI0_2/d__5_ XI11_4/XI0/XI0_2/d_5_ DECAP_INV_G11
XG8456 XI11_4/XI0/XI0_2/d__4_ XI11_4/XI0/XI0_2/d_4_ DECAP_INV_G11
XG8457 XI11_4/XI0/XI0_2/d__3_ XI11_4/XI0/XI0_2/d_3_ DECAP_INV_G11
XG8458 XI11_4/XI0/XI0_2/d__2_ XI11_4/XI0/XI0_2/d_2_ DECAP_INV_G11
XG8459 XI11_4/XI0/XI0_2/d__1_ XI11_4/XI0/XI0_2/d_1_ DECAP_INV_G11
XG8460 XI11_4/XI0/XI0_2/d__0_ XI11_4/XI0/XI0_2/d_0_ DECAP_INV_G11
XG8461 XI11_4/XI0/XI0_2/d_15_ XI11_4/XI0/XI0_2/d__15_ DECAP_INV_G11
XG8462 XI11_4/XI0/XI0_2/d_14_ XI11_4/XI0/XI0_2/d__14_ DECAP_INV_G11
XG8463 XI11_4/XI0/XI0_2/d_13_ XI11_4/XI0/XI0_2/d__13_ DECAP_INV_G11
XG8464 XI11_4/XI0/XI0_2/d_12_ XI11_4/XI0/XI0_2/d__12_ DECAP_INV_G11
XG8465 XI11_4/XI0/XI0_2/d_11_ XI11_4/XI0/XI0_2/d__11_ DECAP_INV_G11
XG8466 XI11_4/XI0/XI0_2/d_10_ XI11_4/XI0/XI0_2/d__10_ DECAP_INV_G11
XG8467 XI11_4/XI0/XI0_2/d_9_ XI11_4/XI0/XI0_2/d__9_ DECAP_INV_G11
XG8468 XI11_4/XI0/XI0_2/d_8_ XI11_4/XI0/XI0_2/d__8_ DECAP_INV_G11
XG8469 XI11_4/XI0/XI0_2/d_7_ XI11_4/XI0/XI0_2/d__7_ DECAP_INV_G11
XG8470 XI11_4/XI0/XI0_2/d_6_ XI11_4/XI0/XI0_2/d__6_ DECAP_INV_G11
XG8471 XI11_4/XI0/XI0_2/d_5_ XI11_4/XI0/XI0_2/d__5_ DECAP_INV_G11
XG8472 XI11_4/XI0/XI0_2/d_4_ XI11_4/XI0/XI0_2/d__4_ DECAP_INV_G11
XG8473 XI11_4/XI0/XI0_2/d_3_ XI11_4/XI0/XI0_2/d__3_ DECAP_INV_G11
XG8474 XI11_4/XI0/XI0_2/d_2_ XI11_4/XI0/XI0_2/d__2_ DECAP_INV_G11
XG8475 XI11_4/XI0/XI0_2/d_1_ XI11_4/XI0/XI0_2/d__1_ DECAP_INV_G11
XG8476 XI11_4/XI0/XI0_2/d_0_ XI11_4/XI0/XI0_2/d__0_ DECAP_INV_G11
XG8477 XI11_4/XI0/XI0_1/d__15_ XI11_4/XI0/XI0_1/d_15_ DECAP_INV_G11
XG8478 XI11_4/XI0/XI0_1/d__14_ XI11_4/XI0/XI0_1/d_14_ DECAP_INV_G11
XG8479 XI11_4/XI0/XI0_1/d__13_ XI11_4/XI0/XI0_1/d_13_ DECAP_INV_G11
XG8480 XI11_4/XI0/XI0_1/d__12_ XI11_4/XI0/XI0_1/d_12_ DECAP_INV_G11
XG8481 XI11_4/XI0/XI0_1/d__11_ XI11_4/XI0/XI0_1/d_11_ DECAP_INV_G11
XG8482 XI11_4/XI0/XI0_1/d__10_ XI11_4/XI0/XI0_1/d_10_ DECAP_INV_G11
XG8483 XI11_4/XI0/XI0_1/d__9_ XI11_4/XI0/XI0_1/d_9_ DECAP_INV_G11
XG8484 XI11_4/XI0/XI0_1/d__8_ XI11_4/XI0/XI0_1/d_8_ DECAP_INV_G11
XG8485 XI11_4/XI0/XI0_1/d__7_ XI11_4/XI0/XI0_1/d_7_ DECAP_INV_G11
XG8486 XI11_4/XI0/XI0_1/d__6_ XI11_4/XI0/XI0_1/d_6_ DECAP_INV_G11
XG8487 XI11_4/XI0/XI0_1/d__5_ XI11_4/XI0/XI0_1/d_5_ DECAP_INV_G11
XG8488 XI11_4/XI0/XI0_1/d__4_ XI11_4/XI0/XI0_1/d_4_ DECAP_INV_G11
XG8489 XI11_4/XI0/XI0_1/d__3_ XI11_4/XI0/XI0_1/d_3_ DECAP_INV_G11
XG8490 XI11_4/XI0/XI0_1/d__2_ XI11_4/XI0/XI0_1/d_2_ DECAP_INV_G11
XG8491 XI11_4/XI0/XI0_1/d__1_ XI11_4/XI0/XI0_1/d_1_ DECAP_INV_G11
XG8492 XI11_4/XI0/XI0_1/d__0_ XI11_4/XI0/XI0_1/d_0_ DECAP_INV_G11
XG8493 XI11_4/XI0/XI0_1/d_15_ XI11_4/XI0/XI0_1/d__15_ DECAP_INV_G11
XG8494 XI11_4/XI0/XI0_1/d_14_ XI11_4/XI0/XI0_1/d__14_ DECAP_INV_G11
XG8495 XI11_4/XI0/XI0_1/d_13_ XI11_4/XI0/XI0_1/d__13_ DECAP_INV_G11
XG8496 XI11_4/XI0/XI0_1/d_12_ XI11_4/XI0/XI0_1/d__12_ DECAP_INV_G11
XG8497 XI11_4/XI0/XI0_1/d_11_ XI11_4/XI0/XI0_1/d__11_ DECAP_INV_G11
XG8498 XI11_4/XI0/XI0_1/d_10_ XI11_4/XI0/XI0_1/d__10_ DECAP_INV_G11
XG8499 XI11_4/XI0/XI0_1/d_9_ XI11_4/XI0/XI0_1/d__9_ DECAP_INV_G11
XG8500 XI11_4/XI0/XI0_1/d_8_ XI11_4/XI0/XI0_1/d__8_ DECAP_INV_G11
XG8501 XI11_4/XI0/XI0_1/d_7_ XI11_4/XI0/XI0_1/d__7_ DECAP_INV_G11
XG8502 XI11_4/XI0/XI0_1/d_6_ XI11_4/XI0/XI0_1/d__6_ DECAP_INV_G11
XG8503 XI11_4/XI0/XI0_1/d_5_ XI11_4/XI0/XI0_1/d__5_ DECAP_INV_G11
XG8504 XI11_4/XI0/XI0_1/d_4_ XI11_4/XI0/XI0_1/d__4_ DECAP_INV_G11
XG8505 XI11_4/XI0/XI0_1/d_3_ XI11_4/XI0/XI0_1/d__3_ DECAP_INV_G11
XG8506 XI11_4/XI0/XI0_1/d_2_ XI11_4/XI0/XI0_1/d__2_ DECAP_INV_G11
XG8507 XI11_4/XI0/XI0_1/d_1_ XI11_4/XI0/XI0_1/d__1_ DECAP_INV_G11
XG8508 XI11_4/XI0/XI0_1/d_0_ XI11_4/XI0/XI0_1/d__0_ DECAP_INV_G11
XG8509 XI11_4/XI0/XI0_0/d__15_ XI11_4/XI0/XI0_0/d_15_ DECAP_INV_G11
XG8510 XI11_4/XI0/XI0_0/d__14_ XI11_4/XI0/XI0_0/d_14_ DECAP_INV_G11
XG8511 XI11_4/XI0/XI0_0/d__13_ XI11_4/XI0/XI0_0/d_13_ DECAP_INV_G11
XG8512 XI11_4/XI0/XI0_0/d__12_ XI11_4/XI0/XI0_0/d_12_ DECAP_INV_G11
XG8513 XI11_4/XI0/XI0_0/d__11_ XI11_4/XI0/XI0_0/d_11_ DECAP_INV_G11
XG8514 XI11_4/XI0/XI0_0/d__10_ XI11_4/XI0/XI0_0/d_10_ DECAP_INV_G11
XG8515 XI11_4/XI0/XI0_0/d__9_ XI11_4/XI0/XI0_0/d_9_ DECAP_INV_G11
XG8516 XI11_4/XI0/XI0_0/d__8_ XI11_4/XI0/XI0_0/d_8_ DECAP_INV_G11
XG8517 XI11_4/XI0/XI0_0/d__7_ XI11_4/XI0/XI0_0/d_7_ DECAP_INV_G11
XG8518 XI11_4/XI0/XI0_0/d__6_ XI11_4/XI0/XI0_0/d_6_ DECAP_INV_G11
XG8519 XI11_4/XI0/XI0_0/d__5_ XI11_4/XI0/XI0_0/d_5_ DECAP_INV_G11
XG8520 XI11_4/XI0/XI0_0/d__4_ XI11_4/XI0/XI0_0/d_4_ DECAP_INV_G11
XG8521 XI11_4/XI0/XI0_0/d__3_ XI11_4/XI0/XI0_0/d_3_ DECAP_INV_G11
XG8522 XI11_4/XI0/XI0_0/d__2_ XI11_4/XI0/XI0_0/d_2_ DECAP_INV_G11
XG8523 XI11_4/XI0/XI0_0/d__1_ XI11_4/XI0/XI0_0/d_1_ DECAP_INV_G11
XG8524 XI11_4/XI0/XI0_0/d__0_ XI11_4/XI0/XI0_0/d_0_ DECAP_INV_G11
XG8525 XI11_4/XI0/XI0_0/d_15_ XI11_4/XI0/XI0_0/d__15_ DECAP_INV_G11
XG8526 XI11_4/XI0/XI0_0/d_14_ XI11_4/XI0/XI0_0/d__14_ DECAP_INV_G11
XG8527 XI11_4/XI0/XI0_0/d_13_ XI11_4/XI0/XI0_0/d__13_ DECAP_INV_G11
XG8528 XI11_4/XI0/XI0_0/d_12_ XI11_4/XI0/XI0_0/d__12_ DECAP_INV_G11
XG8529 XI11_4/XI0/XI0_0/d_11_ XI11_4/XI0/XI0_0/d__11_ DECAP_INV_G11
XG8530 XI11_4/XI0/XI0_0/d_10_ XI11_4/XI0/XI0_0/d__10_ DECAP_INV_G11
XG8531 XI11_4/XI0/XI0_0/d_9_ XI11_4/XI0/XI0_0/d__9_ DECAP_INV_G11
XG8532 XI11_4/XI0/XI0_0/d_8_ XI11_4/XI0/XI0_0/d__8_ DECAP_INV_G11
XG8533 XI11_4/XI0/XI0_0/d_7_ XI11_4/XI0/XI0_0/d__7_ DECAP_INV_G11
XG8534 XI11_4/XI0/XI0_0/d_6_ XI11_4/XI0/XI0_0/d__6_ DECAP_INV_G11
XG8535 XI11_4/XI0/XI0_0/d_5_ XI11_4/XI0/XI0_0/d__5_ DECAP_INV_G11
XG8536 XI11_4/XI0/XI0_0/d_4_ XI11_4/XI0/XI0_0/d__4_ DECAP_INV_G11
XG8537 XI11_4/XI0/XI0_0/d_3_ XI11_4/XI0/XI0_0/d__3_ DECAP_INV_G11
XG8538 XI11_4/XI0/XI0_0/d_2_ XI11_4/XI0/XI0_0/d__2_ DECAP_INV_G11
XG8539 XI11_4/XI0/XI0_0/d_1_ XI11_4/XI0/XI0_0/d__1_ DECAP_INV_G11
XG8540 XI11_4/XI0/XI0_0/d_0_ XI11_4/XI0/XI0_0/d__0_ DECAP_INV_G11
XG8541 XI11_3/XI3/net17 XI11_3/XI3/net5 DECAP_INV_G7
XG8542 XI11_3/XI3/net5 XI11_3/preck DECAP_INV_G8
XG8543 sck_bar XI11_3/XI3/net018 DECAP_INV_G9
XG8544 XI11_3/XI3/net018 XI11_3/XI3/net012 DECAP_INV_G9
XG8545 XI11_3/XI3/net014 XI11_3/XI3/net7 DECAP_INV_G9
XG8546 XI11_3/XI3/net012 XI11_3/XI3/net014 DECAP_INV_G9
XG8547 XI11_3/XI4/net063 XI11_3/XI4/net0112 DECAP_INV_G10
XG8548 XI11_3/XI4/net26 XI11_3/XI4/net089 DECAP_INV_G10
XG8549 XI11_3/XI4/data_out XI11_3/XI4/data_out_ DECAP_INV_G10
XG8550 XI11_3/XI4/net20 XI11_3/XI4/net0103 DECAP_INV_G10
XG8551 XI11_3/net12 XI11_3/XI4/net32 DECAP_INV_G7
XG8552 XI11_3/net9 XI11_3/XI4/net52 DECAP_INV_G7
XG8553 XI11_3/XI4/data_out_ XI11_3/XI4/data_out DECAP_INV_G10
XG8554 XI11_3/XI0/XI0_63/d__15_ XI11_3/XI0/XI0_63/d_15_ DECAP_INV_G11
XG8555 XI11_3/XI0/XI0_63/d__14_ XI11_3/XI0/XI0_63/d_14_ DECAP_INV_G11
XG8556 XI11_3/XI0/XI0_63/d__13_ XI11_3/XI0/XI0_63/d_13_ DECAP_INV_G11
XG8557 XI11_3/XI0/XI0_63/d__12_ XI11_3/XI0/XI0_63/d_12_ DECAP_INV_G11
XG8558 XI11_3/XI0/XI0_63/d__11_ XI11_3/XI0/XI0_63/d_11_ DECAP_INV_G11
XG8559 XI11_3/XI0/XI0_63/d__10_ XI11_3/XI0/XI0_63/d_10_ DECAP_INV_G11
XG8560 XI11_3/XI0/XI0_63/d__9_ XI11_3/XI0/XI0_63/d_9_ DECAP_INV_G11
XG8561 XI11_3/XI0/XI0_63/d__8_ XI11_3/XI0/XI0_63/d_8_ DECAP_INV_G11
XG8562 XI11_3/XI0/XI0_63/d__7_ XI11_3/XI0/XI0_63/d_7_ DECAP_INV_G11
XG8563 XI11_3/XI0/XI0_63/d__6_ XI11_3/XI0/XI0_63/d_6_ DECAP_INV_G11
XG8564 XI11_3/XI0/XI0_63/d__5_ XI11_3/XI0/XI0_63/d_5_ DECAP_INV_G11
XG8565 XI11_3/XI0/XI0_63/d__4_ XI11_3/XI0/XI0_63/d_4_ DECAP_INV_G11
XG8566 XI11_3/XI0/XI0_63/d__3_ XI11_3/XI0/XI0_63/d_3_ DECAP_INV_G11
XG8567 XI11_3/XI0/XI0_63/d__2_ XI11_3/XI0/XI0_63/d_2_ DECAP_INV_G11
XG8568 XI11_3/XI0/XI0_63/d__1_ XI11_3/XI0/XI0_63/d_1_ DECAP_INV_G11
XG8569 XI11_3/XI0/XI0_63/d__0_ XI11_3/XI0/XI0_63/d_0_ DECAP_INV_G11
XG8570 XI11_3/XI0/XI0_63/d_15_ XI11_3/XI0/XI0_63/d__15_ DECAP_INV_G11
XG8571 XI11_3/XI0/XI0_63/d_14_ XI11_3/XI0/XI0_63/d__14_ DECAP_INV_G11
XG8572 XI11_3/XI0/XI0_63/d_13_ XI11_3/XI0/XI0_63/d__13_ DECAP_INV_G11
XG8573 XI11_3/XI0/XI0_63/d_12_ XI11_3/XI0/XI0_63/d__12_ DECAP_INV_G11
XG8574 XI11_3/XI0/XI0_63/d_11_ XI11_3/XI0/XI0_63/d__11_ DECAP_INV_G11
XG8575 XI11_3/XI0/XI0_63/d_10_ XI11_3/XI0/XI0_63/d__10_ DECAP_INV_G11
XG8576 XI11_3/XI0/XI0_63/d_9_ XI11_3/XI0/XI0_63/d__9_ DECAP_INV_G11
XG8577 XI11_3/XI0/XI0_63/d_8_ XI11_3/XI0/XI0_63/d__8_ DECAP_INV_G11
XG8578 XI11_3/XI0/XI0_63/d_7_ XI11_3/XI0/XI0_63/d__7_ DECAP_INV_G11
XG8579 XI11_3/XI0/XI0_63/d_6_ XI11_3/XI0/XI0_63/d__6_ DECAP_INV_G11
XG8580 XI11_3/XI0/XI0_63/d_5_ XI11_3/XI0/XI0_63/d__5_ DECAP_INV_G11
XG8581 XI11_3/XI0/XI0_63/d_4_ XI11_3/XI0/XI0_63/d__4_ DECAP_INV_G11
XG8582 XI11_3/XI0/XI0_63/d_3_ XI11_3/XI0/XI0_63/d__3_ DECAP_INV_G11
XG8583 XI11_3/XI0/XI0_63/d_2_ XI11_3/XI0/XI0_63/d__2_ DECAP_INV_G11
XG8584 XI11_3/XI0/XI0_63/d_1_ XI11_3/XI0/XI0_63/d__1_ DECAP_INV_G11
XG8585 XI11_3/XI0/XI0_63/d_0_ XI11_3/XI0/XI0_63/d__0_ DECAP_INV_G11
XG8586 XI11_3/XI0/XI0_62/d__15_ XI11_3/XI0/XI0_62/d_15_ DECAP_INV_G11
XG8587 XI11_3/XI0/XI0_62/d__14_ XI11_3/XI0/XI0_62/d_14_ DECAP_INV_G11
XG8588 XI11_3/XI0/XI0_62/d__13_ XI11_3/XI0/XI0_62/d_13_ DECAP_INV_G11
XG8589 XI11_3/XI0/XI0_62/d__12_ XI11_3/XI0/XI0_62/d_12_ DECAP_INV_G11
XG8590 XI11_3/XI0/XI0_62/d__11_ XI11_3/XI0/XI0_62/d_11_ DECAP_INV_G11
XG8591 XI11_3/XI0/XI0_62/d__10_ XI11_3/XI0/XI0_62/d_10_ DECAP_INV_G11
XG8592 XI11_3/XI0/XI0_62/d__9_ XI11_3/XI0/XI0_62/d_9_ DECAP_INV_G11
XG8593 XI11_3/XI0/XI0_62/d__8_ XI11_3/XI0/XI0_62/d_8_ DECAP_INV_G11
XG8594 XI11_3/XI0/XI0_62/d__7_ XI11_3/XI0/XI0_62/d_7_ DECAP_INV_G11
XG8595 XI11_3/XI0/XI0_62/d__6_ XI11_3/XI0/XI0_62/d_6_ DECAP_INV_G11
XG8596 XI11_3/XI0/XI0_62/d__5_ XI11_3/XI0/XI0_62/d_5_ DECAP_INV_G11
XG8597 XI11_3/XI0/XI0_62/d__4_ XI11_3/XI0/XI0_62/d_4_ DECAP_INV_G11
XG8598 XI11_3/XI0/XI0_62/d__3_ XI11_3/XI0/XI0_62/d_3_ DECAP_INV_G11
XG8599 XI11_3/XI0/XI0_62/d__2_ XI11_3/XI0/XI0_62/d_2_ DECAP_INV_G11
XG8600 XI11_3/XI0/XI0_62/d__1_ XI11_3/XI0/XI0_62/d_1_ DECAP_INV_G11
XG8601 XI11_3/XI0/XI0_62/d__0_ XI11_3/XI0/XI0_62/d_0_ DECAP_INV_G11
XG8602 XI11_3/XI0/XI0_62/d_15_ XI11_3/XI0/XI0_62/d__15_ DECAP_INV_G11
XG8603 XI11_3/XI0/XI0_62/d_14_ XI11_3/XI0/XI0_62/d__14_ DECAP_INV_G11
XG8604 XI11_3/XI0/XI0_62/d_13_ XI11_3/XI0/XI0_62/d__13_ DECAP_INV_G11
XG8605 XI11_3/XI0/XI0_62/d_12_ XI11_3/XI0/XI0_62/d__12_ DECAP_INV_G11
XG8606 XI11_3/XI0/XI0_62/d_11_ XI11_3/XI0/XI0_62/d__11_ DECAP_INV_G11
XG8607 XI11_3/XI0/XI0_62/d_10_ XI11_3/XI0/XI0_62/d__10_ DECAP_INV_G11
XG8608 XI11_3/XI0/XI0_62/d_9_ XI11_3/XI0/XI0_62/d__9_ DECAP_INV_G11
XG8609 XI11_3/XI0/XI0_62/d_8_ XI11_3/XI0/XI0_62/d__8_ DECAP_INV_G11
XG8610 XI11_3/XI0/XI0_62/d_7_ XI11_3/XI0/XI0_62/d__7_ DECAP_INV_G11
XG8611 XI11_3/XI0/XI0_62/d_6_ XI11_3/XI0/XI0_62/d__6_ DECAP_INV_G11
XG8612 XI11_3/XI0/XI0_62/d_5_ XI11_3/XI0/XI0_62/d__5_ DECAP_INV_G11
XG8613 XI11_3/XI0/XI0_62/d_4_ XI11_3/XI0/XI0_62/d__4_ DECAP_INV_G11
XG8614 XI11_3/XI0/XI0_62/d_3_ XI11_3/XI0/XI0_62/d__3_ DECAP_INV_G11
XG8615 XI11_3/XI0/XI0_62/d_2_ XI11_3/XI0/XI0_62/d__2_ DECAP_INV_G11
XG8616 XI11_3/XI0/XI0_62/d_1_ XI11_3/XI0/XI0_62/d__1_ DECAP_INV_G11
XG8617 XI11_3/XI0/XI0_62/d_0_ XI11_3/XI0/XI0_62/d__0_ DECAP_INV_G11
XG8618 XI11_3/XI0/XI0_61/d__15_ XI11_3/XI0/XI0_61/d_15_ DECAP_INV_G11
XG8619 XI11_3/XI0/XI0_61/d__14_ XI11_3/XI0/XI0_61/d_14_ DECAP_INV_G11
XG8620 XI11_3/XI0/XI0_61/d__13_ XI11_3/XI0/XI0_61/d_13_ DECAP_INV_G11
XG8621 XI11_3/XI0/XI0_61/d__12_ XI11_3/XI0/XI0_61/d_12_ DECAP_INV_G11
XG8622 XI11_3/XI0/XI0_61/d__11_ XI11_3/XI0/XI0_61/d_11_ DECAP_INV_G11
XG8623 XI11_3/XI0/XI0_61/d__10_ XI11_3/XI0/XI0_61/d_10_ DECAP_INV_G11
XG8624 XI11_3/XI0/XI0_61/d__9_ XI11_3/XI0/XI0_61/d_9_ DECAP_INV_G11
XG8625 XI11_3/XI0/XI0_61/d__8_ XI11_3/XI0/XI0_61/d_8_ DECAP_INV_G11
XG8626 XI11_3/XI0/XI0_61/d__7_ XI11_3/XI0/XI0_61/d_7_ DECAP_INV_G11
XG8627 XI11_3/XI0/XI0_61/d__6_ XI11_3/XI0/XI0_61/d_6_ DECAP_INV_G11
XG8628 XI11_3/XI0/XI0_61/d__5_ XI11_3/XI0/XI0_61/d_5_ DECAP_INV_G11
XG8629 XI11_3/XI0/XI0_61/d__4_ XI11_3/XI0/XI0_61/d_4_ DECAP_INV_G11
XG8630 XI11_3/XI0/XI0_61/d__3_ XI11_3/XI0/XI0_61/d_3_ DECAP_INV_G11
XG8631 XI11_3/XI0/XI0_61/d__2_ XI11_3/XI0/XI0_61/d_2_ DECAP_INV_G11
XG8632 XI11_3/XI0/XI0_61/d__1_ XI11_3/XI0/XI0_61/d_1_ DECAP_INV_G11
XG8633 XI11_3/XI0/XI0_61/d__0_ XI11_3/XI0/XI0_61/d_0_ DECAP_INV_G11
XG8634 XI11_3/XI0/XI0_61/d_15_ XI11_3/XI0/XI0_61/d__15_ DECAP_INV_G11
XG8635 XI11_3/XI0/XI0_61/d_14_ XI11_3/XI0/XI0_61/d__14_ DECAP_INV_G11
XG8636 XI11_3/XI0/XI0_61/d_13_ XI11_3/XI0/XI0_61/d__13_ DECAP_INV_G11
XG8637 XI11_3/XI0/XI0_61/d_12_ XI11_3/XI0/XI0_61/d__12_ DECAP_INV_G11
XG8638 XI11_3/XI0/XI0_61/d_11_ XI11_3/XI0/XI0_61/d__11_ DECAP_INV_G11
XG8639 XI11_3/XI0/XI0_61/d_10_ XI11_3/XI0/XI0_61/d__10_ DECAP_INV_G11
XG8640 XI11_3/XI0/XI0_61/d_9_ XI11_3/XI0/XI0_61/d__9_ DECAP_INV_G11
XG8641 XI11_3/XI0/XI0_61/d_8_ XI11_3/XI0/XI0_61/d__8_ DECAP_INV_G11
XG8642 XI11_3/XI0/XI0_61/d_7_ XI11_3/XI0/XI0_61/d__7_ DECAP_INV_G11
XG8643 XI11_3/XI0/XI0_61/d_6_ XI11_3/XI0/XI0_61/d__6_ DECAP_INV_G11
XG8644 XI11_3/XI0/XI0_61/d_5_ XI11_3/XI0/XI0_61/d__5_ DECAP_INV_G11
XG8645 XI11_3/XI0/XI0_61/d_4_ XI11_3/XI0/XI0_61/d__4_ DECAP_INV_G11
XG8646 XI11_3/XI0/XI0_61/d_3_ XI11_3/XI0/XI0_61/d__3_ DECAP_INV_G11
XG8647 XI11_3/XI0/XI0_61/d_2_ XI11_3/XI0/XI0_61/d__2_ DECAP_INV_G11
XG8648 XI11_3/XI0/XI0_61/d_1_ XI11_3/XI0/XI0_61/d__1_ DECAP_INV_G11
XG8649 XI11_3/XI0/XI0_61/d_0_ XI11_3/XI0/XI0_61/d__0_ DECAP_INV_G11
XG8650 XI11_3/XI0/XI0_60/d__15_ XI11_3/XI0/XI0_60/d_15_ DECAP_INV_G11
XG8651 XI11_3/XI0/XI0_60/d__14_ XI11_3/XI0/XI0_60/d_14_ DECAP_INV_G11
XG8652 XI11_3/XI0/XI0_60/d__13_ XI11_3/XI0/XI0_60/d_13_ DECAP_INV_G11
XG8653 XI11_3/XI0/XI0_60/d__12_ XI11_3/XI0/XI0_60/d_12_ DECAP_INV_G11
XG8654 XI11_3/XI0/XI0_60/d__11_ XI11_3/XI0/XI0_60/d_11_ DECAP_INV_G11
XG8655 XI11_3/XI0/XI0_60/d__10_ XI11_3/XI0/XI0_60/d_10_ DECAP_INV_G11
XG8656 XI11_3/XI0/XI0_60/d__9_ XI11_3/XI0/XI0_60/d_9_ DECAP_INV_G11
XG8657 XI11_3/XI0/XI0_60/d__8_ XI11_3/XI0/XI0_60/d_8_ DECAP_INV_G11
XG8658 XI11_3/XI0/XI0_60/d__7_ XI11_3/XI0/XI0_60/d_7_ DECAP_INV_G11
XG8659 XI11_3/XI0/XI0_60/d__6_ XI11_3/XI0/XI0_60/d_6_ DECAP_INV_G11
XG8660 XI11_3/XI0/XI0_60/d__5_ XI11_3/XI0/XI0_60/d_5_ DECAP_INV_G11
XG8661 XI11_3/XI0/XI0_60/d__4_ XI11_3/XI0/XI0_60/d_4_ DECAP_INV_G11
XG8662 XI11_3/XI0/XI0_60/d__3_ XI11_3/XI0/XI0_60/d_3_ DECAP_INV_G11
XG8663 XI11_3/XI0/XI0_60/d__2_ XI11_3/XI0/XI0_60/d_2_ DECAP_INV_G11
XG8664 XI11_3/XI0/XI0_60/d__1_ XI11_3/XI0/XI0_60/d_1_ DECAP_INV_G11
XG8665 XI11_3/XI0/XI0_60/d__0_ XI11_3/XI0/XI0_60/d_0_ DECAP_INV_G11
XG8666 XI11_3/XI0/XI0_60/d_15_ XI11_3/XI0/XI0_60/d__15_ DECAP_INV_G11
XG8667 XI11_3/XI0/XI0_60/d_14_ XI11_3/XI0/XI0_60/d__14_ DECAP_INV_G11
XG8668 XI11_3/XI0/XI0_60/d_13_ XI11_3/XI0/XI0_60/d__13_ DECAP_INV_G11
XG8669 XI11_3/XI0/XI0_60/d_12_ XI11_3/XI0/XI0_60/d__12_ DECAP_INV_G11
XG8670 XI11_3/XI0/XI0_60/d_11_ XI11_3/XI0/XI0_60/d__11_ DECAP_INV_G11
XG8671 XI11_3/XI0/XI0_60/d_10_ XI11_3/XI0/XI0_60/d__10_ DECAP_INV_G11
XG8672 XI11_3/XI0/XI0_60/d_9_ XI11_3/XI0/XI0_60/d__9_ DECAP_INV_G11
XG8673 XI11_3/XI0/XI0_60/d_8_ XI11_3/XI0/XI0_60/d__8_ DECAP_INV_G11
XG8674 XI11_3/XI0/XI0_60/d_7_ XI11_3/XI0/XI0_60/d__7_ DECAP_INV_G11
XG8675 XI11_3/XI0/XI0_60/d_6_ XI11_3/XI0/XI0_60/d__6_ DECAP_INV_G11
XG8676 XI11_3/XI0/XI0_60/d_5_ XI11_3/XI0/XI0_60/d__5_ DECAP_INV_G11
XG8677 XI11_3/XI0/XI0_60/d_4_ XI11_3/XI0/XI0_60/d__4_ DECAP_INV_G11
XG8678 XI11_3/XI0/XI0_60/d_3_ XI11_3/XI0/XI0_60/d__3_ DECAP_INV_G11
XG8679 XI11_3/XI0/XI0_60/d_2_ XI11_3/XI0/XI0_60/d__2_ DECAP_INV_G11
XG8680 XI11_3/XI0/XI0_60/d_1_ XI11_3/XI0/XI0_60/d__1_ DECAP_INV_G11
XG8681 XI11_3/XI0/XI0_60/d_0_ XI11_3/XI0/XI0_60/d__0_ DECAP_INV_G11
XG8682 XI11_3/XI0/XI0_59/d__15_ XI11_3/XI0/XI0_59/d_15_ DECAP_INV_G11
XG8683 XI11_3/XI0/XI0_59/d__14_ XI11_3/XI0/XI0_59/d_14_ DECAP_INV_G11
XG8684 XI11_3/XI0/XI0_59/d__13_ XI11_3/XI0/XI0_59/d_13_ DECAP_INV_G11
XG8685 XI11_3/XI0/XI0_59/d__12_ XI11_3/XI0/XI0_59/d_12_ DECAP_INV_G11
XG8686 XI11_3/XI0/XI0_59/d__11_ XI11_3/XI0/XI0_59/d_11_ DECAP_INV_G11
XG8687 XI11_3/XI0/XI0_59/d__10_ XI11_3/XI0/XI0_59/d_10_ DECAP_INV_G11
XG8688 XI11_3/XI0/XI0_59/d__9_ XI11_3/XI0/XI0_59/d_9_ DECAP_INV_G11
XG8689 XI11_3/XI0/XI0_59/d__8_ XI11_3/XI0/XI0_59/d_8_ DECAP_INV_G11
XG8690 XI11_3/XI0/XI0_59/d__7_ XI11_3/XI0/XI0_59/d_7_ DECAP_INV_G11
XG8691 XI11_3/XI0/XI0_59/d__6_ XI11_3/XI0/XI0_59/d_6_ DECAP_INV_G11
XG8692 XI11_3/XI0/XI0_59/d__5_ XI11_3/XI0/XI0_59/d_5_ DECAP_INV_G11
XG8693 XI11_3/XI0/XI0_59/d__4_ XI11_3/XI0/XI0_59/d_4_ DECAP_INV_G11
XG8694 XI11_3/XI0/XI0_59/d__3_ XI11_3/XI0/XI0_59/d_3_ DECAP_INV_G11
XG8695 XI11_3/XI0/XI0_59/d__2_ XI11_3/XI0/XI0_59/d_2_ DECAP_INV_G11
XG8696 XI11_3/XI0/XI0_59/d__1_ XI11_3/XI0/XI0_59/d_1_ DECAP_INV_G11
XG8697 XI11_3/XI0/XI0_59/d__0_ XI11_3/XI0/XI0_59/d_0_ DECAP_INV_G11
XG8698 XI11_3/XI0/XI0_59/d_15_ XI11_3/XI0/XI0_59/d__15_ DECAP_INV_G11
XG8699 XI11_3/XI0/XI0_59/d_14_ XI11_3/XI0/XI0_59/d__14_ DECAP_INV_G11
XG8700 XI11_3/XI0/XI0_59/d_13_ XI11_3/XI0/XI0_59/d__13_ DECAP_INV_G11
XG8701 XI11_3/XI0/XI0_59/d_12_ XI11_3/XI0/XI0_59/d__12_ DECAP_INV_G11
XG8702 XI11_3/XI0/XI0_59/d_11_ XI11_3/XI0/XI0_59/d__11_ DECAP_INV_G11
XG8703 XI11_3/XI0/XI0_59/d_10_ XI11_3/XI0/XI0_59/d__10_ DECAP_INV_G11
XG8704 XI11_3/XI0/XI0_59/d_9_ XI11_3/XI0/XI0_59/d__9_ DECAP_INV_G11
XG8705 XI11_3/XI0/XI0_59/d_8_ XI11_3/XI0/XI0_59/d__8_ DECAP_INV_G11
XG8706 XI11_3/XI0/XI0_59/d_7_ XI11_3/XI0/XI0_59/d__7_ DECAP_INV_G11
XG8707 XI11_3/XI0/XI0_59/d_6_ XI11_3/XI0/XI0_59/d__6_ DECAP_INV_G11
XG8708 XI11_3/XI0/XI0_59/d_5_ XI11_3/XI0/XI0_59/d__5_ DECAP_INV_G11
XG8709 XI11_3/XI0/XI0_59/d_4_ XI11_3/XI0/XI0_59/d__4_ DECAP_INV_G11
XG8710 XI11_3/XI0/XI0_59/d_3_ XI11_3/XI0/XI0_59/d__3_ DECAP_INV_G11
XG8711 XI11_3/XI0/XI0_59/d_2_ XI11_3/XI0/XI0_59/d__2_ DECAP_INV_G11
XG8712 XI11_3/XI0/XI0_59/d_1_ XI11_3/XI0/XI0_59/d__1_ DECAP_INV_G11
XG8713 XI11_3/XI0/XI0_59/d_0_ XI11_3/XI0/XI0_59/d__0_ DECAP_INV_G11
XG8714 XI11_3/XI0/XI0_58/d__15_ XI11_3/XI0/XI0_58/d_15_ DECAP_INV_G11
XG8715 XI11_3/XI0/XI0_58/d__14_ XI11_3/XI0/XI0_58/d_14_ DECAP_INV_G11
XG8716 XI11_3/XI0/XI0_58/d__13_ XI11_3/XI0/XI0_58/d_13_ DECAP_INV_G11
XG8717 XI11_3/XI0/XI0_58/d__12_ XI11_3/XI0/XI0_58/d_12_ DECAP_INV_G11
XG8718 XI11_3/XI0/XI0_58/d__11_ XI11_3/XI0/XI0_58/d_11_ DECAP_INV_G11
XG8719 XI11_3/XI0/XI0_58/d__10_ XI11_3/XI0/XI0_58/d_10_ DECAP_INV_G11
XG8720 XI11_3/XI0/XI0_58/d__9_ XI11_3/XI0/XI0_58/d_9_ DECAP_INV_G11
XG8721 XI11_3/XI0/XI0_58/d__8_ XI11_3/XI0/XI0_58/d_8_ DECAP_INV_G11
XG8722 XI11_3/XI0/XI0_58/d__7_ XI11_3/XI0/XI0_58/d_7_ DECAP_INV_G11
XG8723 XI11_3/XI0/XI0_58/d__6_ XI11_3/XI0/XI0_58/d_6_ DECAP_INV_G11
XG8724 XI11_3/XI0/XI0_58/d__5_ XI11_3/XI0/XI0_58/d_5_ DECAP_INV_G11
XG8725 XI11_3/XI0/XI0_58/d__4_ XI11_3/XI0/XI0_58/d_4_ DECAP_INV_G11
XG8726 XI11_3/XI0/XI0_58/d__3_ XI11_3/XI0/XI0_58/d_3_ DECAP_INV_G11
XG8727 XI11_3/XI0/XI0_58/d__2_ XI11_3/XI0/XI0_58/d_2_ DECAP_INV_G11
XG8728 XI11_3/XI0/XI0_58/d__1_ XI11_3/XI0/XI0_58/d_1_ DECAP_INV_G11
XG8729 XI11_3/XI0/XI0_58/d__0_ XI11_3/XI0/XI0_58/d_0_ DECAP_INV_G11
XG8730 XI11_3/XI0/XI0_58/d_15_ XI11_3/XI0/XI0_58/d__15_ DECAP_INV_G11
XG8731 XI11_3/XI0/XI0_58/d_14_ XI11_3/XI0/XI0_58/d__14_ DECAP_INV_G11
XG8732 XI11_3/XI0/XI0_58/d_13_ XI11_3/XI0/XI0_58/d__13_ DECAP_INV_G11
XG8733 XI11_3/XI0/XI0_58/d_12_ XI11_3/XI0/XI0_58/d__12_ DECAP_INV_G11
XG8734 XI11_3/XI0/XI0_58/d_11_ XI11_3/XI0/XI0_58/d__11_ DECAP_INV_G11
XG8735 XI11_3/XI0/XI0_58/d_10_ XI11_3/XI0/XI0_58/d__10_ DECAP_INV_G11
XG8736 XI11_3/XI0/XI0_58/d_9_ XI11_3/XI0/XI0_58/d__9_ DECAP_INV_G11
XG8737 XI11_3/XI0/XI0_58/d_8_ XI11_3/XI0/XI0_58/d__8_ DECAP_INV_G11
XG8738 XI11_3/XI0/XI0_58/d_7_ XI11_3/XI0/XI0_58/d__7_ DECAP_INV_G11
XG8739 XI11_3/XI0/XI0_58/d_6_ XI11_3/XI0/XI0_58/d__6_ DECAP_INV_G11
XG8740 XI11_3/XI0/XI0_58/d_5_ XI11_3/XI0/XI0_58/d__5_ DECAP_INV_G11
XG8741 XI11_3/XI0/XI0_58/d_4_ XI11_3/XI0/XI0_58/d__4_ DECAP_INV_G11
XG8742 XI11_3/XI0/XI0_58/d_3_ XI11_3/XI0/XI0_58/d__3_ DECAP_INV_G11
XG8743 XI11_3/XI0/XI0_58/d_2_ XI11_3/XI0/XI0_58/d__2_ DECAP_INV_G11
XG8744 XI11_3/XI0/XI0_58/d_1_ XI11_3/XI0/XI0_58/d__1_ DECAP_INV_G11
XG8745 XI11_3/XI0/XI0_58/d_0_ XI11_3/XI0/XI0_58/d__0_ DECAP_INV_G11
XG8746 XI11_3/XI0/XI0_57/d__15_ XI11_3/XI0/XI0_57/d_15_ DECAP_INV_G11
XG8747 XI11_3/XI0/XI0_57/d__14_ XI11_3/XI0/XI0_57/d_14_ DECAP_INV_G11
XG8748 XI11_3/XI0/XI0_57/d__13_ XI11_3/XI0/XI0_57/d_13_ DECAP_INV_G11
XG8749 XI11_3/XI0/XI0_57/d__12_ XI11_3/XI0/XI0_57/d_12_ DECAP_INV_G11
XG8750 XI11_3/XI0/XI0_57/d__11_ XI11_3/XI0/XI0_57/d_11_ DECAP_INV_G11
XG8751 XI11_3/XI0/XI0_57/d__10_ XI11_3/XI0/XI0_57/d_10_ DECAP_INV_G11
XG8752 XI11_3/XI0/XI0_57/d__9_ XI11_3/XI0/XI0_57/d_9_ DECAP_INV_G11
XG8753 XI11_3/XI0/XI0_57/d__8_ XI11_3/XI0/XI0_57/d_8_ DECAP_INV_G11
XG8754 XI11_3/XI0/XI0_57/d__7_ XI11_3/XI0/XI0_57/d_7_ DECAP_INV_G11
XG8755 XI11_3/XI0/XI0_57/d__6_ XI11_3/XI0/XI0_57/d_6_ DECAP_INV_G11
XG8756 XI11_3/XI0/XI0_57/d__5_ XI11_3/XI0/XI0_57/d_5_ DECAP_INV_G11
XG8757 XI11_3/XI0/XI0_57/d__4_ XI11_3/XI0/XI0_57/d_4_ DECAP_INV_G11
XG8758 XI11_3/XI0/XI0_57/d__3_ XI11_3/XI0/XI0_57/d_3_ DECAP_INV_G11
XG8759 XI11_3/XI0/XI0_57/d__2_ XI11_3/XI0/XI0_57/d_2_ DECAP_INV_G11
XG8760 XI11_3/XI0/XI0_57/d__1_ XI11_3/XI0/XI0_57/d_1_ DECAP_INV_G11
XG8761 XI11_3/XI0/XI0_57/d__0_ XI11_3/XI0/XI0_57/d_0_ DECAP_INV_G11
XG8762 XI11_3/XI0/XI0_57/d_15_ XI11_3/XI0/XI0_57/d__15_ DECAP_INV_G11
XG8763 XI11_3/XI0/XI0_57/d_14_ XI11_3/XI0/XI0_57/d__14_ DECAP_INV_G11
XG8764 XI11_3/XI0/XI0_57/d_13_ XI11_3/XI0/XI0_57/d__13_ DECAP_INV_G11
XG8765 XI11_3/XI0/XI0_57/d_12_ XI11_3/XI0/XI0_57/d__12_ DECAP_INV_G11
XG8766 XI11_3/XI0/XI0_57/d_11_ XI11_3/XI0/XI0_57/d__11_ DECAP_INV_G11
XG8767 XI11_3/XI0/XI0_57/d_10_ XI11_3/XI0/XI0_57/d__10_ DECAP_INV_G11
XG8768 XI11_3/XI0/XI0_57/d_9_ XI11_3/XI0/XI0_57/d__9_ DECAP_INV_G11
XG8769 XI11_3/XI0/XI0_57/d_8_ XI11_3/XI0/XI0_57/d__8_ DECAP_INV_G11
XG8770 XI11_3/XI0/XI0_57/d_7_ XI11_3/XI0/XI0_57/d__7_ DECAP_INV_G11
XG8771 XI11_3/XI0/XI0_57/d_6_ XI11_3/XI0/XI0_57/d__6_ DECAP_INV_G11
XG8772 XI11_3/XI0/XI0_57/d_5_ XI11_3/XI0/XI0_57/d__5_ DECAP_INV_G11
XG8773 XI11_3/XI0/XI0_57/d_4_ XI11_3/XI0/XI0_57/d__4_ DECAP_INV_G11
XG8774 XI11_3/XI0/XI0_57/d_3_ XI11_3/XI0/XI0_57/d__3_ DECAP_INV_G11
XG8775 XI11_3/XI0/XI0_57/d_2_ XI11_3/XI0/XI0_57/d__2_ DECAP_INV_G11
XG8776 XI11_3/XI0/XI0_57/d_1_ XI11_3/XI0/XI0_57/d__1_ DECAP_INV_G11
XG8777 XI11_3/XI0/XI0_57/d_0_ XI11_3/XI0/XI0_57/d__0_ DECAP_INV_G11
XG8778 XI11_3/XI0/XI0_56/d__15_ XI11_3/XI0/XI0_56/d_15_ DECAP_INV_G11
XG8779 XI11_3/XI0/XI0_56/d__14_ XI11_3/XI0/XI0_56/d_14_ DECAP_INV_G11
XG8780 XI11_3/XI0/XI0_56/d__13_ XI11_3/XI0/XI0_56/d_13_ DECAP_INV_G11
XG8781 XI11_3/XI0/XI0_56/d__12_ XI11_3/XI0/XI0_56/d_12_ DECAP_INV_G11
XG8782 XI11_3/XI0/XI0_56/d__11_ XI11_3/XI0/XI0_56/d_11_ DECAP_INV_G11
XG8783 XI11_3/XI0/XI0_56/d__10_ XI11_3/XI0/XI0_56/d_10_ DECAP_INV_G11
XG8784 XI11_3/XI0/XI0_56/d__9_ XI11_3/XI0/XI0_56/d_9_ DECAP_INV_G11
XG8785 XI11_3/XI0/XI0_56/d__8_ XI11_3/XI0/XI0_56/d_8_ DECAP_INV_G11
XG8786 XI11_3/XI0/XI0_56/d__7_ XI11_3/XI0/XI0_56/d_7_ DECAP_INV_G11
XG8787 XI11_3/XI0/XI0_56/d__6_ XI11_3/XI0/XI0_56/d_6_ DECAP_INV_G11
XG8788 XI11_3/XI0/XI0_56/d__5_ XI11_3/XI0/XI0_56/d_5_ DECAP_INV_G11
XG8789 XI11_3/XI0/XI0_56/d__4_ XI11_3/XI0/XI0_56/d_4_ DECAP_INV_G11
XG8790 XI11_3/XI0/XI0_56/d__3_ XI11_3/XI0/XI0_56/d_3_ DECAP_INV_G11
XG8791 XI11_3/XI0/XI0_56/d__2_ XI11_3/XI0/XI0_56/d_2_ DECAP_INV_G11
XG8792 XI11_3/XI0/XI0_56/d__1_ XI11_3/XI0/XI0_56/d_1_ DECAP_INV_G11
XG8793 XI11_3/XI0/XI0_56/d__0_ XI11_3/XI0/XI0_56/d_0_ DECAP_INV_G11
XG8794 XI11_3/XI0/XI0_56/d_15_ XI11_3/XI0/XI0_56/d__15_ DECAP_INV_G11
XG8795 XI11_3/XI0/XI0_56/d_14_ XI11_3/XI0/XI0_56/d__14_ DECAP_INV_G11
XG8796 XI11_3/XI0/XI0_56/d_13_ XI11_3/XI0/XI0_56/d__13_ DECAP_INV_G11
XG8797 XI11_3/XI0/XI0_56/d_12_ XI11_3/XI0/XI0_56/d__12_ DECAP_INV_G11
XG8798 XI11_3/XI0/XI0_56/d_11_ XI11_3/XI0/XI0_56/d__11_ DECAP_INV_G11
XG8799 XI11_3/XI0/XI0_56/d_10_ XI11_3/XI0/XI0_56/d__10_ DECAP_INV_G11
XG8800 XI11_3/XI0/XI0_56/d_9_ XI11_3/XI0/XI0_56/d__9_ DECAP_INV_G11
XG8801 XI11_3/XI0/XI0_56/d_8_ XI11_3/XI0/XI0_56/d__8_ DECAP_INV_G11
XG8802 XI11_3/XI0/XI0_56/d_7_ XI11_3/XI0/XI0_56/d__7_ DECAP_INV_G11
XG8803 XI11_3/XI0/XI0_56/d_6_ XI11_3/XI0/XI0_56/d__6_ DECAP_INV_G11
XG8804 XI11_3/XI0/XI0_56/d_5_ XI11_3/XI0/XI0_56/d__5_ DECAP_INV_G11
XG8805 XI11_3/XI0/XI0_56/d_4_ XI11_3/XI0/XI0_56/d__4_ DECAP_INV_G11
XG8806 XI11_3/XI0/XI0_56/d_3_ XI11_3/XI0/XI0_56/d__3_ DECAP_INV_G11
XG8807 XI11_3/XI0/XI0_56/d_2_ XI11_3/XI0/XI0_56/d__2_ DECAP_INV_G11
XG8808 XI11_3/XI0/XI0_56/d_1_ XI11_3/XI0/XI0_56/d__1_ DECAP_INV_G11
XG8809 XI11_3/XI0/XI0_56/d_0_ XI11_3/XI0/XI0_56/d__0_ DECAP_INV_G11
XG8810 XI11_3/XI0/XI0_55/d__15_ XI11_3/XI0/XI0_55/d_15_ DECAP_INV_G11
XG8811 XI11_3/XI0/XI0_55/d__14_ XI11_3/XI0/XI0_55/d_14_ DECAP_INV_G11
XG8812 XI11_3/XI0/XI0_55/d__13_ XI11_3/XI0/XI0_55/d_13_ DECAP_INV_G11
XG8813 XI11_3/XI0/XI0_55/d__12_ XI11_3/XI0/XI0_55/d_12_ DECAP_INV_G11
XG8814 XI11_3/XI0/XI0_55/d__11_ XI11_3/XI0/XI0_55/d_11_ DECAP_INV_G11
XG8815 XI11_3/XI0/XI0_55/d__10_ XI11_3/XI0/XI0_55/d_10_ DECAP_INV_G11
XG8816 XI11_3/XI0/XI0_55/d__9_ XI11_3/XI0/XI0_55/d_9_ DECAP_INV_G11
XG8817 XI11_3/XI0/XI0_55/d__8_ XI11_3/XI0/XI0_55/d_8_ DECAP_INV_G11
XG8818 XI11_3/XI0/XI0_55/d__7_ XI11_3/XI0/XI0_55/d_7_ DECAP_INV_G11
XG8819 XI11_3/XI0/XI0_55/d__6_ XI11_3/XI0/XI0_55/d_6_ DECAP_INV_G11
XG8820 XI11_3/XI0/XI0_55/d__5_ XI11_3/XI0/XI0_55/d_5_ DECAP_INV_G11
XG8821 XI11_3/XI0/XI0_55/d__4_ XI11_3/XI0/XI0_55/d_4_ DECAP_INV_G11
XG8822 XI11_3/XI0/XI0_55/d__3_ XI11_3/XI0/XI0_55/d_3_ DECAP_INV_G11
XG8823 XI11_3/XI0/XI0_55/d__2_ XI11_3/XI0/XI0_55/d_2_ DECAP_INV_G11
XG8824 XI11_3/XI0/XI0_55/d__1_ XI11_3/XI0/XI0_55/d_1_ DECAP_INV_G11
XG8825 XI11_3/XI0/XI0_55/d__0_ XI11_3/XI0/XI0_55/d_0_ DECAP_INV_G11
XG8826 XI11_3/XI0/XI0_55/d_15_ XI11_3/XI0/XI0_55/d__15_ DECAP_INV_G11
XG8827 XI11_3/XI0/XI0_55/d_14_ XI11_3/XI0/XI0_55/d__14_ DECAP_INV_G11
XG8828 XI11_3/XI0/XI0_55/d_13_ XI11_3/XI0/XI0_55/d__13_ DECAP_INV_G11
XG8829 XI11_3/XI0/XI0_55/d_12_ XI11_3/XI0/XI0_55/d__12_ DECAP_INV_G11
XG8830 XI11_3/XI0/XI0_55/d_11_ XI11_3/XI0/XI0_55/d__11_ DECAP_INV_G11
XG8831 XI11_3/XI0/XI0_55/d_10_ XI11_3/XI0/XI0_55/d__10_ DECAP_INV_G11
XG8832 XI11_3/XI0/XI0_55/d_9_ XI11_3/XI0/XI0_55/d__9_ DECAP_INV_G11
XG8833 XI11_3/XI0/XI0_55/d_8_ XI11_3/XI0/XI0_55/d__8_ DECAP_INV_G11
XG8834 XI11_3/XI0/XI0_55/d_7_ XI11_3/XI0/XI0_55/d__7_ DECAP_INV_G11
XG8835 XI11_3/XI0/XI0_55/d_6_ XI11_3/XI0/XI0_55/d__6_ DECAP_INV_G11
XG8836 XI11_3/XI0/XI0_55/d_5_ XI11_3/XI0/XI0_55/d__5_ DECAP_INV_G11
XG8837 XI11_3/XI0/XI0_55/d_4_ XI11_3/XI0/XI0_55/d__4_ DECAP_INV_G11
XG8838 XI11_3/XI0/XI0_55/d_3_ XI11_3/XI0/XI0_55/d__3_ DECAP_INV_G11
XG8839 XI11_3/XI0/XI0_55/d_2_ XI11_3/XI0/XI0_55/d__2_ DECAP_INV_G11
XG8840 XI11_3/XI0/XI0_55/d_1_ XI11_3/XI0/XI0_55/d__1_ DECAP_INV_G11
XG8841 XI11_3/XI0/XI0_55/d_0_ XI11_3/XI0/XI0_55/d__0_ DECAP_INV_G11
XG8842 XI11_3/XI0/XI0_54/d__15_ XI11_3/XI0/XI0_54/d_15_ DECAP_INV_G11
XG8843 XI11_3/XI0/XI0_54/d__14_ XI11_3/XI0/XI0_54/d_14_ DECAP_INV_G11
XG8844 XI11_3/XI0/XI0_54/d__13_ XI11_3/XI0/XI0_54/d_13_ DECAP_INV_G11
XG8845 XI11_3/XI0/XI0_54/d__12_ XI11_3/XI0/XI0_54/d_12_ DECAP_INV_G11
XG8846 XI11_3/XI0/XI0_54/d__11_ XI11_3/XI0/XI0_54/d_11_ DECAP_INV_G11
XG8847 XI11_3/XI0/XI0_54/d__10_ XI11_3/XI0/XI0_54/d_10_ DECAP_INV_G11
XG8848 XI11_3/XI0/XI0_54/d__9_ XI11_3/XI0/XI0_54/d_9_ DECAP_INV_G11
XG8849 XI11_3/XI0/XI0_54/d__8_ XI11_3/XI0/XI0_54/d_8_ DECAP_INV_G11
XG8850 XI11_3/XI0/XI0_54/d__7_ XI11_3/XI0/XI0_54/d_7_ DECAP_INV_G11
XG8851 XI11_3/XI0/XI0_54/d__6_ XI11_3/XI0/XI0_54/d_6_ DECAP_INV_G11
XG8852 XI11_3/XI0/XI0_54/d__5_ XI11_3/XI0/XI0_54/d_5_ DECAP_INV_G11
XG8853 XI11_3/XI0/XI0_54/d__4_ XI11_3/XI0/XI0_54/d_4_ DECAP_INV_G11
XG8854 XI11_3/XI0/XI0_54/d__3_ XI11_3/XI0/XI0_54/d_3_ DECAP_INV_G11
XG8855 XI11_3/XI0/XI0_54/d__2_ XI11_3/XI0/XI0_54/d_2_ DECAP_INV_G11
XG8856 XI11_3/XI0/XI0_54/d__1_ XI11_3/XI0/XI0_54/d_1_ DECAP_INV_G11
XG8857 XI11_3/XI0/XI0_54/d__0_ XI11_3/XI0/XI0_54/d_0_ DECAP_INV_G11
XG8858 XI11_3/XI0/XI0_54/d_15_ XI11_3/XI0/XI0_54/d__15_ DECAP_INV_G11
XG8859 XI11_3/XI0/XI0_54/d_14_ XI11_3/XI0/XI0_54/d__14_ DECAP_INV_G11
XG8860 XI11_3/XI0/XI0_54/d_13_ XI11_3/XI0/XI0_54/d__13_ DECAP_INV_G11
XG8861 XI11_3/XI0/XI0_54/d_12_ XI11_3/XI0/XI0_54/d__12_ DECAP_INV_G11
XG8862 XI11_3/XI0/XI0_54/d_11_ XI11_3/XI0/XI0_54/d__11_ DECAP_INV_G11
XG8863 XI11_3/XI0/XI0_54/d_10_ XI11_3/XI0/XI0_54/d__10_ DECAP_INV_G11
XG8864 XI11_3/XI0/XI0_54/d_9_ XI11_3/XI0/XI0_54/d__9_ DECAP_INV_G11
XG8865 XI11_3/XI0/XI0_54/d_8_ XI11_3/XI0/XI0_54/d__8_ DECAP_INV_G11
XG8866 XI11_3/XI0/XI0_54/d_7_ XI11_3/XI0/XI0_54/d__7_ DECAP_INV_G11
XG8867 XI11_3/XI0/XI0_54/d_6_ XI11_3/XI0/XI0_54/d__6_ DECAP_INV_G11
XG8868 XI11_3/XI0/XI0_54/d_5_ XI11_3/XI0/XI0_54/d__5_ DECAP_INV_G11
XG8869 XI11_3/XI0/XI0_54/d_4_ XI11_3/XI0/XI0_54/d__4_ DECAP_INV_G11
XG8870 XI11_3/XI0/XI0_54/d_3_ XI11_3/XI0/XI0_54/d__3_ DECAP_INV_G11
XG8871 XI11_3/XI0/XI0_54/d_2_ XI11_3/XI0/XI0_54/d__2_ DECAP_INV_G11
XG8872 XI11_3/XI0/XI0_54/d_1_ XI11_3/XI0/XI0_54/d__1_ DECAP_INV_G11
XG8873 XI11_3/XI0/XI0_54/d_0_ XI11_3/XI0/XI0_54/d__0_ DECAP_INV_G11
XG8874 XI11_3/XI0/XI0_53/d__15_ XI11_3/XI0/XI0_53/d_15_ DECAP_INV_G11
XG8875 XI11_3/XI0/XI0_53/d__14_ XI11_3/XI0/XI0_53/d_14_ DECAP_INV_G11
XG8876 XI11_3/XI0/XI0_53/d__13_ XI11_3/XI0/XI0_53/d_13_ DECAP_INV_G11
XG8877 XI11_3/XI0/XI0_53/d__12_ XI11_3/XI0/XI0_53/d_12_ DECAP_INV_G11
XG8878 XI11_3/XI0/XI0_53/d__11_ XI11_3/XI0/XI0_53/d_11_ DECAP_INV_G11
XG8879 XI11_3/XI0/XI0_53/d__10_ XI11_3/XI0/XI0_53/d_10_ DECAP_INV_G11
XG8880 XI11_3/XI0/XI0_53/d__9_ XI11_3/XI0/XI0_53/d_9_ DECAP_INV_G11
XG8881 XI11_3/XI0/XI0_53/d__8_ XI11_3/XI0/XI0_53/d_8_ DECAP_INV_G11
XG8882 XI11_3/XI0/XI0_53/d__7_ XI11_3/XI0/XI0_53/d_7_ DECAP_INV_G11
XG8883 XI11_3/XI0/XI0_53/d__6_ XI11_3/XI0/XI0_53/d_6_ DECAP_INV_G11
XG8884 XI11_3/XI0/XI0_53/d__5_ XI11_3/XI0/XI0_53/d_5_ DECAP_INV_G11
XG8885 XI11_3/XI0/XI0_53/d__4_ XI11_3/XI0/XI0_53/d_4_ DECAP_INV_G11
XG8886 XI11_3/XI0/XI0_53/d__3_ XI11_3/XI0/XI0_53/d_3_ DECAP_INV_G11
XG8887 XI11_3/XI0/XI0_53/d__2_ XI11_3/XI0/XI0_53/d_2_ DECAP_INV_G11
XG8888 XI11_3/XI0/XI0_53/d__1_ XI11_3/XI0/XI0_53/d_1_ DECAP_INV_G11
XG8889 XI11_3/XI0/XI0_53/d__0_ XI11_3/XI0/XI0_53/d_0_ DECAP_INV_G11
XG8890 XI11_3/XI0/XI0_53/d_15_ XI11_3/XI0/XI0_53/d__15_ DECAP_INV_G11
XG8891 XI11_3/XI0/XI0_53/d_14_ XI11_3/XI0/XI0_53/d__14_ DECAP_INV_G11
XG8892 XI11_3/XI0/XI0_53/d_13_ XI11_3/XI0/XI0_53/d__13_ DECAP_INV_G11
XG8893 XI11_3/XI0/XI0_53/d_12_ XI11_3/XI0/XI0_53/d__12_ DECAP_INV_G11
XG8894 XI11_3/XI0/XI0_53/d_11_ XI11_3/XI0/XI0_53/d__11_ DECAP_INV_G11
XG8895 XI11_3/XI0/XI0_53/d_10_ XI11_3/XI0/XI0_53/d__10_ DECAP_INV_G11
XG8896 XI11_3/XI0/XI0_53/d_9_ XI11_3/XI0/XI0_53/d__9_ DECAP_INV_G11
XG8897 XI11_3/XI0/XI0_53/d_8_ XI11_3/XI0/XI0_53/d__8_ DECAP_INV_G11
XG8898 XI11_3/XI0/XI0_53/d_7_ XI11_3/XI0/XI0_53/d__7_ DECAP_INV_G11
XG8899 XI11_3/XI0/XI0_53/d_6_ XI11_3/XI0/XI0_53/d__6_ DECAP_INV_G11
XG8900 XI11_3/XI0/XI0_53/d_5_ XI11_3/XI0/XI0_53/d__5_ DECAP_INV_G11
XG8901 XI11_3/XI0/XI0_53/d_4_ XI11_3/XI0/XI0_53/d__4_ DECAP_INV_G11
XG8902 XI11_3/XI0/XI0_53/d_3_ XI11_3/XI0/XI0_53/d__3_ DECAP_INV_G11
XG8903 XI11_3/XI0/XI0_53/d_2_ XI11_3/XI0/XI0_53/d__2_ DECAP_INV_G11
XG8904 XI11_3/XI0/XI0_53/d_1_ XI11_3/XI0/XI0_53/d__1_ DECAP_INV_G11
XG8905 XI11_3/XI0/XI0_53/d_0_ XI11_3/XI0/XI0_53/d__0_ DECAP_INV_G11
XG8906 XI11_3/XI0/XI0_52/d__15_ XI11_3/XI0/XI0_52/d_15_ DECAP_INV_G11
XG8907 XI11_3/XI0/XI0_52/d__14_ XI11_3/XI0/XI0_52/d_14_ DECAP_INV_G11
XG8908 XI11_3/XI0/XI0_52/d__13_ XI11_3/XI0/XI0_52/d_13_ DECAP_INV_G11
XG8909 XI11_3/XI0/XI0_52/d__12_ XI11_3/XI0/XI0_52/d_12_ DECAP_INV_G11
XG8910 XI11_3/XI0/XI0_52/d__11_ XI11_3/XI0/XI0_52/d_11_ DECAP_INV_G11
XG8911 XI11_3/XI0/XI0_52/d__10_ XI11_3/XI0/XI0_52/d_10_ DECAP_INV_G11
XG8912 XI11_3/XI0/XI0_52/d__9_ XI11_3/XI0/XI0_52/d_9_ DECAP_INV_G11
XG8913 XI11_3/XI0/XI0_52/d__8_ XI11_3/XI0/XI0_52/d_8_ DECAP_INV_G11
XG8914 XI11_3/XI0/XI0_52/d__7_ XI11_3/XI0/XI0_52/d_7_ DECAP_INV_G11
XG8915 XI11_3/XI0/XI0_52/d__6_ XI11_3/XI0/XI0_52/d_6_ DECAP_INV_G11
XG8916 XI11_3/XI0/XI0_52/d__5_ XI11_3/XI0/XI0_52/d_5_ DECAP_INV_G11
XG8917 XI11_3/XI0/XI0_52/d__4_ XI11_3/XI0/XI0_52/d_4_ DECAP_INV_G11
XG8918 XI11_3/XI0/XI0_52/d__3_ XI11_3/XI0/XI0_52/d_3_ DECAP_INV_G11
XG8919 XI11_3/XI0/XI0_52/d__2_ XI11_3/XI0/XI0_52/d_2_ DECAP_INV_G11
XG8920 XI11_3/XI0/XI0_52/d__1_ XI11_3/XI0/XI0_52/d_1_ DECAP_INV_G11
XG8921 XI11_3/XI0/XI0_52/d__0_ XI11_3/XI0/XI0_52/d_0_ DECAP_INV_G11
XG8922 XI11_3/XI0/XI0_52/d_15_ XI11_3/XI0/XI0_52/d__15_ DECAP_INV_G11
XG8923 XI11_3/XI0/XI0_52/d_14_ XI11_3/XI0/XI0_52/d__14_ DECAP_INV_G11
XG8924 XI11_3/XI0/XI0_52/d_13_ XI11_3/XI0/XI0_52/d__13_ DECAP_INV_G11
XG8925 XI11_3/XI0/XI0_52/d_12_ XI11_3/XI0/XI0_52/d__12_ DECAP_INV_G11
XG8926 XI11_3/XI0/XI0_52/d_11_ XI11_3/XI0/XI0_52/d__11_ DECAP_INV_G11
XG8927 XI11_3/XI0/XI0_52/d_10_ XI11_3/XI0/XI0_52/d__10_ DECAP_INV_G11
XG8928 XI11_3/XI0/XI0_52/d_9_ XI11_3/XI0/XI0_52/d__9_ DECAP_INV_G11
XG8929 XI11_3/XI0/XI0_52/d_8_ XI11_3/XI0/XI0_52/d__8_ DECAP_INV_G11
XG8930 XI11_3/XI0/XI0_52/d_7_ XI11_3/XI0/XI0_52/d__7_ DECAP_INV_G11
XG8931 XI11_3/XI0/XI0_52/d_6_ XI11_3/XI0/XI0_52/d__6_ DECAP_INV_G11
XG8932 XI11_3/XI0/XI0_52/d_5_ XI11_3/XI0/XI0_52/d__5_ DECAP_INV_G11
XG8933 XI11_3/XI0/XI0_52/d_4_ XI11_3/XI0/XI0_52/d__4_ DECAP_INV_G11
XG8934 XI11_3/XI0/XI0_52/d_3_ XI11_3/XI0/XI0_52/d__3_ DECAP_INV_G11
XG8935 XI11_3/XI0/XI0_52/d_2_ XI11_3/XI0/XI0_52/d__2_ DECAP_INV_G11
XG8936 XI11_3/XI0/XI0_52/d_1_ XI11_3/XI0/XI0_52/d__1_ DECAP_INV_G11
XG8937 XI11_3/XI0/XI0_52/d_0_ XI11_3/XI0/XI0_52/d__0_ DECAP_INV_G11
XG8938 XI11_3/XI0/XI0_51/d__15_ XI11_3/XI0/XI0_51/d_15_ DECAP_INV_G11
XG8939 XI11_3/XI0/XI0_51/d__14_ XI11_3/XI0/XI0_51/d_14_ DECAP_INV_G11
XG8940 XI11_3/XI0/XI0_51/d__13_ XI11_3/XI0/XI0_51/d_13_ DECAP_INV_G11
XG8941 XI11_3/XI0/XI0_51/d__12_ XI11_3/XI0/XI0_51/d_12_ DECAP_INV_G11
XG8942 XI11_3/XI0/XI0_51/d__11_ XI11_3/XI0/XI0_51/d_11_ DECAP_INV_G11
XG8943 XI11_3/XI0/XI0_51/d__10_ XI11_3/XI0/XI0_51/d_10_ DECAP_INV_G11
XG8944 XI11_3/XI0/XI0_51/d__9_ XI11_3/XI0/XI0_51/d_9_ DECAP_INV_G11
XG8945 XI11_3/XI0/XI0_51/d__8_ XI11_3/XI0/XI0_51/d_8_ DECAP_INV_G11
XG8946 XI11_3/XI0/XI0_51/d__7_ XI11_3/XI0/XI0_51/d_7_ DECAP_INV_G11
XG8947 XI11_3/XI0/XI0_51/d__6_ XI11_3/XI0/XI0_51/d_6_ DECAP_INV_G11
XG8948 XI11_3/XI0/XI0_51/d__5_ XI11_3/XI0/XI0_51/d_5_ DECAP_INV_G11
XG8949 XI11_3/XI0/XI0_51/d__4_ XI11_3/XI0/XI0_51/d_4_ DECAP_INV_G11
XG8950 XI11_3/XI0/XI0_51/d__3_ XI11_3/XI0/XI0_51/d_3_ DECAP_INV_G11
XG8951 XI11_3/XI0/XI0_51/d__2_ XI11_3/XI0/XI0_51/d_2_ DECAP_INV_G11
XG8952 XI11_3/XI0/XI0_51/d__1_ XI11_3/XI0/XI0_51/d_1_ DECAP_INV_G11
XG8953 XI11_3/XI0/XI0_51/d__0_ XI11_3/XI0/XI0_51/d_0_ DECAP_INV_G11
XG8954 XI11_3/XI0/XI0_51/d_15_ XI11_3/XI0/XI0_51/d__15_ DECAP_INV_G11
XG8955 XI11_3/XI0/XI0_51/d_14_ XI11_3/XI0/XI0_51/d__14_ DECAP_INV_G11
XG8956 XI11_3/XI0/XI0_51/d_13_ XI11_3/XI0/XI0_51/d__13_ DECAP_INV_G11
XG8957 XI11_3/XI0/XI0_51/d_12_ XI11_3/XI0/XI0_51/d__12_ DECAP_INV_G11
XG8958 XI11_3/XI0/XI0_51/d_11_ XI11_3/XI0/XI0_51/d__11_ DECAP_INV_G11
XG8959 XI11_3/XI0/XI0_51/d_10_ XI11_3/XI0/XI0_51/d__10_ DECAP_INV_G11
XG8960 XI11_3/XI0/XI0_51/d_9_ XI11_3/XI0/XI0_51/d__9_ DECAP_INV_G11
XG8961 XI11_3/XI0/XI0_51/d_8_ XI11_3/XI0/XI0_51/d__8_ DECAP_INV_G11
XG8962 XI11_3/XI0/XI0_51/d_7_ XI11_3/XI0/XI0_51/d__7_ DECAP_INV_G11
XG8963 XI11_3/XI0/XI0_51/d_6_ XI11_3/XI0/XI0_51/d__6_ DECAP_INV_G11
XG8964 XI11_3/XI0/XI0_51/d_5_ XI11_3/XI0/XI0_51/d__5_ DECAP_INV_G11
XG8965 XI11_3/XI0/XI0_51/d_4_ XI11_3/XI0/XI0_51/d__4_ DECAP_INV_G11
XG8966 XI11_3/XI0/XI0_51/d_3_ XI11_3/XI0/XI0_51/d__3_ DECAP_INV_G11
XG8967 XI11_3/XI0/XI0_51/d_2_ XI11_3/XI0/XI0_51/d__2_ DECAP_INV_G11
XG8968 XI11_3/XI0/XI0_51/d_1_ XI11_3/XI0/XI0_51/d__1_ DECAP_INV_G11
XG8969 XI11_3/XI0/XI0_51/d_0_ XI11_3/XI0/XI0_51/d__0_ DECAP_INV_G11
XG8970 XI11_3/XI0/XI0_50/d__15_ XI11_3/XI0/XI0_50/d_15_ DECAP_INV_G11
XG8971 XI11_3/XI0/XI0_50/d__14_ XI11_3/XI0/XI0_50/d_14_ DECAP_INV_G11
XG8972 XI11_3/XI0/XI0_50/d__13_ XI11_3/XI0/XI0_50/d_13_ DECAP_INV_G11
XG8973 XI11_3/XI0/XI0_50/d__12_ XI11_3/XI0/XI0_50/d_12_ DECAP_INV_G11
XG8974 XI11_3/XI0/XI0_50/d__11_ XI11_3/XI0/XI0_50/d_11_ DECAP_INV_G11
XG8975 XI11_3/XI0/XI0_50/d__10_ XI11_3/XI0/XI0_50/d_10_ DECAP_INV_G11
XG8976 XI11_3/XI0/XI0_50/d__9_ XI11_3/XI0/XI0_50/d_9_ DECAP_INV_G11
XG8977 XI11_3/XI0/XI0_50/d__8_ XI11_3/XI0/XI0_50/d_8_ DECAP_INV_G11
XG8978 XI11_3/XI0/XI0_50/d__7_ XI11_3/XI0/XI0_50/d_7_ DECAP_INV_G11
XG8979 XI11_3/XI0/XI0_50/d__6_ XI11_3/XI0/XI0_50/d_6_ DECAP_INV_G11
XG8980 XI11_3/XI0/XI0_50/d__5_ XI11_3/XI0/XI0_50/d_5_ DECAP_INV_G11
XG8981 XI11_3/XI0/XI0_50/d__4_ XI11_3/XI0/XI0_50/d_4_ DECAP_INV_G11
XG8982 XI11_3/XI0/XI0_50/d__3_ XI11_3/XI0/XI0_50/d_3_ DECAP_INV_G11
XG8983 XI11_3/XI0/XI0_50/d__2_ XI11_3/XI0/XI0_50/d_2_ DECAP_INV_G11
XG8984 XI11_3/XI0/XI0_50/d__1_ XI11_3/XI0/XI0_50/d_1_ DECAP_INV_G11
XG8985 XI11_3/XI0/XI0_50/d__0_ XI11_3/XI0/XI0_50/d_0_ DECAP_INV_G11
XG8986 XI11_3/XI0/XI0_50/d_15_ XI11_3/XI0/XI0_50/d__15_ DECAP_INV_G11
XG8987 XI11_3/XI0/XI0_50/d_14_ XI11_3/XI0/XI0_50/d__14_ DECAP_INV_G11
XG8988 XI11_3/XI0/XI0_50/d_13_ XI11_3/XI0/XI0_50/d__13_ DECAP_INV_G11
XG8989 XI11_3/XI0/XI0_50/d_12_ XI11_3/XI0/XI0_50/d__12_ DECAP_INV_G11
XG8990 XI11_3/XI0/XI0_50/d_11_ XI11_3/XI0/XI0_50/d__11_ DECAP_INV_G11
XG8991 XI11_3/XI0/XI0_50/d_10_ XI11_3/XI0/XI0_50/d__10_ DECAP_INV_G11
XG8992 XI11_3/XI0/XI0_50/d_9_ XI11_3/XI0/XI0_50/d__9_ DECAP_INV_G11
XG8993 XI11_3/XI0/XI0_50/d_8_ XI11_3/XI0/XI0_50/d__8_ DECAP_INV_G11
XG8994 XI11_3/XI0/XI0_50/d_7_ XI11_3/XI0/XI0_50/d__7_ DECAP_INV_G11
XG8995 XI11_3/XI0/XI0_50/d_6_ XI11_3/XI0/XI0_50/d__6_ DECAP_INV_G11
XG8996 XI11_3/XI0/XI0_50/d_5_ XI11_3/XI0/XI0_50/d__5_ DECAP_INV_G11
XG8997 XI11_3/XI0/XI0_50/d_4_ XI11_3/XI0/XI0_50/d__4_ DECAP_INV_G11
XG8998 XI11_3/XI0/XI0_50/d_3_ XI11_3/XI0/XI0_50/d__3_ DECAP_INV_G11
XG8999 XI11_3/XI0/XI0_50/d_2_ XI11_3/XI0/XI0_50/d__2_ DECAP_INV_G11
XG9000 XI11_3/XI0/XI0_50/d_1_ XI11_3/XI0/XI0_50/d__1_ DECAP_INV_G11
XG9001 XI11_3/XI0/XI0_50/d_0_ XI11_3/XI0/XI0_50/d__0_ DECAP_INV_G11
XG9002 XI11_3/XI0/XI0_49/d__15_ XI11_3/XI0/XI0_49/d_15_ DECAP_INV_G11
XG9003 XI11_3/XI0/XI0_49/d__14_ XI11_3/XI0/XI0_49/d_14_ DECAP_INV_G11
XG9004 XI11_3/XI0/XI0_49/d__13_ XI11_3/XI0/XI0_49/d_13_ DECAP_INV_G11
XG9005 XI11_3/XI0/XI0_49/d__12_ XI11_3/XI0/XI0_49/d_12_ DECAP_INV_G11
XG9006 XI11_3/XI0/XI0_49/d__11_ XI11_3/XI0/XI0_49/d_11_ DECAP_INV_G11
XG9007 XI11_3/XI0/XI0_49/d__10_ XI11_3/XI0/XI0_49/d_10_ DECAP_INV_G11
XG9008 XI11_3/XI0/XI0_49/d__9_ XI11_3/XI0/XI0_49/d_9_ DECAP_INV_G11
XG9009 XI11_3/XI0/XI0_49/d__8_ XI11_3/XI0/XI0_49/d_8_ DECAP_INV_G11
XG9010 XI11_3/XI0/XI0_49/d__7_ XI11_3/XI0/XI0_49/d_7_ DECAP_INV_G11
XG9011 XI11_3/XI0/XI0_49/d__6_ XI11_3/XI0/XI0_49/d_6_ DECAP_INV_G11
XG9012 XI11_3/XI0/XI0_49/d__5_ XI11_3/XI0/XI0_49/d_5_ DECAP_INV_G11
XG9013 XI11_3/XI0/XI0_49/d__4_ XI11_3/XI0/XI0_49/d_4_ DECAP_INV_G11
XG9014 XI11_3/XI0/XI0_49/d__3_ XI11_3/XI0/XI0_49/d_3_ DECAP_INV_G11
XG9015 XI11_3/XI0/XI0_49/d__2_ XI11_3/XI0/XI0_49/d_2_ DECAP_INV_G11
XG9016 XI11_3/XI0/XI0_49/d__1_ XI11_3/XI0/XI0_49/d_1_ DECAP_INV_G11
XG9017 XI11_3/XI0/XI0_49/d__0_ XI11_3/XI0/XI0_49/d_0_ DECAP_INV_G11
XG9018 XI11_3/XI0/XI0_49/d_15_ XI11_3/XI0/XI0_49/d__15_ DECAP_INV_G11
XG9019 XI11_3/XI0/XI0_49/d_14_ XI11_3/XI0/XI0_49/d__14_ DECAP_INV_G11
XG9020 XI11_3/XI0/XI0_49/d_13_ XI11_3/XI0/XI0_49/d__13_ DECAP_INV_G11
XG9021 XI11_3/XI0/XI0_49/d_12_ XI11_3/XI0/XI0_49/d__12_ DECAP_INV_G11
XG9022 XI11_3/XI0/XI0_49/d_11_ XI11_3/XI0/XI0_49/d__11_ DECAP_INV_G11
XG9023 XI11_3/XI0/XI0_49/d_10_ XI11_3/XI0/XI0_49/d__10_ DECAP_INV_G11
XG9024 XI11_3/XI0/XI0_49/d_9_ XI11_3/XI0/XI0_49/d__9_ DECAP_INV_G11
XG9025 XI11_3/XI0/XI0_49/d_8_ XI11_3/XI0/XI0_49/d__8_ DECAP_INV_G11
XG9026 XI11_3/XI0/XI0_49/d_7_ XI11_3/XI0/XI0_49/d__7_ DECAP_INV_G11
XG9027 XI11_3/XI0/XI0_49/d_6_ XI11_3/XI0/XI0_49/d__6_ DECAP_INV_G11
XG9028 XI11_3/XI0/XI0_49/d_5_ XI11_3/XI0/XI0_49/d__5_ DECAP_INV_G11
XG9029 XI11_3/XI0/XI0_49/d_4_ XI11_3/XI0/XI0_49/d__4_ DECAP_INV_G11
XG9030 XI11_3/XI0/XI0_49/d_3_ XI11_3/XI0/XI0_49/d__3_ DECAP_INV_G11
XG9031 XI11_3/XI0/XI0_49/d_2_ XI11_3/XI0/XI0_49/d__2_ DECAP_INV_G11
XG9032 XI11_3/XI0/XI0_49/d_1_ XI11_3/XI0/XI0_49/d__1_ DECAP_INV_G11
XG9033 XI11_3/XI0/XI0_49/d_0_ XI11_3/XI0/XI0_49/d__0_ DECAP_INV_G11
XG9034 XI11_3/XI0/XI0_48/d__15_ XI11_3/XI0/XI0_48/d_15_ DECAP_INV_G11
XG9035 XI11_3/XI0/XI0_48/d__14_ XI11_3/XI0/XI0_48/d_14_ DECAP_INV_G11
XG9036 XI11_3/XI0/XI0_48/d__13_ XI11_3/XI0/XI0_48/d_13_ DECAP_INV_G11
XG9037 XI11_3/XI0/XI0_48/d__12_ XI11_3/XI0/XI0_48/d_12_ DECAP_INV_G11
XG9038 XI11_3/XI0/XI0_48/d__11_ XI11_3/XI0/XI0_48/d_11_ DECAP_INV_G11
XG9039 XI11_3/XI0/XI0_48/d__10_ XI11_3/XI0/XI0_48/d_10_ DECAP_INV_G11
XG9040 XI11_3/XI0/XI0_48/d__9_ XI11_3/XI0/XI0_48/d_9_ DECAP_INV_G11
XG9041 XI11_3/XI0/XI0_48/d__8_ XI11_3/XI0/XI0_48/d_8_ DECAP_INV_G11
XG9042 XI11_3/XI0/XI0_48/d__7_ XI11_3/XI0/XI0_48/d_7_ DECAP_INV_G11
XG9043 XI11_3/XI0/XI0_48/d__6_ XI11_3/XI0/XI0_48/d_6_ DECAP_INV_G11
XG9044 XI11_3/XI0/XI0_48/d__5_ XI11_3/XI0/XI0_48/d_5_ DECAP_INV_G11
XG9045 XI11_3/XI0/XI0_48/d__4_ XI11_3/XI0/XI0_48/d_4_ DECAP_INV_G11
XG9046 XI11_3/XI0/XI0_48/d__3_ XI11_3/XI0/XI0_48/d_3_ DECAP_INV_G11
XG9047 XI11_3/XI0/XI0_48/d__2_ XI11_3/XI0/XI0_48/d_2_ DECAP_INV_G11
XG9048 XI11_3/XI0/XI0_48/d__1_ XI11_3/XI0/XI0_48/d_1_ DECAP_INV_G11
XG9049 XI11_3/XI0/XI0_48/d__0_ XI11_3/XI0/XI0_48/d_0_ DECAP_INV_G11
XG9050 XI11_3/XI0/XI0_48/d_15_ XI11_3/XI0/XI0_48/d__15_ DECAP_INV_G11
XG9051 XI11_3/XI0/XI0_48/d_14_ XI11_3/XI0/XI0_48/d__14_ DECAP_INV_G11
XG9052 XI11_3/XI0/XI0_48/d_13_ XI11_3/XI0/XI0_48/d__13_ DECAP_INV_G11
XG9053 XI11_3/XI0/XI0_48/d_12_ XI11_3/XI0/XI0_48/d__12_ DECAP_INV_G11
XG9054 XI11_3/XI0/XI0_48/d_11_ XI11_3/XI0/XI0_48/d__11_ DECAP_INV_G11
XG9055 XI11_3/XI0/XI0_48/d_10_ XI11_3/XI0/XI0_48/d__10_ DECAP_INV_G11
XG9056 XI11_3/XI0/XI0_48/d_9_ XI11_3/XI0/XI0_48/d__9_ DECAP_INV_G11
XG9057 XI11_3/XI0/XI0_48/d_8_ XI11_3/XI0/XI0_48/d__8_ DECAP_INV_G11
XG9058 XI11_3/XI0/XI0_48/d_7_ XI11_3/XI0/XI0_48/d__7_ DECAP_INV_G11
XG9059 XI11_3/XI0/XI0_48/d_6_ XI11_3/XI0/XI0_48/d__6_ DECAP_INV_G11
XG9060 XI11_3/XI0/XI0_48/d_5_ XI11_3/XI0/XI0_48/d__5_ DECAP_INV_G11
XG9061 XI11_3/XI0/XI0_48/d_4_ XI11_3/XI0/XI0_48/d__4_ DECAP_INV_G11
XG9062 XI11_3/XI0/XI0_48/d_3_ XI11_3/XI0/XI0_48/d__3_ DECAP_INV_G11
XG9063 XI11_3/XI0/XI0_48/d_2_ XI11_3/XI0/XI0_48/d__2_ DECAP_INV_G11
XG9064 XI11_3/XI0/XI0_48/d_1_ XI11_3/XI0/XI0_48/d__1_ DECAP_INV_G11
XG9065 XI11_3/XI0/XI0_48/d_0_ XI11_3/XI0/XI0_48/d__0_ DECAP_INV_G11
XG9066 XI11_3/XI0/XI0_47/d__15_ XI11_3/XI0/XI0_47/d_15_ DECAP_INV_G11
XG9067 XI11_3/XI0/XI0_47/d__14_ XI11_3/XI0/XI0_47/d_14_ DECAP_INV_G11
XG9068 XI11_3/XI0/XI0_47/d__13_ XI11_3/XI0/XI0_47/d_13_ DECAP_INV_G11
XG9069 XI11_3/XI0/XI0_47/d__12_ XI11_3/XI0/XI0_47/d_12_ DECAP_INV_G11
XG9070 XI11_3/XI0/XI0_47/d__11_ XI11_3/XI0/XI0_47/d_11_ DECAP_INV_G11
XG9071 XI11_3/XI0/XI0_47/d__10_ XI11_3/XI0/XI0_47/d_10_ DECAP_INV_G11
XG9072 XI11_3/XI0/XI0_47/d__9_ XI11_3/XI0/XI0_47/d_9_ DECAP_INV_G11
XG9073 XI11_3/XI0/XI0_47/d__8_ XI11_3/XI0/XI0_47/d_8_ DECAP_INV_G11
XG9074 XI11_3/XI0/XI0_47/d__7_ XI11_3/XI0/XI0_47/d_7_ DECAP_INV_G11
XG9075 XI11_3/XI0/XI0_47/d__6_ XI11_3/XI0/XI0_47/d_6_ DECAP_INV_G11
XG9076 XI11_3/XI0/XI0_47/d__5_ XI11_3/XI0/XI0_47/d_5_ DECAP_INV_G11
XG9077 XI11_3/XI0/XI0_47/d__4_ XI11_3/XI0/XI0_47/d_4_ DECAP_INV_G11
XG9078 XI11_3/XI0/XI0_47/d__3_ XI11_3/XI0/XI0_47/d_3_ DECAP_INV_G11
XG9079 XI11_3/XI0/XI0_47/d__2_ XI11_3/XI0/XI0_47/d_2_ DECAP_INV_G11
XG9080 XI11_3/XI0/XI0_47/d__1_ XI11_3/XI0/XI0_47/d_1_ DECAP_INV_G11
XG9081 XI11_3/XI0/XI0_47/d__0_ XI11_3/XI0/XI0_47/d_0_ DECAP_INV_G11
XG9082 XI11_3/XI0/XI0_47/d_15_ XI11_3/XI0/XI0_47/d__15_ DECAP_INV_G11
XG9083 XI11_3/XI0/XI0_47/d_14_ XI11_3/XI0/XI0_47/d__14_ DECAP_INV_G11
XG9084 XI11_3/XI0/XI0_47/d_13_ XI11_3/XI0/XI0_47/d__13_ DECAP_INV_G11
XG9085 XI11_3/XI0/XI0_47/d_12_ XI11_3/XI0/XI0_47/d__12_ DECAP_INV_G11
XG9086 XI11_3/XI0/XI0_47/d_11_ XI11_3/XI0/XI0_47/d__11_ DECAP_INV_G11
XG9087 XI11_3/XI0/XI0_47/d_10_ XI11_3/XI0/XI0_47/d__10_ DECAP_INV_G11
XG9088 XI11_3/XI0/XI0_47/d_9_ XI11_3/XI0/XI0_47/d__9_ DECAP_INV_G11
XG9089 XI11_3/XI0/XI0_47/d_8_ XI11_3/XI0/XI0_47/d__8_ DECAP_INV_G11
XG9090 XI11_3/XI0/XI0_47/d_7_ XI11_3/XI0/XI0_47/d__7_ DECAP_INV_G11
XG9091 XI11_3/XI0/XI0_47/d_6_ XI11_3/XI0/XI0_47/d__6_ DECAP_INV_G11
XG9092 XI11_3/XI0/XI0_47/d_5_ XI11_3/XI0/XI0_47/d__5_ DECAP_INV_G11
XG9093 XI11_3/XI0/XI0_47/d_4_ XI11_3/XI0/XI0_47/d__4_ DECAP_INV_G11
XG9094 XI11_3/XI0/XI0_47/d_3_ XI11_3/XI0/XI0_47/d__3_ DECAP_INV_G11
XG9095 XI11_3/XI0/XI0_47/d_2_ XI11_3/XI0/XI0_47/d__2_ DECAP_INV_G11
XG9096 XI11_3/XI0/XI0_47/d_1_ XI11_3/XI0/XI0_47/d__1_ DECAP_INV_G11
XG9097 XI11_3/XI0/XI0_47/d_0_ XI11_3/XI0/XI0_47/d__0_ DECAP_INV_G11
XG9098 XI11_3/XI0/XI0_46/d__15_ XI11_3/XI0/XI0_46/d_15_ DECAP_INV_G11
XG9099 XI11_3/XI0/XI0_46/d__14_ XI11_3/XI0/XI0_46/d_14_ DECAP_INV_G11
XG9100 XI11_3/XI0/XI0_46/d__13_ XI11_3/XI0/XI0_46/d_13_ DECAP_INV_G11
XG9101 XI11_3/XI0/XI0_46/d__12_ XI11_3/XI0/XI0_46/d_12_ DECAP_INV_G11
XG9102 XI11_3/XI0/XI0_46/d__11_ XI11_3/XI0/XI0_46/d_11_ DECAP_INV_G11
XG9103 XI11_3/XI0/XI0_46/d__10_ XI11_3/XI0/XI0_46/d_10_ DECAP_INV_G11
XG9104 XI11_3/XI0/XI0_46/d__9_ XI11_3/XI0/XI0_46/d_9_ DECAP_INV_G11
XG9105 XI11_3/XI0/XI0_46/d__8_ XI11_3/XI0/XI0_46/d_8_ DECAP_INV_G11
XG9106 XI11_3/XI0/XI0_46/d__7_ XI11_3/XI0/XI0_46/d_7_ DECAP_INV_G11
XG9107 XI11_3/XI0/XI0_46/d__6_ XI11_3/XI0/XI0_46/d_6_ DECAP_INV_G11
XG9108 XI11_3/XI0/XI0_46/d__5_ XI11_3/XI0/XI0_46/d_5_ DECAP_INV_G11
XG9109 XI11_3/XI0/XI0_46/d__4_ XI11_3/XI0/XI0_46/d_4_ DECAP_INV_G11
XG9110 XI11_3/XI0/XI0_46/d__3_ XI11_3/XI0/XI0_46/d_3_ DECAP_INV_G11
XG9111 XI11_3/XI0/XI0_46/d__2_ XI11_3/XI0/XI0_46/d_2_ DECAP_INV_G11
XG9112 XI11_3/XI0/XI0_46/d__1_ XI11_3/XI0/XI0_46/d_1_ DECAP_INV_G11
XG9113 XI11_3/XI0/XI0_46/d__0_ XI11_3/XI0/XI0_46/d_0_ DECAP_INV_G11
XG9114 XI11_3/XI0/XI0_46/d_15_ XI11_3/XI0/XI0_46/d__15_ DECAP_INV_G11
XG9115 XI11_3/XI0/XI0_46/d_14_ XI11_3/XI0/XI0_46/d__14_ DECAP_INV_G11
XG9116 XI11_3/XI0/XI0_46/d_13_ XI11_3/XI0/XI0_46/d__13_ DECAP_INV_G11
XG9117 XI11_3/XI0/XI0_46/d_12_ XI11_3/XI0/XI0_46/d__12_ DECAP_INV_G11
XG9118 XI11_3/XI0/XI0_46/d_11_ XI11_3/XI0/XI0_46/d__11_ DECAP_INV_G11
XG9119 XI11_3/XI0/XI0_46/d_10_ XI11_3/XI0/XI0_46/d__10_ DECAP_INV_G11
XG9120 XI11_3/XI0/XI0_46/d_9_ XI11_3/XI0/XI0_46/d__9_ DECAP_INV_G11
XG9121 XI11_3/XI0/XI0_46/d_8_ XI11_3/XI0/XI0_46/d__8_ DECAP_INV_G11
XG9122 XI11_3/XI0/XI0_46/d_7_ XI11_3/XI0/XI0_46/d__7_ DECAP_INV_G11
XG9123 XI11_3/XI0/XI0_46/d_6_ XI11_3/XI0/XI0_46/d__6_ DECAP_INV_G11
XG9124 XI11_3/XI0/XI0_46/d_5_ XI11_3/XI0/XI0_46/d__5_ DECAP_INV_G11
XG9125 XI11_3/XI0/XI0_46/d_4_ XI11_3/XI0/XI0_46/d__4_ DECAP_INV_G11
XG9126 XI11_3/XI0/XI0_46/d_3_ XI11_3/XI0/XI0_46/d__3_ DECAP_INV_G11
XG9127 XI11_3/XI0/XI0_46/d_2_ XI11_3/XI0/XI0_46/d__2_ DECAP_INV_G11
XG9128 XI11_3/XI0/XI0_46/d_1_ XI11_3/XI0/XI0_46/d__1_ DECAP_INV_G11
XG9129 XI11_3/XI0/XI0_46/d_0_ XI11_3/XI0/XI0_46/d__0_ DECAP_INV_G11
XG9130 XI11_3/XI0/XI0_45/d__15_ XI11_3/XI0/XI0_45/d_15_ DECAP_INV_G11
XG9131 XI11_3/XI0/XI0_45/d__14_ XI11_3/XI0/XI0_45/d_14_ DECAP_INV_G11
XG9132 XI11_3/XI0/XI0_45/d__13_ XI11_3/XI0/XI0_45/d_13_ DECAP_INV_G11
XG9133 XI11_3/XI0/XI0_45/d__12_ XI11_3/XI0/XI0_45/d_12_ DECAP_INV_G11
XG9134 XI11_3/XI0/XI0_45/d__11_ XI11_3/XI0/XI0_45/d_11_ DECAP_INV_G11
XG9135 XI11_3/XI0/XI0_45/d__10_ XI11_3/XI0/XI0_45/d_10_ DECAP_INV_G11
XG9136 XI11_3/XI0/XI0_45/d__9_ XI11_3/XI0/XI0_45/d_9_ DECAP_INV_G11
XG9137 XI11_3/XI0/XI0_45/d__8_ XI11_3/XI0/XI0_45/d_8_ DECAP_INV_G11
XG9138 XI11_3/XI0/XI0_45/d__7_ XI11_3/XI0/XI0_45/d_7_ DECAP_INV_G11
XG9139 XI11_3/XI0/XI0_45/d__6_ XI11_3/XI0/XI0_45/d_6_ DECAP_INV_G11
XG9140 XI11_3/XI0/XI0_45/d__5_ XI11_3/XI0/XI0_45/d_5_ DECAP_INV_G11
XG9141 XI11_3/XI0/XI0_45/d__4_ XI11_3/XI0/XI0_45/d_4_ DECAP_INV_G11
XG9142 XI11_3/XI0/XI0_45/d__3_ XI11_3/XI0/XI0_45/d_3_ DECAP_INV_G11
XG9143 XI11_3/XI0/XI0_45/d__2_ XI11_3/XI0/XI0_45/d_2_ DECAP_INV_G11
XG9144 XI11_3/XI0/XI0_45/d__1_ XI11_3/XI0/XI0_45/d_1_ DECAP_INV_G11
XG9145 XI11_3/XI0/XI0_45/d__0_ XI11_3/XI0/XI0_45/d_0_ DECAP_INV_G11
XG9146 XI11_3/XI0/XI0_45/d_15_ XI11_3/XI0/XI0_45/d__15_ DECAP_INV_G11
XG9147 XI11_3/XI0/XI0_45/d_14_ XI11_3/XI0/XI0_45/d__14_ DECAP_INV_G11
XG9148 XI11_3/XI0/XI0_45/d_13_ XI11_3/XI0/XI0_45/d__13_ DECAP_INV_G11
XG9149 XI11_3/XI0/XI0_45/d_12_ XI11_3/XI0/XI0_45/d__12_ DECAP_INV_G11
XG9150 XI11_3/XI0/XI0_45/d_11_ XI11_3/XI0/XI0_45/d__11_ DECAP_INV_G11
XG9151 XI11_3/XI0/XI0_45/d_10_ XI11_3/XI0/XI0_45/d__10_ DECAP_INV_G11
XG9152 XI11_3/XI0/XI0_45/d_9_ XI11_3/XI0/XI0_45/d__9_ DECAP_INV_G11
XG9153 XI11_3/XI0/XI0_45/d_8_ XI11_3/XI0/XI0_45/d__8_ DECAP_INV_G11
XG9154 XI11_3/XI0/XI0_45/d_7_ XI11_3/XI0/XI0_45/d__7_ DECAP_INV_G11
XG9155 XI11_3/XI0/XI0_45/d_6_ XI11_3/XI0/XI0_45/d__6_ DECAP_INV_G11
XG9156 XI11_3/XI0/XI0_45/d_5_ XI11_3/XI0/XI0_45/d__5_ DECAP_INV_G11
XG9157 XI11_3/XI0/XI0_45/d_4_ XI11_3/XI0/XI0_45/d__4_ DECAP_INV_G11
XG9158 XI11_3/XI0/XI0_45/d_3_ XI11_3/XI0/XI0_45/d__3_ DECAP_INV_G11
XG9159 XI11_3/XI0/XI0_45/d_2_ XI11_3/XI0/XI0_45/d__2_ DECAP_INV_G11
XG9160 XI11_3/XI0/XI0_45/d_1_ XI11_3/XI0/XI0_45/d__1_ DECAP_INV_G11
XG9161 XI11_3/XI0/XI0_45/d_0_ XI11_3/XI0/XI0_45/d__0_ DECAP_INV_G11
XG9162 XI11_3/XI0/XI0_44/d__15_ XI11_3/XI0/XI0_44/d_15_ DECAP_INV_G11
XG9163 XI11_3/XI0/XI0_44/d__14_ XI11_3/XI0/XI0_44/d_14_ DECAP_INV_G11
XG9164 XI11_3/XI0/XI0_44/d__13_ XI11_3/XI0/XI0_44/d_13_ DECAP_INV_G11
XG9165 XI11_3/XI0/XI0_44/d__12_ XI11_3/XI0/XI0_44/d_12_ DECAP_INV_G11
XG9166 XI11_3/XI0/XI0_44/d__11_ XI11_3/XI0/XI0_44/d_11_ DECAP_INV_G11
XG9167 XI11_3/XI0/XI0_44/d__10_ XI11_3/XI0/XI0_44/d_10_ DECAP_INV_G11
XG9168 XI11_3/XI0/XI0_44/d__9_ XI11_3/XI0/XI0_44/d_9_ DECAP_INV_G11
XG9169 XI11_3/XI0/XI0_44/d__8_ XI11_3/XI0/XI0_44/d_8_ DECAP_INV_G11
XG9170 XI11_3/XI0/XI0_44/d__7_ XI11_3/XI0/XI0_44/d_7_ DECAP_INV_G11
XG9171 XI11_3/XI0/XI0_44/d__6_ XI11_3/XI0/XI0_44/d_6_ DECAP_INV_G11
XG9172 XI11_3/XI0/XI0_44/d__5_ XI11_3/XI0/XI0_44/d_5_ DECAP_INV_G11
XG9173 XI11_3/XI0/XI0_44/d__4_ XI11_3/XI0/XI0_44/d_4_ DECAP_INV_G11
XG9174 XI11_3/XI0/XI0_44/d__3_ XI11_3/XI0/XI0_44/d_3_ DECAP_INV_G11
XG9175 XI11_3/XI0/XI0_44/d__2_ XI11_3/XI0/XI0_44/d_2_ DECAP_INV_G11
XG9176 XI11_3/XI0/XI0_44/d__1_ XI11_3/XI0/XI0_44/d_1_ DECAP_INV_G11
XG9177 XI11_3/XI0/XI0_44/d__0_ XI11_3/XI0/XI0_44/d_0_ DECAP_INV_G11
XG9178 XI11_3/XI0/XI0_44/d_15_ XI11_3/XI0/XI0_44/d__15_ DECAP_INV_G11
XG9179 XI11_3/XI0/XI0_44/d_14_ XI11_3/XI0/XI0_44/d__14_ DECAP_INV_G11
XG9180 XI11_3/XI0/XI0_44/d_13_ XI11_3/XI0/XI0_44/d__13_ DECAP_INV_G11
XG9181 XI11_3/XI0/XI0_44/d_12_ XI11_3/XI0/XI0_44/d__12_ DECAP_INV_G11
XG9182 XI11_3/XI0/XI0_44/d_11_ XI11_3/XI0/XI0_44/d__11_ DECAP_INV_G11
XG9183 XI11_3/XI0/XI0_44/d_10_ XI11_3/XI0/XI0_44/d__10_ DECAP_INV_G11
XG9184 XI11_3/XI0/XI0_44/d_9_ XI11_3/XI0/XI0_44/d__9_ DECAP_INV_G11
XG9185 XI11_3/XI0/XI0_44/d_8_ XI11_3/XI0/XI0_44/d__8_ DECAP_INV_G11
XG9186 XI11_3/XI0/XI0_44/d_7_ XI11_3/XI0/XI0_44/d__7_ DECAP_INV_G11
XG9187 XI11_3/XI0/XI0_44/d_6_ XI11_3/XI0/XI0_44/d__6_ DECAP_INV_G11
XG9188 XI11_3/XI0/XI0_44/d_5_ XI11_3/XI0/XI0_44/d__5_ DECAP_INV_G11
XG9189 XI11_3/XI0/XI0_44/d_4_ XI11_3/XI0/XI0_44/d__4_ DECAP_INV_G11
XG9190 XI11_3/XI0/XI0_44/d_3_ XI11_3/XI0/XI0_44/d__3_ DECAP_INV_G11
XG9191 XI11_3/XI0/XI0_44/d_2_ XI11_3/XI0/XI0_44/d__2_ DECAP_INV_G11
XG9192 XI11_3/XI0/XI0_44/d_1_ XI11_3/XI0/XI0_44/d__1_ DECAP_INV_G11
XG9193 XI11_3/XI0/XI0_44/d_0_ XI11_3/XI0/XI0_44/d__0_ DECAP_INV_G11
XG9194 XI11_3/XI0/XI0_43/d__15_ XI11_3/XI0/XI0_43/d_15_ DECAP_INV_G11
XG9195 XI11_3/XI0/XI0_43/d__14_ XI11_3/XI0/XI0_43/d_14_ DECAP_INV_G11
XG9196 XI11_3/XI0/XI0_43/d__13_ XI11_3/XI0/XI0_43/d_13_ DECAP_INV_G11
XG9197 XI11_3/XI0/XI0_43/d__12_ XI11_3/XI0/XI0_43/d_12_ DECAP_INV_G11
XG9198 XI11_3/XI0/XI0_43/d__11_ XI11_3/XI0/XI0_43/d_11_ DECAP_INV_G11
XG9199 XI11_3/XI0/XI0_43/d__10_ XI11_3/XI0/XI0_43/d_10_ DECAP_INV_G11
XG9200 XI11_3/XI0/XI0_43/d__9_ XI11_3/XI0/XI0_43/d_9_ DECAP_INV_G11
XG9201 XI11_3/XI0/XI0_43/d__8_ XI11_3/XI0/XI0_43/d_8_ DECAP_INV_G11
XG9202 XI11_3/XI0/XI0_43/d__7_ XI11_3/XI0/XI0_43/d_7_ DECAP_INV_G11
XG9203 XI11_3/XI0/XI0_43/d__6_ XI11_3/XI0/XI0_43/d_6_ DECAP_INV_G11
XG9204 XI11_3/XI0/XI0_43/d__5_ XI11_3/XI0/XI0_43/d_5_ DECAP_INV_G11
XG9205 XI11_3/XI0/XI0_43/d__4_ XI11_3/XI0/XI0_43/d_4_ DECAP_INV_G11
XG9206 XI11_3/XI0/XI0_43/d__3_ XI11_3/XI0/XI0_43/d_3_ DECAP_INV_G11
XG9207 XI11_3/XI0/XI0_43/d__2_ XI11_3/XI0/XI0_43/d_2_ DECAP_INV_G11
XG9208 XI11_3/XI0/XI0_43/d__1_ XI11_3/XI0/XI0_43/d_1_ DECAP_INV_G11
XG9209 XI11_3/XI0/XI0_43/d__0_ XI11_3/XI0/XI0_43/d_0_ DECAP_INV_G11
XG9210 XI11_3/XI0/XI0_43/d_15_ XI11_3/XI0/XI0_43/d__15_ DECAP_INV_G11
XG9211 XI11_3/XI0/XI0_43/d_14_ XI11_3/XI0/XI0_43/d__14_ DECAP_INV_G11
XG9212 XI11_3/XI0/XI0_43/d_13_ XI11_3/XI0/XI0_43/d__13_ DECAP_INV_G11
XG9213 XI11_3/XI0/XI0_43/d_12_ XI11_3/XI0/XI0_43/d__12_ DECAP_INV_G11
XG9214 XI11_3/XI0/XI0_43/d_11_ XI11_3/XI0/XI0_43/d__11_ DECAP_INV_G11
XG9215 XI11_3/XI0/XI0_43/d_10_ XI11_3/XI0/XI0_43/d__10_ DECAP_INV_G11
XG9216 XI11_3/XI0/XI0_43/d_9_ XI11_3/XI0/XI0_43/d__9_ DECAP_INV_G11
XG9217 XI11_3/XI0/XI0_43/d_8_ XI11_3/XI0/XI0_43/d__8_ DECAP_INV_G11
XG9218 XI11_3/XI0/XI0_43/d_7_ XI11_3/XI0/XI0_43/d__7_ DECAP_INV_G11
XG9219 XI11_3/XI0/XI0_43/d_6_ XI11_3/XI0/XI0_43/d__6_ DECAP_INV_G11
XG9220 XI11_3/XI0/XI0_43/d_5_ XI11_3/XI0/XI0_43/d__5_ DECAP_INV_G11
XG9221 XI11_3/XI0/XI0_43/d_4_ XI11_3/XI0/XI0_43/d__4_ DECAP_INV_G11
XG9222 XI11_3/XI0/XI0_43/d_3_ XI11_3/XI0/XI0_43/d__3_ DECAP_INV_G11
XG9223 XI11_3/XI0/XI0_43/d_2_ XI11_3/XI0/XI0_43/d__2_ DECAP_INV_G11
XG9224 XI11_3/XI0/XI0_43/d_1_ XI11_3/XI0/XI0_43/d__1_ DECAP_INV_G11
XG9225 XI11_3/XI0/XI0_43/d_0_ XI11_3/XI0/XI0_43/d__0_ DECAP_INV_G11
XG9226 XI11_3/XI0/XI0_42/d__15_ XI11_3/XI0/XI0_42/d_15_ DECAP_INV_G11
XG9227 XI11_3/XI0/XI0_42/d__14_ XI11_3/XI0/XI0_42/d_14_ DECAP_INV_G11
XG9228 XI11_3/XI0/XI0_42/d__13_ XI11_3/XI0/XI0_42/d_13_ DECAP_INV_G11
XG9229 XI11_3/XI0/XI0_42/d__12_ XI11_3/XI0/XI0_42/d_12_ DECAP_INV_G11
XG9230 XI11_3/XI0/XI0_42/d__11_ XI11_3/XI0/XI0_42/d_11_ DECAP_INV_G11
XG9231 XI11_3/XI0/XI0_42/d__10_ XI11_3/XI0/XI0_42/d_10_ DECAP_INV_G11
XG9232 XI11_3/XI0/XI0_42/d__9_ XI11_3/XI0/XI0_42/d_9_ DECAP_INV_G11
XG9233 XI11_3/XI0/XI0_42/d__8_ XI11_3/XI0/XI0_42/d_8_ DECAP_INV_G11
XG9234 XI11_3/XI0/XI0_42/d__7_ XI11_3/XI0/XI0_42/d_7_ DECAP_INV_G11
XG9235 XI11_3/XI0/XI0_42/d__6_ XI11_3/XI0/XI0_42/d_6_ DECAP_INV_G11
XG9236 XI11_3/XI0/XI0_42/d__5_ XI11_3/XI0/XI0_42/d_5_ DECAP_INV_G11
XG9237 XI11_3/XI0/XI0_42/d__4_ XI11_3/XI0/XI0_42/d_4_ DECAP_INV_G11
XG9238 XI11_3/XI0/XI0_42/d__3_ XI11_3/XI0/XI0_42/d_3_ DECAP_INV_G11
XG9239 XI11_3/XI0/XI0_42/d__2_ XI11_3/XI0/XI0_42/d_2_ DECAP_INV_G11
XG9240 XI11_3/XI0/XI0_42/d__1_ XI11_3/XI0/XI0_42/d_1_ DECAP_INV_G11
XG9241 XI11_3/XI0/XI0_42/d__0_ XI11_3/XI0/XI0_42/d_0_ DECAP_INV_G11
XG9242 XI11_3/XI0/XI0_42/d_15_ XI11_3/XI0/XI0_42/d__15_ DECAP_INV_G11
XG9243 XI11_3/XI0/XI0_42/d_14_ XI11_3/XI0/XI0_42/d__14_ DECAP_INV_G11
XG9244 XI11_3/XI0/XI0_42/d_13_ XI11_3/XI0/XI0_42/d__13_ DECAP_INV_G11
XG9245 XI11_3/XI0/XI0_42/d_12_ XI11_3/XI0/XI0_42/d__12_ DECAP_INV_G11
XG9246 XI11_3/XI0/XI0_42/d_11_ XI11_3/XI0/XI0_42/d__11_ DECAP_INV_G11
XG9247 XI11_3/XI0/XI0_42/d_10_ XI11_3/XI0/XI0_42/d__10_ DECAP_INV_G11
XG9248 XI11_3/XI0/XI0_42/d_9_ XI11_3/XI0/XI0_42/d__9_ DECAP_INV_G11
XG9249 XI11_3/XI0/XI0_42/d_8_ XI11_3/XI0/XI0_42/d__8_ DECAP_INV_G11
XG9250 XI11_3/XI0/XI0_42/d_7_ XI11_3/XI0/XI0_42/d__7_ DECAP_INV_G11
XG9251 XI11_3/XI0/XI0_42/d_6_ XI11_3/XI0/XI0_42/d__6_ DECAP_INV_G11
XG9252 XI11_3/XI0/XI0_42/d_5_ XI11_3/XI0/XI0_42/d__5_ DECAP_INV_G11
XG9253 XI11_3/XI0/XI0_42/d_4_ XI11_3/XI0/XI0_42/d__4_ DECAP_INV_G11
XG9254 XI11_3/XI0/XI0_42/d_3_ XI11_3/XI0/XI0_42/d__3_ DECAP_INV_G11
XG9255 XI11_3/XI0/XI0_42/d_2_ XI11_3/XI0/XI0_42/d__2_ DECAP_INV_G11
XG9256 XI11_3/XI0/XI0_42/d_1_ XI11_3/XI0/XI0_42/d__1_ DECAP_INV_G11
XG9257 XI11_3/XI0/XI0_42/d_0_ XI11_3/XI0/XI0_42/d__0_ DECAP_INV_G11
XG9258 XI11_3/XI0/XI0_41/d__15_ XI11_3/XI0/XI0_41/d_15_ DECAP_INV_G11
XG9259 XI11_3/XI0/XI0_41/d__14_ XI11_3/XI0/XI0_41/d_14_ DECAP_INV_G11
XG9260 XI11_3/XI0/XI0_41/d__13_ XI11_3/XI0/XI0_41/d_13_ DECAP_INV_G11
XG9261 XI11_3/XI0/XI0_41/d__12_ XI11_3/XI0/XI0_41/d_12_ DECAP_INV_G11
XG9262 XI11_3/XI0/XI0_41/d__11_ XI11_3/XI0/XI0_41/d_11_ DECAP_INV_G11
XG9263 XI11_3/XI0/XI0_41/d__10_ XI11_3/XI0/XI0_41/d_10_ DECAP_INV_G11
XG9264 XI11_3/XI0/XI0_41/d__9_ XI11_3/XI0/XI0_41/d_9_ DECAP_INV_G11
XG9265 XI11_3/XI0/XI0_41/d__8_ XI11_3/XI0/XI0_41/d_8_ DECAP_INV_G11
XG9266 XI11_3/XI0/XI0_41/d__7_ XI11_3/XI0/XI0_41/d_7_ DECAP_INV_G11
XG9267 XI11_3/XI0/XI0_41/d__6_ XI11_3/XI0/XI0_41/d_6_ DECAP_INV_G11
XG9268 XI11_3/XI0/XI0_41/d__5_ XI11_3/XI0/XI0_41/d_5_ DECAP_INV_G11
XG9269 XI11_3/XI0/XI0_41/d__4_ XI11_3/XI0/XI0_41/d_4_ DECAP_INV_G11
XG9270 XI11_3/XI0/XI0_41/d__3_ XI11_3/XI0/XI0_41/d_3_ DECAP_INV_G11
XG9271 XI11_3/XI0/XI0_41/d__2_ XI11_3/XI0/XI0_41/d_2_ DECAP_INV_G11
XG9272 XI11_3/XI0/XI0_41/d__1_ XI11_3/XI0/XI0_41/d_1_ DECAP_INV_G11
XG9273 XI11_3/XI0/XI0_41/d__0_ XI11_3/XI0/XI0_41/d_0_ DECAP_INV_G11
XG9274 XI11_3/XI0/XI0_41/d_15_ XI11_3/XI0/XI0_41/d__15_ DECAP_INV_G11
XG9275 XI11_3/XI0/XI0_41/d_14_ XI11_3/XI0/XI0_41/d__14_ DECAP_INV_G11
XG9276 XI11_3/XI0/XI0_41/d_13_ XI11_3/XI0/XI0_41/d__13_ DECAP_INV_G11
XG9277 XI11_3/XI0/XI0_41/d_12_ XI11_3/XI0/XI0_41/d__12_ DECAP_INV_G11
XG9278 XI11_3/XI0/XI0_41/d_11_ XI11_3/XI0/XI0_41/d__11_ DECAP_INV_G11
XG9279 XI11_3/XI0/XI0_41/d_10_ XI11_3/XI0/XI0_41/d__10_ DECAP_INV_G11
XG9280 XI11_3/XI0/XI0_41/d_9_ XI11_3/XI0/XI0_41/d__9_ DECAP_INV_G11
XG9281 XI11_3/XI0/XI0_41/d_8_ XI11_3/XI0/XI0_41/d__8_ DECAP_INV_G11
XG9282 XI11_3/XI0/XI0_41/d_7_ XI11_3/XI0/XI0_41/d__7_ DECAP_INV_G11
XG9283 XI11_3/XI0/XI0_41/d_6_ XI11_3/XI0/XI0_41/d__6_ DECAP_INV_G11
XG9284 XI11_3/XI0/XI0_41/d_5_ XI11_3/XI0/XI0_41/d__5_ DECAP_INV_G11
XG9285 XI11_3/XI0/XI0_41/d_4_ XI11_3/XI0/XI0_41/d__4_ DECAP_INV_G11
XG9286 XI11_3/XI0/XI0_41/d_3_ XI11_3/XI0/XI0_41/d__3_ DECAP_INV_G11
XG9287 XI11_3/XI0/XI0_41/d_2_ XI11_3/XI0/XI0_41/d__2_ DECAP_INV_G11
XG9288 XI11_3/XI0/XI0_41/d_1_ XI11_3/XI0/XI0_41/d__1_ DECAP_INV_G11
XG9289 XI11_3/XI0/XI0_41/d_0_ XI11_3/XI0/XI0_41/d__0_ DECAP_INV_G11
XG9290 XI11_3/XI0/XI0_40/d__15_ XI11_3/XI0/XI0_40/d_15_ DECAP_INV_G11
XG9291 XI11_3/XI0/XI0_40/d__14_ XI11_3/XI0/XI0_40/d_14_ DECAP_INV_G11
XG9292 XI11_3/XI0/XI0_40/d__13_ XI11_3/XI0/XI0_40/d_13_ DECAP_INV_G11
XG9293 XI11_3/XI0/XI0_40/d__12_ XI11_3/XI0/XI0_40/d_12_ DECAP_INV_G11
XG9294 XI11_3/XI0/XI0_40/d__11_ XI11_3/XI0/XI0_40/d_11_ DECAP_INV_G11
XG9295 XI11_3/XI0/XI0_40/d__10_ XI11_3/XI0/XI0_40/d_10_ DECAP_INV_G11
XG9296 XI11_3/XI0/XI0_40/d__9_ XI11_3/XI0/XI0_40/d_9_ DECAP_INV_G11
XG9297 XI11_3/XI0/XI0_40/d__8_ XI11_3/XI0/XI0_40/d_8_ DECAP_INV_G11
XG9298 XI11_3/XI0/XI0_40/d__7_ XI11_3/XI0/XI0_40/d_7_ DECAP_INV_G11
XG9299 XI11_3/XI0/XI0_40/d__6_ XI11_3/XI0/XI0_40/d_6_ DECAP_INV_G11
XG9300 XI11_3/XI0/XI0_40/d__5_ XI11_3/XI0/XI0_40/d_5_ DECAP_INV_G11
XG9301 XI11_3/XI0/XI0_40/d__4_ XI11_3/XI0/XI0_40/d_4_ DECAP_INV_G11
XG9302 XI11_3/XI0/XI0_40/d__3_ XI11_3/XI0/XI0_40/d_3_ DECAP_INV_G11
XG9303 XI11_3/XI0/XI0_40/d__2_ XI11_3/XI0/XI0_40/d_2_ DECAP_INV_G11
XG9304 XI11_3/XI0/XI0_40/d__1_ XI11_3/XI0/XI0_40/d_1_ DECAP_INV_G11
XG9305 XI11_3/XI0/XI0_40/d__0_ XI11_3/XI0/XI0_40/d_0_ DECAP_INV_G11
XG9306 XI11_3/XI0/XI0_40/d_15_ XI11_3/XI0/XI0_40/d__15_ DECAP_INV_G11
XG9307 XI11_3/XI0/XI0_40/d_14_ XI11_3/XI0/XI0_40/d__14_ DECAP_INV_G11
XG9308 XI11_3/XI0/XI0_40/d_13_ XI11_3/XI0/XI0_40/d__13_ DECAP_INV_G11
XG9309 XI11_3/XI0/XI0_40/d_12_ XI11_3/XI0/XI0_40/d__12_ DECAP_INV_G11
XG9310 XI11_3/XI0/XI0_40/d_11_ XI11_3/XI0/XI0_40/d__11_ DECAP_INV_G11
XG9311 XI11_3/XI0/XI0_40/d_10_ XI11_3/XI0/XI0_40/d__10_ DECAP_INV_G11
XG9312 XI11_3/XI0/XI0_40/d_9_ XI11_3/XI0/XI0_40/d__9_ DECAP_INV_G11
XG9313 XI11_3/XI0/XI0_40/d_8_ XI11_3/XI0/XI0_40/d__8_ DECAP_INV_G11
XG9314 XI11_3/XI0/XI0_40/d_7_ XI11_3/XI0/XI0_40/d__7_ DECAP_INV_G11
XG9315 XI11_3/XI0/XI0_40/d_6_ XI11_3/XI0/XI0_40/d__6_ DECAP_INV_G11
XG9316 XI11_3/XI0/XI0_40/d_5_ XI11_3/XI0/XI0_40/d__5_ DECAP_INV_G11
XG9317 XI11_3/XI0/XI0_40/d_4_ XI11_3/XI0/XI0_40/d__4_ DECAP_INV_G11
XG9318 XI11_3/XI0/XI0_40/d_3_ XI11_3/XI0/XI0_40/d__3_ DECAP_INV_G11
XG9319 XI11_3/XI0/XI0_40/d_2_ XI11_3/XI0/XI0_40/d__2_ DECAP_INV_G11
XG9320 XI11_3/XI0/XI0_40/d_1_ XI11_3/XI0/XI0_40/d__1_ DECAP_INV_G11
XG9321 XI11_3/XI0/XI0_40/d_0_ XI11_3/XI0/XI0_40/d__0_ DECAP_INV_G11
XG9322 XI11_3/XI0/XI0_39/d__15_ XI11_3/XI0/XI0_39/d_15_ DECAP_INV_G11
XG9323 XI11_3/XI0/XI0_39/d__14_ XI11_3/XI0/XI0_39/d_14_ DECAP_INV_G11
XG9324 XI11_3/XI0/XI0_39/d__13_ XI11_3/XI0/XI0_39/d_13_ DECAP_INV_G11
XG9325 XI11_3/XI0/XI0_39/d__12_ XI11_3/XI0/XI0_39/d_12_ DECAP_INV_G11
XG9326 XI11_3/XI0/XI0_39/d__11_ XI11_3/XI0/XI0_39/d_11_ DECAP_INV_G11
XG9327 XI11_3/XI0/XI0_39/d__10_ XI11_3/XI0/XI0_39/d_10_ DECAP_INV_G11
XG9328 XI11_3/XI0/XI0_39/d__9_ XI11_3/XI0/XI0_39/d_9_ DECAP_INV_G11
XG9329 XI11_3/XI0/XI0_39/d__8_ XI11_3/XI0/XI0_39/d_8_ DECAP_INV_G11
XG9330 XI11_3/XI0/XI0_39/d__7_ XI11_3/XI0/XI0_39/d_7_ DECAP_INV_G11
XG9331 XI11_3/XI0/XI0_39/d__6_ XI11_3/XI0/XI0_39/d_6_ DECAP_INV_G11
XG9332 XI11_3/XI0/XI0_39/d__5_ XI11_3/XI0/XI0_39/d_5_ DECAP_INV_G11
XG9333 XI11_3/XI0/XI0_39/d__4_ XI11_3/XI0/XI0_39/d_4_ DECAP_INV_G11
XG9334 XI11_3/XI0/XI0_39/d__3_ XI11_3/XI0/XI0_39/d_3_ DECAP_INV_G11
XG9335 XI11_3/XI0/XI0_39/d__2_ XI11_3/XI0/XI0_39/d_2_ DECAP_INV_G11
XG9336 XI11_3/XI0/XI0_39/d__1_ XI11_3/XI0/XI0_39/d_1_ DECAP_INV_G11
XG9337 XI11_3/XI0/XI0_39/d__0_ XI11_3/XI0/XI0_39/d_0_ DECAP_INV_G11
XG9338 XI11_3/XI0/XI0_39/d_15_ XI11_3/XI0/XI0_39/d__15_ DECAP_INV_G11
XG9339 XI11_3/XI0/XI0_39/d_14_ XI11_3/XI0/XI0_39/d__14_ DECAP_INV_G11
XG9340 XI11_3/XI0/XI0_39/d_13_ XI11_3/XI0/XI0_39/d__13_ DECAP_INV_G11
XG9341 XI11_3/XI0/XI0_39/d_12_ XI11_3/XI0/XI0_39/d__12_ DECAP_INV_G11
XG9342 XI11_3/XI0/XI0_39/d_11_ XI11_3/XI0/XI0_39/d__11_ DECAP_INV_G11
XG9343 XI11_3/XI0/XI0_39/d_10_ XI11_3/XI0/XI0_39/d__10_ DECAP_INV_G11
XG9344 XI11_3/XI0/XI0_39/d_9_ XI11_3/XI0/XI0_39/d__9_ DECAP_INV_G11
XG9345 XI11_3/XI0/XI0_39/d_8_ XI11_3/XI0/XI0_39/d__8_ DECAP_INV_G11
XG9346 XI11_3/XI0/XI0_39/d_7_ XI11_3/XI0/XI0_39/d__7_ DECAP_INV_G11
XG9347 XI11_3/XI0/XI0_39/d_6_ XI11_3/XI0/XI0_39/d__6_ DECAP_INV_G11
XG9348 XI11_3/XI0/XI0_39/d_5_ XI11_3/XI0/XI0_39/d__5_ DECAP_INV_G11
XG9349 XI11_3/XI0/XI0_39/d_4_ XI11_3/XI0/XI0_39/d__4_ DECAP_INV_G11
XG9350 XI11_3/XI0/XI0_39/d_3_ XI11_3/XI0/XI0_39/d__3_ DECAP_INV_G11
XG9351 XI11_3/XI0/XI0_39/d_2_ XI11_3/XI0/XI0_39/d__2_ DECAP_INV_G11
XG9352 XI11_3/XI0/XI0_39/d_1_ XI11_3/XI0/XI0_39/d__1_ DECAP_INV_G11
XG9353 XI11_3/XI0/XI0_39/d_0_ XI11_3/XI0/XI0_39/d__0_ DECAP_INV_G11
XG9354 XI11_3/XI0/XI0_38/d__15_ XI11_3/XI0/XI0_38/d_15_ DECAP_INV_G11
XG9355 XI11_3/XI0/XI0_38/d__14_ XI11_3/XI0/XI0_38/d_14_ DECAP_INV_G11
XG9356 XI11_3/XI0/XI0_38/d__13_ XI11_3/XI0/XI0_38/d_13_ DECAP_INV_G11
XG9357 XI11_3/XI0/XI0_38/d__12_ XI11_3/XI0/XI0_38/d_12_ DECAP_INV_G11
XG9358 XI11_3/XI0/XI0_38/d__11_ XI11_3/XI0/XI0_38/d_11_ DECAP_INV_G11
XG9359 XI11_3/XI0/XI0_38/d__10_ XI11_3/XI0/XI0_38/d_10_ DECAP_INV_G11
XG9360 XI11_3/XI0/XI0_38/d__9_ XI11_3/XI0/XI0_38/d_9_ DECAP_INV_G11
XG9361 XI11_3/XI0/XI0_38/d__8_ XI11_3/XI0/XI0_38/d_8_ DECAP_INV_G11
XG9362 XI11_3/XI0/XI0_38/d__7_ XI11_3/XI0/XI0_38/d_7_ DECAP_INV_G11
XG9363 XI11_3/XI0/XI0_38/d__6_ XI11_3/XI0/XI0_38/d_6_ DECAP_INV_G11
XG9364 XI11_3/XI0/XI0_38/d__5_ XI11_3/XI0/XI0_38/d_5_ DECAP_INV_G11
XG9365 XI11_3/XI0/XI0_38/d__4_ XI11_3/XI0/XI0_38/d_4_ DECAP_INV_G11
XG9366 XI11_3/XI0/XI0_38/d__3_ XI11_3/XI0/XI0_38/d_3_ DECAP_INV_G11
XG9367 XI11_3/XI0/XI0_38/d__2_ XI11_3/XI0/XI0_38/d_2_ DECAP_INV_G11
XG9368 XI11_3/XI0/XI0_38/d__1_ XI11_3/XI0/XI0_38/d_1_ DECAP_INV_G11
XG9369 XI11_3/XI0/XI0_38/d__0_ XI11_3/XI0/XI0_38/d_0_ DECAP_INV_G11
XG9370 XI11_3/XI0/XI0_38/d_15_ XI11_3/XI0/XI0_38/d__15_ DECAP_INV_G11
XG9371 XI11_3/XI0/XI0_38/d_14_ XI11_3/XI0/XI0_38/d__14_ DECAP_INV_G11
XG9372 XI11_3/XI0/XI0_38/d_13_ XI11_3/XI0/XI0_38/d__13_ DECAP_INV_G11
XG9373 XI11_3/XI0/XI0_38/d_12_ XI11_3/XI0/XI0_38/d__12_ DECAP_INV_G11
XG9374 XI11_3/XI0/XI0_38/d_11_ XI11_3/XI0/XI0_38/d__11_ DECAP_INV_G11
XG9375 XI11_3/XI0/XI0_38/d_10_ XI11_3/XI0/XI0_38/d__10_ DECAP_INV_G11
XG9376 XI11_3/XI0/XI0_38/d_9_ XI11_3/XI0/XI0_38/d__9_ DECAP_INV_G11
XG9377 XI11_3/XI0/XI0_38/d_8_ XI11_3/XI0/XI0_38/d__8_ DECAP_INV_G11
XG9378 XI11_3/XI0/XI0_38/d_7_ XI11_3/XI0/XI0_38/d__7_ DECAP_INV_G11
XG9379 XI11_3/XI0/XI0_38/d_6_ XI11_3/XI0/XI0_38/d__6_ DECAP_INV_G11
XG9380 XI11_3/XI0/XI0_38/d_5_ XI11_3/XI0/XI0_38/d__5_ DECAP_INV_G11
XG9381 XI11_3/XI0/XI0_38/d_4_ XI11_3/XI0/XI0_38/d__4_ DECAP_INV_G11
XG9382 XI11_3/XI0/XI0_38/d_3_ XI11_3/XI0/XI0_38/d__3_ DECAP_INV_G11
XG9383 XI11_3/XI0/XI0_38/d_2_ XI11_3/XI0/XI0_38/d__2_ DECAP_INV_G11
XG9384 XI11_3/XI0/XI0_38/d_1_ XI11_3/XI0/XI0_38/d__1_ DECAP_INV_G11
XG9385 XI11_3/XI0/XI0_38/d_0_ XI11_3/XI0/XI0_38/d__0_ DECAP_INV_G11
XG9386 XI11_3/XI0/XI0_37/d__15_ XI11_3/XI0/XI0_37/d_15_ DECAP_INV_G11
XG9387 XI11_3/XI0/XI0_37/d__14_ XI11_3/XI0/XI0_37/d_14_ DECAP_INV_G11
XG9388 XI11_3/XI0/XI0_37/d__13_ XI11_3/XI0/XI0_37/d_13_ DECAP_INV_G11
XG9389 XI11_3/XI0/XI0_37/d__12_ XI11_3/XI0/XI0_37/d_12_ DECAP_INV_G11
XG9390 XI11_3/XI0/XI0_37/d__11_ XI11_3/XI0/XI0_37/d_11_ DECAP_INV_G11
XG9391 XI11_3/XI0/XI0_37/d__10_ XI11_3/XI0/XI0_37/d_10_ DECAP_INV_G11
XG9392 XI11_3/XI0/XI0_37/d__9_ XI11_3/XI0/XI0_37/d_9_ DECAP_INV_G11
XG9393 XI11_3/XI0/XI0_37/d__8_ XI11_3/XI0/XI0_37/d_8_ DECAP_INV_G11
XG9394 XI11_3/XI0/XI0_37/d__7_ XI11_3/XI0/XI0_37/d_7_ DECAP_INV_G11
XG9395 XI11_3/XI0/XI0_37/d__6_ XI11_3/XI0/XI0_37/d_6_ DECAP_INV_G11
XG9396 XI11_3/XI0/XI0_37/d__5_ XI11_3/XI0/XI0_37/d_5_ DECAP_INV_G11
XG9397 XI11_3/XI0/XI0_37/d__4_ XI11_3/XI0/XI0_37/d_4_ DECAP_INV_G11
XG9398 XI11_3/XI0/XI0_37/d__3_ XI11_3/XI0/XI0_37/d_3_ DECAP_INV_G11
XG9399 XI11_3/XI0/XI0_37/d__2_ XI11_3/XI0/XI0_37/d_2_ DECAP_INV_G11
XG9400 XI11_3/XI0/XI0_37/d__1_ XI11_3/XI0/XI0_37/d_1_ DECAP_INV_G11
XG9401 XI11_3/XI0/XI0_37/d__0_ XI11_3/XI0/XI0_37/d_0_ DECAP_INV_G11
XG9402 XI11_3/XI0/XI0_37/d_15_ XI11_3/XI0/XI0_37/d__15_ DECAP_INV_G11
XG9403 XI11_3/XI0/XI0_37/d_14_ XI11_3/XI0/XI0_37/d__14_ DECAP_INV_G11
XG9404 XI11_3/XI0/XI0_37/d_13_ XI11_3/XI0/XI0_37/d__13_ DECAP_INV_G11
XG9405 XI11_3/XI0/XI0_37/d_12_ XI11_3/XI0/XI0_37/d__12_ DECAP_INV_G11
XG9406 XI11_3/XI0/XI0_37/d_11_ XI11_3/XI0/XI0_37/d__11_ DECAP_INV_G11
XG9407 XI11_3/XI0/XI0_37/d_10_ XI11_3/XI0/XI0_37/d__10_ DECAP_INV_G11
XG9408 XI11_3/XI0/XI0_37/d_9_ XI11_3/XI0/XI0_37/d__9_ DECAP_INV_G11
XG9409 XI11_3/XI0/XI0_37/d_8_ XI11_3/XI0/XI0_37/d__8_ DECAP_INV_G11
XG9410 XI11_3/XI0/XI0_37/d_7_ XI11_3/XI0/XI0_37/d__7_ DECAP_INV_G11
XG9411 XI11_3/XI0/XI0_37/d_6_ XI11_3/XI0/XI0_37/d__6_ DECAP_INV_G11
XG9412 XI11_3/XI0/XI0_37/d_5_ XI11_3/XI0/XI0_37/d__5_ DECAP_INV_G11
XG9413 XI11_3/XI0/XI0_37/d_4_ XI11_3/XI0/XI0_37/d__4_ DECAP_INV_G11
XG9414 XI11_3/XI0/XI0_37/d_3_ XI11_3/XI0/XI0_37/d__3_ DECAP_INV_G11
XG9415 XI11_3/XI0/XI0_37/d_2_ XI11_3/XI0/XI0_37/d__2_ DECAP_INV_G11
XG9416 XI11_3/XI0/XI0_37/d_1_ XI11_3/XI0/XI0_37/d__1_ DECAP_INV_G11
XG9417 XI11_3/XI0/XI0_37/d_0_ XI11_3/XI0/XI0_37/d__0_ DECAP_INV_G11
XG9418 XI11_3/XI0/XI0_36/d__15_ XI11_3/XI0/XI0_36/d_15_ DECAP_INV_G11
XG9419 XI11_3/XI0/XI0_36/d__14_ XI11_3/XI0/XI0_36/d_14_ DECAP_INV_G11
XG9420 XI11_3/XI0/XI0_36/d__13_ XI11_3/XI0/XI0_36/d_13_ DECAP_INV_G11
XG9421 XI11_3/XI0/XI0_36/d__12_ XI11_3/XI0/XI0_36/d_12_ DECAP_INV_G11
XG9422 XI11_3/XI0/XI0_36/d__11_ XI11_3/XI0/XI0_36/d_11_ DECAP_INV_G11
XG9423 XI11_3/XI0/XI0_36/d__10_ XI11_3/XI0/XI0_36/d_10_ DECAP_INV_G11
XG9424 XI11_3/XI0/XI0_36/d__9_ XI11_3/XI0/XI0_36/d_9_ DECAP_INV_G11
XG9425 XI11_3/XI0/XI0_36/d__8_ XI11_3/XI0/XI0_36/d_8_ DECAP_INV_G11
XG9426 XI11_3/XI0/XI0_36/d__7_ XI11_3/XI0/XI0_36/d_7_ DECAP_INV_G11
XG9427 XI11_3/XI0/XI0_36/d__6_ XI11_3/XI0/XI0_36/d_6_ DECAP_INV_G11
XG9428 XI11_3/XI0/XI0_36/d__5_ XI11_3/XI0/XI0_36/d_5_ DECAP_INV_G11
XG9429 XI11_3/XI0/XI0_36/d__4_ XI11_3/XI0/XI0_36/d_4_ DECAP_INV_G11
XG9430 XI11_3/XI0/XI0_36/d__3_ XI11_3/XI0/XI0_36/d_3_ DECAP_INV_G11
XG9431 XI11_3/XI0/XI0_36/d__2_ XI11_3/XI0/XI0_36/d_2_ DECAP_INV_G11
XG9432 XI11_3/XI0/XI0_36/d__1_ XI11_3/XI0/XI0_36/d_1_ DECAP_INV_G11
XG9433 XI11_3/XI0/XI0_36/d__0_ XI11_3/XI0/XI0_36/d_0_ DECAP_INV_G11
XG9434 XI11_3/XI0/XI0_36/d_15_ XI11_3/XI0/XI0_36/d__15_ DECAP_INV_G11
XG9435 XI11_3/XI0/XI0_36/d_14_ XI11_3/XI0/XI0_36/d__14_ DECAP_INV_G11
XG9436 XI11_3/XI0/XI0_36/d_13_ XI11_3/XI0/XI0_36/d__13_ DECAP_INV_G11
XG9437 XI11_3/XI0/XI0_36/d_12_ XI11_3/XI0/XI0_36/d__12_ DECAP_INV_G11
XG9438 XI11_3/XI0/XI0_36/d_11_ XI11_3/XI0/XI0_36/d__11_ DECAP_INV_G11
XG9439 XI11_3/XI0/XI0_36/d_10_ XI11_3/XI0/XI0_36/d__10_ DECAP_INV_G11
XG9440 XI11_3/XI0/XI0_36/d_9_ XI11_3/XI0/XI0_36/d__9_ DECAP_INV_G11
XG9441 XI11_3/XI0/XI0_36/d_8_ XI11_3/XI0/XI0_36/d__8_ DECAP_INV_G11
XG9442 XI11_3/XI0/XI0_36/d_7_ XI11_3/XI0/XI0_36/d__7_ DECAP_INV_G11
XG9443 XI11_3/XI0/XI0_36/d_6_ XI11_3/XI0/XI0_36/d__6_ DECAP_INV_G11
XG9444 XI11_3/XI0/XI0_36/d_5_ XI11_3/XI0/XI0_36/d__5_ DECAP_INV_G11
XG9445 XI11_3/XI0/XI0_36/d_4_ XI11_3/XI0/XI0_36/d__4_ DECAP_INV_G11
XG9446 XI11_3/XI0/XI0_36/d_3_ XI11_3/XI0/XI0_36/d__3_ DECAP_INV_G11
XG9447 XI11_3/XI0/XI0_36/d_2_ XI11_3/XI0/XI0_36/d__2_ DECAP_INV_G11
XG9448 XI11_3/XI0/XI0_36/d_1_ XI11_3/XI0/XI0_36/d__1_ DECAP_INV_G11
XG9449 XI11_3/XI0/XI0_36/d_0_ XI11_3/XI0/XI0_36/d__0_ DECAP_INV_G11
XG9450 XI11_3/XI0/XI0_35/d__15_ XI11_3/XI0/XI0_35/d_15_ DECAP_INV_G11
XG9451 XI11_3/XI0/XI0_35/d__14_ XI11_3/XI0/XI0_35/d_14_ DECAP_INV_G11
XG9452 XI11_3/XI0/XI0_35/d__13_ XI11_3/XI0/XI0_35/d_13_ DECAP_INV_G11
XG9453 XI11_3/XI0/XI0_35/d__12_ XI11_3/XI0/XI0_35/d_12_ DECAP_INV_G11
XG9454 XI11_3/XI0/XI0_35/d__11_ XI11_3/XI0/XI0_35/d_11_ DECAP_INV_G11
XG9455 XI11_3/XI0/XI0_35/d__10_ XI11_3/XI0/XI0_35/d_10_ DECAP_INV_G11
XG9456 XI11_3/XI0/XI0_35/d__9_ XI11_3/XI0/XI0_35/d_9_ DECAP_INV_G11
XG9457 XI11_3/XI0/XI0_35/d__8_ XI11_3/XI0/XI0_35/d_8_ DECAP_INV_G11
XG9458 XI11_3/XI0/XI0_35/d__7_ XI11_3/XI0/XI0_35/d_7_ DECAP_INV_G11
XG9459 XI11_3/XI0/XI0_35/d__6_ XI11_3/XI0/XI0_35/d_6_ DECAP_INV_G11
XG9460 XI11_3/XI0/XI0_35/d__5_ XI11_3/XI0/XI0_35/d_5_ DECAP_INV_G11
XG9461 XI11_3/XI0/XI0_35/d__4_ XI11_3/XI0/XI0_35/d_4_ DECAP_INV_G11
XG9462 XI11_3/XI0/XI0_35/d__3_ XI11_3/XI0/XI0_35/d_3_ DECAP_INV_G11
XG9463 XI11_3/XI0/XI0_35/d__2_ XI11_3/XI0/XI0_35/d_2_ DECAP_INV_G11
XG9464 XI11_3/XI0/XI0_35/d__1_ XI11_3/XI0/XI0_35/d_1_ DECAP_INV_G11
XG9465 XI11_3/XI0/XI0_35/d__0_ XI11_3/XI0/XI0_35/d_0_ DECAP_INV_G11
XG9466 XI11_3/XI0/XI0_35/d_15_ XI11_3/XI0/XI0_35/d__15_ DECAP_INV_G11
XG9467 XI11_3/XI0/XI0_35/d_14_ XI11_3/XI0/XI0_35/d__14_ DECAP_INV_G11
XG9468 XI11_3/XI0/XI0_35/d_13_ XI11_3/XI0/XI0_35/d__13_ DECAP_INV_G11
XG9469 XI11_3/XI0/XI0_35/d_12_ XI11_3/XI0/XI0_35/d__12_ DECAP_INV_G11
XG9470 XI11_3/XI0/XI0_35/d_11_ XI11_3/XI0/XI0_35/d__11_ DECAP_INV_G11
XG9471 XI11_3/XI0/XI0_35/d_10_ XI11_3/XI0/XI0_35/d__10_ DECAP_INV_G11
XG9472 XI11_3/XI0/XI0_35/d_9_ XI11_3/XI0/XI0_35/d__9_ DECAP_INV_G11
XG9473 XI11_3/XI0/XI0_35/d_8_ XI11_3/XI0/XI0_35/d__8_ DECAP_INV_G11
XG9474 XI11_3/XI0/XI0_35/d_7_ XI11_3/XI0/XI0_35/d__7_ DECAP_INV_G11
XG9475 XI11_3/XI0/XI0_35/d_6_ XI11_3/XI0/XI0_35/d__6_ DECAP_INV_G11
XG9476 XI11_3/XI0/XI0_35/d_5_ XI11_3/XI0/XI0_35/d__5_ DECAP_INV_G11
XG9477 XI11_3/XI0/XI0_35/d_4_ XI11_3/XI0/XI0_35/d__4_ DECAP_INV_G11
XG9478 XI11_3/XI0/XI0_35/d_3_ XI11_3/XI0/XI0_35/d__3_ DECAP_INV_G11
XG9479 XI11_3/XI0/XI0_35/d_2_ XI11_3/XI0/XI0_35/d__2_ DECAP_INV_G11
XG9480 XI11_3/XI0/XI0_35/d_1_ XI11_3/XI0/XI0_35/d__1_ DECAP_INV_G11
XG9481 XI11_3/XI0/XI0_35/d_0_ XI11_3/XI0/XI0_35/d__0_ DECAP_INV_G11
XG9482 XI11_3/XI0/XI0_34/d__15_ XI11_3/XI0/XI0_34/d_15_ DECAP_INV_G11
XG9483 XI11_3/XI0/XI0_34/d__14_ XI11_3/XI0/XI0_34/d_14_ DECAP_INV_G11
XG9484 XI11_3/XI0/XI0_34/d__13_ XI11_3/XI0/XI0_34/d_13_ DECAP_INV_G11
XG9485 XI11_3/XI0/XI0_34/d__12_ XI11_3/XI0/XI0_34/d_12_ DECAP_INV_G11
XG9486 XI11_3/XI0/XI0_34/d__11_ XI11_3/XI0/XI0_34/d_11_ DECAP_INV_G11
XG9487 XI11_3/XI0/XI0_34/d__10_ XI11_3/XI0/XI0_34/d_10_ DECAP_INV_G11
XG9488 XI11_3/XI0/XI0_34/d__9_ XI11_3/XI0/XI0_34/d_9_ DECAP_INV_G11
XG9489 XI11_3/XI0/XI0_34/d__8_ XI11_3/XI0/XI0_34/d_8_ DECAP_INV_G11
XG9490 XI11_3/XI0/XI0_34/d__7_ XI11_3/XI0/XI0_34/d_7_ DECAP_INV_G11
XG9491 XI11_3/XI0/XI0_34/d__6_ XI11_3/XI0/XI0_34/d_6_ DECAP_INV_G11
XG9492 XI11_3/XI0/XI0_34/d__5_ XI11_3/XI0/XI0_34/d_5_ DECAP_INV_G11
XG9493 XI11_3/XI0/XI0_34/d__4_ XI11_3/XI0/XI0_34/d_4_ DECAP_INV_G11
XG9494 XI11_3/XI0/XI0_34/d__3_ XI11_3/XI0/XI0_34/d_3_ DECAP_INV_G11
XG9495 XI11_3/XI0/XI0_34/d__2_ XI11_3/XI0/XI0_34/d_2_ DECAP_INV_G11
XG9496 XI11_3/XI0/XI0_34/d__1_ XI11_3/XI0/XI0_34/d_1_ DECAP_INV_G11
XG9497 XI11_3/XI0/XI0_34/d__0_ XI11_3/XI0/XI0_34/d_0_ DECAP_INV_G11
XG9498 XI11_3/XI0/XI0_34/d_15_ XI11_3/XI0/XI0_34/d__15_ DECAP_INV_G11
XG9499 XI11_3/XI0/XI0_34/d_14_ XI11_3/XI0/XI0_34/d__14_ DECAP_INV_G11
XG9500 XI11_3/XI0/XI0_34/d_13_ XI11_3/XI0/XI0_34/d__13_ DECAP_INV_G11
XG9501 XI11_3/XI0/XI0_34/d_12_ XI11_3/XI0/XI0_34/d__12_ DECAP_INV_G11
XG9502 XI11_3/XI0/XI0_34/d_11_ XI11_3/XI0/XI0_34/d__11_ DECAP_INV_G11
XG9503 XI11_3/XI0/XI0_34/d_10_ XI11_3/XI0/XI0_34/d__10_ DECAP_INV_G11
XG9504 XI11_3/XI0/XI0_34/d_9_ XI11_3/XI0/XI0_34/d__9_ DECAP_INV_G11
XG9505 XI11_3/XI0/XI0_34/d_8_ XI11_3/XI0/XI0_34/d__8_ DECAP_INV_G11
XG9506 XI11_3/XI0/XI0_34/d_7_ XI11_3/XI0/XI0_34/d__7_ DECAP_INV_G11
XG9507 XI11_3/XI0/XI0_34/d_6_ XI11_3/XI0/XI0_34/d__6_ DECAP_INV_G11
XG9508 XI11_3/XI0/XI0_34/d_5_ XI11_3/XI0/XI0_34/d__5_ DECAP_INV_G11
XG9509 XI11_3/XI0/XI0_34/d_4_ XI11_3/XI0/XI0_34/d__4_ DECAP_INV_G11
XG9510 XI11_3/XI0/XI0_34/d_3_ XI11_3/XI0/XI0_34/d__3_ DECAP_INV_G11
XG9511 XI11_3/XI0/XI0_34/d_2_ XI11_3/XI0/XI0_34/d__2_ DECAP_INV_G11
XG9512 XI11_3/XI0/XI0_34/d_1_ XI11_3/XI0/XI0_34/d__1_ DECAP_INV_G11
XG9513 XI11_3/XI0/XI0_34/d_0_ XI11_3/XI0/XI0_34/d__0_ DECAP_INV_G11
XG9514 XI11_3/XI0/XI0_33/d__15_ XI11_3/XI0/XI0_33/d_15_ DECAP_INV_G11
XG9515 XI11_3/XI0/XI0_33/d__14_ XI11_3/XI0/XI0_33/d_14_ DECAP_INV_G11
XG9516 XI11_3/XI0/XI0_33/d__13_ XI11_3/XI0/XI0_33/d_13_ DECAP_INV_G11
XG9517 XI11_3/XI0/XI0_33/d__12_ XI11_3/XI0/XI0_33/d_12_ DECAP_INV_G11
XG9518 XI11_3/XI0/XI0_33/d__11_ XI11_3/XI0/XI0_33/d_11_ DECAP_INV_G11
XG9519 XI11_3/XI0/XI0_33/d__10_ XI11_3/XI0/XI0_33/d_10_ DECAP_INV_G11
XG9520 XI11_3/XI0/XI0_33/d__9_ XI11_3/XI0/XI0_33/d_9_ DECAP_INV_G11
XG9521 XI11_3/XI0/XI0_33/d__8_ XI11_3/XI0/XI0_33/d_8_ DECAP_INV_G11
XG9522 XI11_3/XI0/XI0_33/d__7_ XI11_3/XI0/XI0_33/d_7_ DECAP_INV_G11
XG9523 XI11_3/XI0/XI0_33/d__6_ XI11_3/XI0/XI0_33/d_6_ DECAP_INV_G11
XG9524 XI11_3/XI0/XI0_33/d__5_ XI11_3/XI0/XI0_33/d_5_ DECAP_INV_G11
XG9525 XI11_3/XI0/XI0_33/d__4_ XI11_3/XI0/XI0_33/d_4_ DECAP_INV_G11
XG9526 XI11_3/XI0/XI0_33/d__3_ XI11_3/XI0/XI0_33/d_3_ DECAP_INV_G11
XG9527 XI11_3/XI0/XI0_33/d__2_ XI11_3/XI0/XI0_33/d_2_ DECAP_INV_G11
XG9528 XI11_3/XI0/XI0_33/d__1_ XI11_3/XI0/XI0_33/d_1_ DECAP_INV_G11
XG9529 XI11_3/XI0/XI0_33/d__0_ XI11_3/XI0/XI0_33/d_0_ DECAP_INV_G11
XG9530 XI11_3/XI0/XI0_33/d_15_ XI11_3/XI0/XI0_33/d__15_ DECAP_INV_G11
XG9531 XI11_3/XI0/XI0_33/d_14_ XI11_3/XI0/XI0_33/d__14_ DECAP_INV_G11
XG9532 XI11_3/XI0/XI0_33/d_13_ XI11_3/XI0/XI0_33/d__13_ DECAP_INV_G11
XG9533 XI11_3/XI0/XI0_33/d_12_ XI11_3/XI0/XI0_33/d__12_ DECAP_INV_G11
XG9534 XI11_3/XI0/XI0_33/d_11_ XI11_3/XI0/XI0_33/d__11_ DECAP_INV_G11
XG9535 XI11_3/XI0/XI0_33/d_10_ XI11_3/XI0/XI0_33/d__10_ DECAP_INV_G11
XG9536 XI11_3/XI0/XI0_33/d_9_ XI11_3/XI0/XI0_33/d__9_ DECAP_INV_G11
XG9537 XI11_3/XI0/XI0_33/d_8_ XI11_3/XI0/XI0_33/d__8_ DECAP_INV_G11
XG9538 XI11_3/XI0/XI0_33/d_7_ XI11_3/XI0/XI0_33/d__7_ DECAP_INV_G11
XG9539 XI11_3/XI0/XI0_33/d_6_ XI11_3/XI0/XI0_33/d__6_ DECAP_INV_G11
XG9540 XI11_3/XI0/XI0_33/d_5_ XI11_3/XI0/XI0_33/d__5_ DECAP_INV_G11
XG9541 XI11_3/XI0/XI0_33/d_4_ XI11_3/XI0/XI0_33/d__4_ DECAP_INV_G11
XG9542 XI11_3/XI0/XI0_33/d_3_ XI11_3/XI0/XI0_33/d__3_ DECAP_INV_G11
XG9543 XI11_3/XI0/XI0_33/d_2_ XI11_3/XI0/XI0_33/d__2_ DECAP_INV_G11
XG9544 XI11_3/XI0/XI0_33/d_1_ XI11_3/XI0/XI0_33/d__1_ DECAP_INV_G11
XG9545 XI11_3/XI0/XI0_33/d_0_ XI11_3/XI0/XI0_33/d__0_ DECAP_INV_G11
XG9546 XI11_3/XI0/XI0_32/d__15_ XI11_3/XI0/XI0_32/d_15_ DECAP_INV_G11
XG9547 XI11_3/XI0/XI0_32/d__14_ XI11_3/XI0/XI0_32/d_14_ DECAP_INV_G11
XG9548 XI11_3/XI0/XI0_32/d__13_ XI11_3/XI0/XI0_32/d_13_ DECAP_INV_G11
XG9549 XI11_3/XI0/XI0_32/d__12_ XI11_3/XI0/XI0_32/d_12_ DECAP_INV_G11
XG9550 XI11_3/XI0/XI0_32/d__11_ XI11_3/XI0/XI0_32/d_11_ DECAP_INV_G11
XG9551 XI11_3/XI0/XI0_32/d__10_ XI11_3/XI0/XI0_32/d_10_ DECAP_INV_G11
XG9552 XI11_3/XI0/XI0_32/d__9_ XI11_3/XI0/XI0_32/d_9_ DECAP_INV_G11
XG9553 XI11_3/XI0/XI0_32/d__8_ XI11_3/XI0/XI0_32/d_8_ DECAP_INV_G11
XG9554 XI11_3/XI0/XI0_32/d__7_ XI11_3/XI0/XI0_32/d_7_ DECAP_INV_G11
XG9555 XI11_3/XI0/XI0_32/d__6_ XI11_3/XI0/XI0_32/d_6_ DECAP_INV_G11
XG9556 XI11_3/XI0/XI0_32/d__5_ XI11_3/XI0/XI0_32/d_5_ DECAP_INV_G11
XG9557 XI11_3/XI0/XI0_32/d__4_ XI11_3/XI0/XI0_32/d_4_ DECAP_INV_G11
XG9558 XI11_3/XI0/XI0_32/d__3_ XI11_3/XI0/XI0_32/d_3_ DECAP_INV_G11
XG9559 XI11_3/XI0/XI0_32/d__2_ XI11_3/XI0/XI0_32/d_2_ DECAP_INV_G11
XG9560 XI11_3/XI0/XI0_32/d__1_ XI11_3/XI0/XI0_32/d_1_ DECAP_INV_G11
XG9561 XI11_3/XI0/XI0_32/d__0_ XI11_3/XI0/XI0_32/d_0_ DECAP_INV_G11
XG9562 XI11_3/XI0/XI0_32/d_15_ XI11_3/XI0/XI0_32/d__15_ DECAP_INV_G11
XG9563 XI11_3/XI0/XI0_32/d_14_ XI11_3/XI0/XI0_32/d__14_ DECAP_INV_G11
XG9564 XI11_3/XI0/XI0_32/d_13_ XI11_3/XI0/XI0_32/d__13_ DECAP_INV_G11
XG9565 XI11_3/XI0/XI0_32/d_12_ XI11_3/XI0/XI0_32/d__12_ DECAP_INV_G11
XG9566 XI11_3/XI0/XI0_32/d_11_ XI11_3/XI0/XI0_32/d__11_ DECAP_INV_G11
XG9567 XI11_3/XI0/XI0_32/d_10_ XI11_3/XI0/XI0_32/d__10_ DECAP_INV_G11
XG9568 XI11_3/XI0/XI0_32/d_9_ XI11_3/XI0/XI0_32/d__9_ DECAP_INV_G11
XG9569 XI11_3/XI0/XI0_32/d_8_ XI11_3/XI0/XI0_32/d__8_ DECAP_INV_G11
XG9570 XI11_3/XI0/XI0_32/d_7_ XI11_3/XI0/XI0_32/d__7_ DECAP_INV_G11
XG9571 XI11_3/XI0/XI0_32/d_6_ XI11_3/XI0/XI0_32/d__6_ DECAP_INV_G11
XG9572 XI11_3/XI0/XI0_32/d_5_ XI11_3/XI0/XI0_32/d__5_ DECAP_INV_G11
XG9573 XI11_3/XI0/XI0_32/d_4_ XI11_3/XI0/XI0_32/d__4_ DECAP_INV_G11
XG9574 XI11_3/XI0/XI0_32/d_3_ XI11_3/XI0/XI0_32/d__3_ DECAP_INV_G11
XG9575 XI11_3/XI0/XI0_32/d_2_ XI11_3/XI0/XI0_32/d__2_ DECAP_INV_G11
XG9576 XI11_3/XI0/XI0_32/d_1_ XI11_3/XI0/XI0_32/d__1_ DECAP_INV_G11
XG9577 XI11_3/XI0/XI0_32/d_0_ XI11_3/XI0/XI0_32/d__0_ DECAP_INV_G11
XG9578 XI11_3/XI0/XI0_31/d__15_ XI11_3/XI0/XI0_31/d_15_ DECAP_INV_G11
XG9579 XI11_3/XI0/XI0_31/d__14_ XI11_3/XI0/XI0_31/d_14_ DECAP_INV_G11
XG9580 XI11_3/XI0/XI0_31/d__13_ XI11_3/XI0/XI0_31/d_13_ DECAP_INV_G11
XG9581 XI11_3/XI0/XI0_31/d__12_ XI11_3/XI0/XI0_31/d_12_ DECAP_INV_G11
XG9582 XI11_3/XI0/XI0_31/d__11_ XI11_3/XI0/XI0_31/d_11_ DECAP_INV_G11
XG9583 XI11_3/XI0/XI0_31/d__10_ XI11_3/XI0/XI0_31/d_10_ DECAP_INV_G11
XG9584 XI11_3/XI0/XI0_31/d__9_ XI11_3/XI0/XI0_31/d_9_ DECAP_INV_G11
XG9585 XI11_3/XI0/XI0_31/d__8_ XI11_3/XI0/XI0_31/d_8_ DECAP_INV_G11
XG9586 XI11_3/XI0/XI0_31/d__7_ XI11_3/XI0/XI0_31/d_7_ DECAP_INV_G11
XG9587 XI11_3/XI0/XI0_31/d__6_ XI11_3/XI0/XI0_31/d_6_ DECAP_INV_G11
XG9588 XI11_3/XI0/XI0_31/d__5_ XI11_3/XI0/XI0_31/d_5_ DECAP_INV_G11
XG9589 XI11_3/XI0/XI0_31/d__4_ XI11_3/XI0/XI0_31/d_4_ DECAP_INV_G11
XG9590 XI11_3/XI0/XI0_31/d__3_ XI11_3/XI0/XI0_31/d_3_ DECAP_INV_G11
XG9591 XI11_3/XI0/XI0_31/d__2_ XI11_3/XI0/XI0_31/d_2_ DECAP_INV_G11
XG9592 XI11_3/XI0/XI0_31/d__1_ XI11_3/XI0/XI0_31/d_1_ DECAP_INV_G11
XG9593 XI11_3/XI0/XI0_31/d__0_ XI11_3/XI0/XI0_31/d_0_ DECAP_INV_G11
XG9594 XI11_3/XI0/XI0_31/d_15_ XI11_3/XI0/XI0_31/d__15_ DECAP_INV_G11
XG9595 XI11_3/XI0/XI0_31/d_14_ XI11_3/XI0/XI0_31/d__14_ DECAP_INV_G11
XG9596 XI11_3/XI0/XI0_31/d_13_ XI11_3/XI0/XI0_31/d__13_ DECAP_INV_G11
XG9597 XI11_3/XI0/XI0_31/d_12_ XI11_3/XI0/XI0_31/d__12_ DECAP_INV_G11
XG9598 XI11_3/XI0/XI0_31/d_11_ XI11_3/XI0/XI0_31/d__11_ DECAP_INV_G11
XG9599 XI11_3/XI0/XI0_31/d_10_ XI11_3/XI0/XI0_31/d__10_ DECAP_INV_G11
XG9600 XI11_3/XI0/XI0_31/d_9_ XI11_3/XI0/XI0_31/d__9_ DECAP_INV_G11
XG9601 XI11_3/XI0/XI0_31/d_8_ XI11_3/XI0/XI0_31/d__8_ DECAP_INV_G11
XG9602 XI11_3/XI0/XI0_31/d_7_ XI11_3/XI0/XI0_31/d__7_ DECAP_INV_G11
XG9603 XI11_3/XI0/XI0_31/d_6_ XI11_3/XI0/XI0_31/d__6_ DECAP_INV_G11
XG9604 XI11_3/XI0/XI0_31/d_5_ XI11_3/XI0/XI0_31/d__5_ DECAP_INV_G11
XG9605 XI11_3/XI0/XI0_31/d_4_ XI11_3/XI0/XI0_31/d__4_ DECAP_INV_G11
XG9606 XI11_3/XI0/XI0_31/d_3_ XI11_3/XI0/XI0_31/d__3_ DECAP_INV_G11
XG9607 XI11_3/XI0/XI0_31/d_2_ XI11_3/XI0/XI0_31/d__2_ DECAP_INV_G11
XG9608 XI11_3/XI0/XI0_31/d_1_ XI11_3/XI0/XI0_31/d__1_ DECAP_INV_G11
XG9609 XI11_3/XI0/XI0_31/d_0_ XI11_3/XI0/XI0_31/d__0_ DECAP_INV_G11
XG9610 XI11_3/XI0/XI0_30/d__15_ XI11_3/XI0/XI0_30/d_15_ DECAP_INV_G11
XG9611 XI11_3/XI0/XI0_30/d__14_ XI11_3/XI0/XI0_30/d_14_ DECAP_INV_G11
XG9612 XI11_3/XI0/XI0_30/d__13_ XI11_3/XI0/XI0_30/d_13_ DECAP_INV_G11
XG9613 XI11_3/XI0/XI0_30/d__12_ XI11_3/XI0/XI0_30/d_12_ DECAP_INV_G11
XG9614 XI11_3/XI0/XI0_30/d__11_ XI11_3/XI0/XI0_30/d_11_ DECAP_INV_G11
XG9615 XI11_3/XI0/XI0_30/d__10_ XI11_3/XI0/XI0_30/d_10_ DECAP_INV_G11
XG9616 XI11_3/XI0/XI0_30/d__9_ XI11_3/XI0/XI0_30/d_9_ DECAP_INV_G11
XG9617 XI11_3/XI0/XI0_30/d__8_ XI11_3/XI0/XI0_30/d_8_ DECAP_INV_G11
XG9618 XI11_3/XI0/XI0_30/d__7_ XI11_3/XI0/XI0_30/d_7_ DECAP_INV_G11
XG9619 XI11_3/XI0/XI0_30/d__6_ XI11_3/XI0/XI0_30/d_6_ DECAP_INV_G11
XG9620 XI11_3/XI0/XI0_30/d__5_ XI11_3/XI0/XI0_30/d_5_ DECAP_INV_G11
XG9621 XI11_3/XI0/XI0_30/d__4_ XI11_3/XI0/XI0_30/d_4_ DECAP_INV_G11
XG9622 XI11_3/XI0/XI0_30/d__3_ XI11_3/XI0/XI0_30/d_3_ DECAP_INV_G11
XG9623 XI11_3/XI0/XI0_30/d__2_ XI11_3/XI0/XI0_30/d_2_ DECAP_INV_G11
XG9624 XI11_3/XI0/XI0_30/d__1_ XI11_3/XI0/XI0_30/d_1_ DECAP_INV_G11
XG9625 XI11_3/XI0/XI0_30/d__0_ XI11_3/XI0/XI0_30/d_0_ DECAP_INV_G11
XG9626 XI11_3/XI0/XI0_30/d_15_ XI11_3/XI0/XI0_30/d__15_ DECAP_INV_G11
XG9627 XI11_3/XI0/XI0_30/d_14_ XI11_3/XI0/XI0_30/d__14_ DECAP_INV_G11
XG9628 XI11_3/XI0/XI0_30/d_13_ XI11_3/XI0/XI0_30/d__13_ DECAP_INV_G11
XG9629 XI11_3/XI0/XI0_30/d_12_ XI11_3/XI0/XI0_30/d__12_ DECAP_INV_G11
XG9630 XI11_3/XI0/XI0_30/d_11_ XI11_3/XI0/XI0_30/d__11_ DECAP_INV_G11
XG9631 XI11_3/XI0/XI0_30/d_10_ XI11_3/XI0/XI0_30/d__10_ DECAP_INV_G11
XG9632 XI11_3/XI0/XI0_30/d_9_ XI11_3/XI0/XI0_30/d__9_ DECAP_INV_G11
XG9633 XI11_3/XI0/XI0_30/d_8_ XI11_3/XI0/XI0_30/d__8_ DECAP_INV_G11
XG9634 XI11_3/XI0/XI0_30/d_7_ XI11_3/XI0/XI0_30/d__7_ DECAP_INV_G11
XG9635 XI11_3/XI0/XI0_30/d_6_ XI11_3/XI0/XI0_30/d__6_ DECAP_INV_G11
XG9636 XI11_3/XI0/XI0_30/d_5_ XI11_3/XI0/XI0_30/d__5_ DECAP_INV_G11
XG9637 XI11_3/XI0/XI0_30/d_4_ XI11_3/XI0/XI0_30/d__4_ DECAP_INV_G11
XG9638 XI11_3/XI0/XI0_30/d_3_ XI11_3/XI0/XI0_30/d__3_ DECAP_INV_G11
XG9639 XI11_3/XI0/XI0_30/d_2_ XI11_3/XI0/XI0_30/d__2_ DECAP_INV_G11
XG9640 XI11_3/XI0/XI0_30/d_1_ XI11_3/XI0/XI0_30/d__1_ DECAP_INV_G11
XG9641 XI11_3/XI0/XI0_30/d_0_ XI11_3/XI0/XI0_30/d__0_ DECAP_INV_G11
XG9642 XI11_3/XI0/XI0_29/d__15_ XI11_3/XI0/XI0_29/d_15_ DECAP_INV_G11
XG9643 XI11_3/XI0/XI0_29/d__14_ XI11_3/XI0/XI0_29/d_14_ DECAP_INV_G11
XG9644 XI11_3/XI0/XI0_29/d__13_ XI11_3/XI0/XI0_29/d_13_ DECAP_INV_G11
XG9645 XI11_3/XI0/XI0_29/d__12_ XI11_3/XI0/XI0_29/d_12_ DECAP_INV_G11
XG9646 XI11_3/XI0/XI0_29/d__11_ XI11_3/XI0/XI0_29/d_11_ DECAP_INV_G11
XG9647 XI11_3/XI0/XI0_29/d__10_ XI11_3/XI0/XI0_29/d_10_ DECAP_INV_G11
XG9648 XI11_3/XI0/XI0_29/d__9_ XI11_3/XI0/XI0_29/d_9_ DECAP_INV_G11
XG9649 XI11_3/XI0/XI0_29/d__8_ XI11_3/XI0/XI0_29/d_8_ DECAP_INV_G11
XG9650 XI11_3/XI0/XI0_29/d__7_ XI11_3/XI0/XI0_29/d_7_ DECAP_INV_G11
XG9651 XI11_3/XI0/XI0_29/d__6_ XI11_3/XI0/XI0_29/d_6_ DECAP_INV_G11
XG9652 XI11_3/XI0/XI0_29/d__5_ XI11_3/XI0/XI0_29/d_5_ DECAP_INV_G11
XG9653 XI11_3/XI0/XI0_29/d__4_ XI11_3/XI0/XI0_29/d_4_ DECAP_INV_G11
XG9654 XI11_3/XI0/XI0_29/d__3_ XI11_3/XI0/XI0_29/d_3_ DECAP_INV_G11
XG9655 XI11_3/XI0/XI0_29/d__2_ XI11_3/XI0/XI0_29/d_2_ DECAP_INV_G11
XG9656 XI11_3/XI0/XI0_29/d__1_ XI11_3/XI0/XI0_29/d_1_ DECAP_INV_G11
XG9657 XI11_3/XI0/XI0_29/d__0_ XI11_3/XI0/XI0_29/d_0_ DECAP_INV_G11
XG9658 XI11_3/XI0/XI0_29/d_15_ XI11_3/XI0/XI0_29/d__15_ DECAP_INV_G11
XG9659 XI11_3/XI0/XI0_29/d_14_ XI11_3/XI0/XI0_29/d__14_ DECAP_INV_G11
XG9660 XI11_3/XI0/XI0_29/d_13_ XI11_3/XI0/XI0_29/d__13_ DECAP_INV_G11
XG9661 XI11_3/XI0/XI0_29/d_12_ XI11_3/XI0/XI0_29/d__12_ DECAP_INV_G11
XG9662 XI11_3/XI0/XI0_29/d_11_ XI11_3/XI0/XI0_29/d__11_ DECAP_INV_G11
XG9663 XI11_3/XI0/XI0_29/d_10_ XI11_3/XI0/XI0_29/d__10_ DECAP_INV_G11
XG9664 XI11_3/XI0/XI0_29/d_9_ XI11_3/XI0/XI0_29/d__9_ DECAP_INV_G11
XG9665 XI11_3/XI0/XI0_29/d_8_ XI11_3/XI0/XI0_29/d__8_ DECAP_INV_G11
XG9666 XI11_3/XI0/XI0_29/d_7_ XI11_3/XI0/XI0_29/d__7_ DECAP_INV_G11
XG9667 XI11_3/XI0/XI0_29/d_6_ XI11_3/XI0/XI0_29/d__6_ DECAP_INV_G11
XG9668 XI11_3/XI0/XI0_29/d_5_ XI11_3/XI0/XI0_29/d__5_ DECAP_INV_G11
XG9669 XI11_3/XI0/XI0_29/d_4_ XI11_3/XI0/XI0_29/d__4_ DECAP_INV_G11
XG9670 XI11_3/XI0/XI0_29/d_3_ XI11_3/XI0/XI0_29/d__3_ DECAP_INV_G11
XG9671 XI11_3/XI0/XI0_29/d_2_ XI11_3/XI0/XI0_29/d__2_ DECAP_INV_G11
XG9672 XI11_3/XI0/XI0_29/d_1_ XI11_3/XI0/XI0_29/d__1_ DECAP_INV_G11
XG9673 XI11_3/XI0/XI0_29/d_0_ XI11_3/XI0/XI0_29/d__0_ DECAP_INV_G11
XG9674 XI11_3/XI0/XI0_28/d__15_ XI11_3/XI0/XI0_28/d_15_ DECAP_INV_G11
XG9675 XI11_3/XI0/XI0_28/d__14_ XI11_3/XI0/XI0_28/d_14_ DECAP_INV_G11
XG9676 XI11_3/XI0/XI0_28/d__13_ XI11_3/XI0/XI0_28/d_13_ DECAP_INV_G11
XG9677 XI11_3/XI0/XI0_28/d__12_ XI11_3/XI0/XI0_28/d_12_ DECAP_INV_G11
XG9678 XI11_3/XI0/XI0_28/d__11_ XI11_3/XI0/XI0_28/d_11_ DECAP_INV_G11
XG9679 XI11_3/XI0/XI0_28/d__10_ XI11_3/XI0/XI0_28/d_10_ DECAP_INV_G11
XG9680 XI11_3/XI0/XI0_28/d__9_ XI11_3/XI0/XI0_28/d_9_ DECAP_INV_G11
XG9681 XI11_3/XI0/XI0_28/d__8_ XI11_3/XI0/XI0_28/d_8_ DECAP_INV_G11
XG9682 XI11_3/XI0/XI0_28/d__7_ XI11_3/XI0/XI0_28/d_7_ DECAP_INV_G11
XG9683 XI11_3/XI0/XI0_28/d__6_ XI11_3/XI0/XI0_28/d_6_ DECAP_INV_G11
XG9684 XI11_3/XI0/XI0_28/d__5_ XI11_3/XI0/XI0_28/d_5_ DECAP_INV_G11
XG9685 XI11_3/XI0/XI0_28/d__4_ XI11_3/XI0/XI0_28/d_4_ DECAP_INV_G11
XG9686 XI11_3/XI0/XI0_28/d__3_ XI11_3/XI0/XI0_28/d_3_ DECAP_INV_G11
XG9687 XI11_3/XI0/XI0_28/d__2_ XI11_3/XI0/XI0_28/d_2_ DECAP_INV_G11
XG9688 XI11_3/XI0/XI0_28/d__1_ XI11_3/XI0/XI0_28/d_1_ DECAP_INV_G11
XG9689 XI11_3/XI0/XI0_28/d__0_ XI11_3/XI0/XI0_28/d_0_ DECAP_INV_G11
XG9690 XI11_3/XI0/XI0_28/d_15_ XI11_3/XI0/XI0_28/d__15_ DECAP_INV_G11
XG9691 XI11_3/XI0/XI0_28/d_14_ XI11_3/XI0/XI0_28/d__14_ DECAP_INV_G11
XG9692 XI11_3/XI0/XI0_28/d_13_ XI11_3/XI0/XI0_28/d__13_ DECAP_INV_G11
XG9693 XI11_3/XI0/XI0_28/d_12_ XI11_3/XI0/XI0_28/d__12_ DECAP_INV_G11
XG9694 XI11_3/XI0/XI0_28/d_11_ XI11_3/XI0/XI0_28/d__11_ DECAP_INV_G11
XG9695 XI11_3/XI0/XI0_28/d_10_ XI11_3/XI0/XI0_28/d__10_ DECAP_INV_G11
XG9696 XI11_3/XI0/XI0_28/d_9_ XI11_3/XI0/XI0_28/d__9_ DECAP_INV_G11
XG9697 XI11_3/XI0/XI0_28/d_8_ XI11_3/XI0/XI0_28/d__8_ DECAP_INV_G11
XG9698 XI11_3/XI0/XI0_28/d_7_ XI11_3/XI0/XI0_28/d__7_ DECAP_INV_G11
XG9699 XI11_3/XI0/XI0_28/d_6_ XI11_3/XI0/XI0_28/d__6_ DECAP_INV_G11
XG9700 XI11_3/XI0/XI0_28/d_5_ XI11_3/XI0/XI0_28/d__5_ DECAP_INV_G11
XG9701 XI11_3/XI0/XI0_28/d_4_ XI11_3/XI0/XI0_28/d__4_ DECAP_INV_G11
XG9702 XI11_3/XI0/XI0_28/d_3_ XI11_3/XI0/XI0_28/d__3_ DECAP_INV_G11
XG9703 XI11_3/XI0/XI0_28/d_2_ XI11_3/XI0/XI0_28/d__2_ DECAP_INV_G11
XG9704 XI11_3/XI0/XI0_28/d_1_ XI11_3/XI0/XI0_28/d__1_ DECAP_INV_G11
XG9705 XI11_3/XI0/XI0_28/d_0_ XI11_3/XI0/XI0_28/d__0_ DECAP_INV_G11
XG9706 XI11_3/XI0/XI0_27/d__15_ XI11_3/XI0/XI0_27/d_15_ DECAP_INV_G11
XG9707 XI11_3/XI0/XI0_27/d__14_ XI11_3/XI0/XI0_27/d_14_ DECAP_INV_G11
XG9708 XI11_3/XI0/XI0_27/d__13_ XI11_3/XI0/XI0_27/d_13_ DECAP_INV_G11
XG9709 XI11_3/XI0/XI0_27/d__12_ XI11_3/XI0/XI0_27/d_12_ DECAP_INV_G11
XG9710 XI11_3/XI0/XI0_27/d__11_ XI11_3/XI0/XI0_27/d_11_ DECAP_INV_G11
XG9711 XI11_3/XI0/XI0_27/d__10_ XI11_3/XI0/XI0_27/d_10_ DECAP_INV_G11
XG9712 XI11_3/XI0/XI0_27/d__9_ XI11_3/XI0/XI0_27/d_9_ DECAP_INV_G11
XG9713 XI11_3/XI0/XI0_27/d__8_ XI11_3/XI0/XI0_27/d_8_ DECAP_INV_G11
XG9714 XI11_3/XI0/XI0_27/d__7_ XI11_3/XI0/XI0_27/d_7_ DECAP_INV_G11
XG9715 XI11_3/XI0/XI0_27/d__6_ XI11_3/XI0/XI0_27/d_6_ DECAP_INV_G11
XG9716 XI11_3/XI0/XI0_27/d__5_ XI11_3/XI0/XI0_27/d_5_ DECAP_INV_G11
XG9717 XI11_3/XI0/XI0_27/d__4_ XI11_3/XI0/XI0_27/d_4_ DECAP_INV_G11
XG9718 XI11_3/XI0/XI0_27/d__3_ XI11_3/XI0/XI0_27/d_3_ DECAP_INV_G11
XG9719 XI11_3/XI0/XI0_27/d__2_ XI11_3/XI0/XI0_27/d_2_ DECAP_INV_G11
XG9720 XI11_3/XI0/XI0_27/d__1_ XI11_3/XI0/XI0_27/d_1_ DECAP_INV_G11
XG9721 XI11_3/XI0/XI0_27/d__0_ XI11_3/XI0/XI0_27/d_0_ DECAP_INV_G11
XG9722 XI11_3/XI0/XI0_27/d_15_ XI11_3/XI0/XI0_27/d__15_ DECAP_INV_G11
XG9723 XI11_3/XI0/XI0_27/d_14_ XI11_3/XI0/XI0_27/d__14_ DECAP_INV_G11
XG9724 XI11_3/XI0/XI0_27/d_13_ XI11_3/XI0/XI0_27/d__13_ DECAP_INV_G11
XG9725 XI11_3/XI0/XI0_27/d_12_ XI11_3/XI0/XI0_27/d__12_ DECAP_INV_G11
XG9726 XI11_3/XI0/XI0_27/d_11_ XI11_3/XI0/XI0_27/d__11_ DECAP_INV_G11
XG9727 XI11_3/XI0/XI0_27/d_10_ XI11_3/XI0/XI0_27/d__10_ DECAP_INV_G11
XG9728 XI11_3/XI0/XI0_27/d_9_ XI11_3/XI0/XI0_27/d__9_ DECAP_INV_G11
XG9729 XI11_3/XI0/XI0_27/d_8_ XI11_3/XI0/XI0_27/d__8_ DECAP_INV_G11
XG9730 XI11_3/XI0/XI0_27/d_7_ XI11_3/XI0/XI0_27/d__7_ DECAP_INV_G11
XG9731 XI11_3/XI0/XI0_27/d_6_ XI11_3/XI0/XI0_27/d__6_ DECAP_INV_G11
XG9732 XI11_3/XI0/XI0_27/d_5_ XI11_3/XI0/XI0_27/d__5_ DECAP_INV_G11
XG9733 XI11_3/XI0/XI0_27/d_4_ XI11_3/XI0/XI0_27/d__4_ DECAP_INV_G11
XG9734 XI11_3/XI0/XI0_27/d_3_ XI11_3/XI0/XI0_27/d__3_ DECAP_INV_G11
XG9735 XI11_3/XI0/XI0_27/d_2_ XI11_3/XI0/XI0_27/d__2_ DECAP_INV_G11
XG9736 XI11_3/XI0/XI0_27/d_1_ XI11_3/XI0/XI0_27/d__1_ DECAP_INV_G11
XG9737 XI11_3/XI0/XI0_27/d_0_ XI11_3/XI0/XI0_27/d__0_ DECAP_INV_G11
XG9738 XI11_3/XI0/XI0_26/d__15_ XI11_3/XI0/XI0_26/d_15_ DECAP_INV_G11
XG9739 XI11_3/XI0/XI0_26/d__14_ XI11_3/XI0/XI0_26/d_14_ DECAP_INV_G11
XG9740 XI11_3/XI0/XI0_26/d__13_ XI11_3/XI0/XI0_26/d_13_ DECAP_INV_G11
XG9741 XI11_3/XI0/XI0_26/d__12_ XI11_3/XI0/XI0_26/d_12_ DECAP_INV_G11
XG9742 XI11_3/XI0/XI0_26/d__11_ XI11_3/XI0/XI0_26/d_11_ DECAP_INV_G11
XG9743 XI11_3/XI0/XI0_26/d__10_ XI11_3/XI0/XI0_26/d_10_ DECAP_INV_G11
XG9744 XI11_3/XI0/XI0_26/d__9_ XI11_3/XI0/XI0_26/d_9_ DECAP_INV_G11
XG9745 XI11_3/XI0/XI0_26/d__8_ XI11_3/XI0/XI0_26/d_8_ DECAP_INV_G11
XG9746 XI11_3/XI0/XI0_26/d__7_ XI11_3/XI0/XI0_26/d_7_ DECAP_INV_G11
XG9747 XI11_3/XI0/XI0_26/d__6_ XI11_3/XI0/XI0_26/d_6_ DECAP_INV_G11
XG9748 XI11_3/XI0/XI0_26/d__5_ XI11_3/XI0/XI0_26/d_5_ DECAP_INV_G11
XG9749 XI11_3/XI0/XI0_26/d__4_ XI11_3/XI0/XI0_26/d_4_ DECAP_INV_G11
XG9750 XI11_3/XI0/XI0_26/d__3_ XI11_3/XI0/XI0_26/d_3_ DECAP_INV_G11
XG9751 XI11_3/XI0/XI0_26/d__2_ XI11_3/XI0/XI0_26/d_2_ DECAP_INV_G11
XG9752 XI11_3/XI0/XI0_26/d__1_ XI11_3/XI0/XI0_26/d_1_ DECAP_INV_G11
XG9753 XI11_3/XI0/XI0_26/d__0_ XI11_3/XI0/XI0_26/d_0_ DECAP_INV_G11
XG9754 XI11_3/XI0/XI0_26/d_15_ XI11_3/XI0/XI0_26/d__15_ DECAP_INV_G11
XG9755 XI11_3/XI0/XI0_26/d_14_ XI11_3/XI0/XI0_26/d__14_ DECAP_INV_G11
XG9756 XI11_3/XI0/XI0_26/d_13_ XI11_3/XI0/XI0_26/d__13_ DECAP_INV_G11
XG9757 XI11_3/XI0/XI0_26/d_12_ XI11_3/XI0/XI0_26/d__12_ DECAP_INV_G11
XG9758 XI11_3/XI0/XI0_26/d_11_ XI11_3/XI0/XI0_26/d__11_ DECAP_INV_G11
XG9759 XI11_3/XI0/XI0_26/d_10_ XI11_3/XI0/XI0_26/d__10_ DECAP_INV_G11
XG9760 XI11_3/XI0/XI0_26/d_9_ XI11_3/XI0/XI0_26/d__9_ DECAP_INV_G11
XG9761 XI11_3/XI0/XI0_26/d_8_ XI11_3/XI0/XI0_26/d__8_ DECAP_INV_G11
XG9762 XI11_3/XI0/XI0_26/d_7_ XI11_3/XI0/XI0_26/d__7_ DECAP_INV_G11
XG9763 XI11_3/XI0/XI0_26/d_6_ XI11_3/XI0/XI0_26/d__6_ DECAP_INV_G11
XG9764 XI11_3/XI0/XI0_26/d_5_ XI11_3/XI0/XI0_26/d__5_ DECAP_INV_G11
XG9765 XI11_3/XI0/XI0_26/d_4_ XI11_3/XI0/XI0_26/d__4_ DECAP_INV_G11
XG9766 XI11_3/XI0/XI0_26/d_3_ XI11_3/XI0/XI0_26/d__3_ DECAP_INV_G11
XG9767 XI11_3/XI0/XI0_26/d_2_ XI11_3/XI0/XI0_26/d__2_ DECAP_INV_G11
XG9768 XI11_3/XI0/XI0_26/d_1_ XI11_3/XI0/XI0_26/d__1_ DECAP_INV_G11
XG9769 XI11_3/XI0/XI0_26/d_0_ XI11_3/XI0/XI0_26/d__0_ DECAP_INV_G11
XG9770 XI11_3/XI0/XI0_25/d__15_ XI11_3/XI0/XI0_25/d_15_ DECAP_INV_G11
XG9771 XI11_3/XI0/XI0_25/d__14_ XI11_3/XI0/XI0_25/d_14_ DECAP_INV_G11
XG9772 XI11_3/XI0/XI0_25/d__13_ XI11_3/XI0/XI0_25/d_13_ DECAP_INV_G11
XG9773 XI11_3/XI0/XI0_25/d__12_ XI11_3/XI0/XI0_25/d_12_ DECAP_INV_G11
XG9774 XI11_3/XI0/XI0_25/d__11_ XI11_3/XI0/XI0_25/d_11_ DECAP_INV_G11
XG9775 XI11_3/XI0/XI0_25/d__10_ XI11_3/XI0/XI0_25/d_10_ DECAP_INV_G11
XG9776 XI11_3/XI0/XI0_25/d__9_ XI11_3/XI0/XI0_25/d_9_ DECAP_INV_G11
XG9777 XI11_3/XI0/XI0_25/d__8_ XI11_3/XI0/XI0_25/d_8_ DECAP_INV_G11
XG9778 XI11_3/XI0/XI0_25/d__7_ XI11_3/XI0/XI0_25/d_7_ DECAP_INV_G11
XG9779 XI11_3/XI0/XI0_25/d__6_ XI11_3/XI0/XI0_25/d_6_ DECAP_INV_G11
XG9780 XI11_3/XI0/XI0_25/d__5_ XI11_3/XI0/XI0_25/d_5_ DECAP_INV_G11
XG9781 XI11_3/XI0/XI0_25/d__4_ XI11_3/XI0/XI0_25/d_4_ DECAP_INV_G11
XG9782 XI11_3/XI0/XI0_25/d__3_ XI11_3/XI0/XI0_25/d_3_ DECAP_INV_G11
XG9783 XI11_3/XI0/XI0_25/d__2_ XI11_3/XI0/XI0_25/d_2_ DECAP_INV_G11
XG9784 XI11_3/XI0/XI0_25/d__1_ XI11_3/XI0/XI0_25/d_1_ DECAP_INV_G11
XG9785 XI11_3/XI0/XI0_25/d__0_ XI11_3/XI0/XI0_25/d_0_ DECAP_INV_G11
XG9786 XI11_3/XI0/XI0_25/d_15_ XI11_3/XI0/XI0_25/d__15_ DECAP_INV_G11
XG9787 XI11_3/XI0/XI0_25/d_14_ XI11_3/XI0/XI0_25/d__14_ DECAP_INV_G11
XG9788 XI11_3/XI0/XI0_25/d_13_ XI11_3/XI0/XI0_25/d__13_ DECAP_INV_G11
XG9789 XI11_3/XI0/XI0_25/d_12_ XI11_3/XI0/XI0_25/d__12_ DECAP_INV_G11
XG9790 XI11_3/XI0/XI0_25/d_11_ XI11_3/XI0/XI0_25/d__11_ DECAP_INV_G11
XG9791 XI11_3/XI0/XI0_25/d_10_ XI11_3/XI0/XI0_25/d__10_ DECAP_INV_G11
XG9792 XI11_3/XI0/XI0_25/d_9_ XI11_3/XI0/XI0_25/d__9_ DECAP_INV_G11
XG9793 XI11_3/XI0/XI0_25/d_8_ XI11_3/XI0/XI0_25/d__8_ DECAP_INV_G11
XG9794 XI11_3/XI0/XI0_25/d_7_ XI11_3/XI0/XI0_25/d__7_ DECAP_INV_G11
XG9795 XI11_3/XI0/XI0_25/d_6_ XI11_3/XI0/XI0_25/d__6_ DECAP_INV_G11
XG9796 XI11_3/XI0/XI0_25/d_5_ XI11_3/XI0/XI0_25/d__5_ DECAP_INV_G11
XG9797 XI11_3/XI0/XI0_25/d_4_ XI11_3/XI0/XI0_25/d__4_ DECAP_INV_G11
XG9798 XI11_3/XI0/XI0_25/d_3_ XI11_3/XI0/XI0_25/d__3_ DECAP_INV_G11
XG9799 XI11_3/XI0/XI0_25/d_2_ XI11_3/XI0/XI0_25/d__2_ DECAP_INV_G11
XG9800 XI11_3/XI0/XI0_25/d_1_ XI11_3/XI0/XI0_25/d__1_ DECAP_INV_G11
XG9801 XI11_3/XI0/XI0_25/d_0_ XI11_3/XI0/XI0_25/d__0_ DECAP_INV_G11
XG9802 XI11_3/XI0/XI0_24/d__15_ XI11_3/XI0/XI0_24/d_15_ DECAP_INV_G11
XG9803 XI11_3/XI0/XI0_24/d__14_ XI11_3/XI0/XI0_24/d_14_ DECAP_INV_G11
XG9804 XI11_3/XI0/XI0_24/d__13_ XI11_3/XI0/XI0_24/d_13_ DECAP_INV_G11
XG9805 XI11_3/XI0/XI0_24/d__12_ XI11_3/XI0/XI0_24/d_12_ DECAP_INV_G11
XG9806 XI11_3/XI0/XI0_24/d__11_ XI11_3/XI0/XI0_24/d_11_ DECAP_INV_G11
XG9807 XI11_3/XI0/XI0_24/d__10_ XI11_3/XI0/XI0_24/d_10_ DECAP_INV_G11
XG9808 XI11_3/XI0/XI0_24/d__9_ XI11_3/XI0/XI0_24/d_9_ DECAP_INV_G11
XG9809 XI11_3/XI0/XI0_24/d__8_ XI11_3/XI0/XI0_24/d_8_ DECAP_INV_G11
XG9810 XI11_3/XI0/XI0_24/d__7_ XI11_3/XI0/XI0_24/d_7_ DECAP_INV_G11
XG9811 XI11_3/XI0/XI0_24/d__6_ XI11_3/XI0/XI0_24/d_6_ DECAP_INV_G11
XG9812 XI11_3/XI0/XI0_24/d__5_ XI11_3/XI0/XI0_24/d_5_ DECAP_INV_G11
XG9813 XI11_3/XI0/XI0_24/d__4_ XI11_3/XI0/XI0_24/d_4_ DECAP_INV_G11
XG9814 XI11_3/XI0/XI0_24/d__3_ XI11_3/XI0/XI0_24/d_3_ DECAP_INV_G11
XG9815 XI11_3/XI0/XI0_24/d__2_ XI11_3/XI0/XI0_24/d_2_ DECAP_INV_G11
XG9816 XI11_3/XI0/XI0_24/d__1_ XI11_3/XI0/XI0_24/d_1_ DECAP_INV_G11
XG9817 XI11_3/XI0/XI0_24/d__0_ XI11_3/XI0/XI0_24/d_0_ DECAP_INV_G11
XG9818 XI11_3/XI0/XI0_24/d_15_ XI11_3/XI0/XI0_24/d__15_ DECAP_INV_G11
XG9819 XI11_3/XI0/XI0_24/d_14_ XI11_3/XI0/XI0_24/d__14_ DECAP_INV_G11
XG9820 XI11_3/XI0/XI0_24/d_13_ XI11_3/XI0/XI0_24/d__13_ DECAP_INV_G11
XG9821 XI11_3/XI0/XI0_24/d_12_ XI11_3/XI0/XI0_24/d__12_ DECAP_INV_G11
XG9822 XI11_3/XI0/XI0_24/d_11_ XI11_3/XI0/XI0_24/d__11_ DECAP_INV_G11
XG9823 XI11_3/XI0/XI0_24/d_10_ XI11_3/XI0/XI0_24/d__10_ DECAP_INV_G11
XG9824 XI11_3/XI0/XI0_24/d_9_ XI11_3/XI0/XI0_24/d__9_ DECAP_INV_G11
XG9825 XI11_3/XI0/XI0_24/d_8_ XI11_3/XI0/XI0_24/d__8_ DECAP_INV_G11
XG9826 XI11_3/XI0/XI0_24/d_7_ XI11_3/XI0/XI0_24/d__7_ DECAP_INV_G11
XG9827 XI11_3/XI0/XI0_24/d_6_ XI11_3/XI0/XI0_24/d__6_ DECAP_INV_G11
XG9828 XI11_3/XI0/XI0_24/d_5_ XI11_3/XI0/XI0_24/d__5_ DECAP_INV_G11
XG9829 XI11_3/XI0/XI0_24/d_4_ XI11_3/XI0/XI0_24/d__4_ DECAP_INV_G11
XG9830 XI11_3/XI0/XI0_24/d_3_ XI11_3/XI0/XI0_24/d__3_ DECAP_INV_G11
XG9831 XI11_3/XI0/XI0_24/d_2_ XI11_3/XI0/XI0_24/d__2_ DECAP_INV_G11
XG9832 XI11_3/XI0/XI0_24/d_1_ XI11_3/XI0/XI0_24/d__1_ DECAP_INV_G11
XG9833 XI11_3/XI0/XI0_24/d_0_ XI11_3/XI0/XI0_24/d__0_ DECAP_INV_G11
XG9834 XI11_3/XI0/XI0_23/d__15_ XI11_3/XI0/XI0_23/d_15_ DECAP_INV_G11
XG9835 XI11_3/XI0/XI0_23/d__14_ XI11_3/XI0/XI0_23/d_14_ DECAP_INV_G11
XG9836 XI11_3/XI0/XI0_23/d__13_ XI11_3/XI0/XI0_23/d_13_ DECAP_INV_G11
XG9837 XI11_3/XI0/XI0_23/d__12_ XI11_3/XI0/XI0_23/d_12_ DECAP_INV_G11
XG9838 XI11_3/XI0/XI0_23/d__11_ XI11_3/XI0/XI0_23/d_11_ DECAP_INV_G11
XG9839 XI11_3/XI0/XI0_23/d__10_ XI11_3/XI0/XI0_23/d_10_ DECAP_INV_G11
XG9840 XI11_3/XI0/XI0_23/d__9_ XI11_3/XI0/XI0_23/d_9_ DECAP_INV_G11
XG9841 XI11_3/XI0/XI0_23/d__8_ XI11_3/XI0/XI0_23/d_8_ DECAP_INV_G11
XG9842 XI11_3/XI0/XI0_23/d__7_ XI11_3/XI0/XI0_23/d_7_ DECAP_INV_G11
XG9843 XI11_3/XI0/XI0_23/d__6_ XI11_3/XI0/XI0_23/d_6_ DECAP_INV_G11
XG9844 XI11_3/XI0/XI0_23/d__5_ XI11_3/XI0/XI0_23/d_5_ DECAP_INV_G11
XG9845 XI11_3/XI0/XI0_23/d__4_ XI11_3/XI0/XI0_23/d_4_ DECAP_INV_G11
XG9846 XI11_3/XI0/XI0_23/d__3_ XI11_3/XI0/XI0_23/d_3_ DECAP_INV_G11
XG9847 XI11_3/XI0/XI0_23/d__2_ XI11_3/XI0/XI0_23/d_2_ DECAP_INV_G11
XG9848 XI11_3/XI0/XI0_23/d__1_ XI11_3/XI0/XI0_23/d_1_ DECAP_INV_G11
XG9849 XI11_3/XI0/XI0_23/d__0_ XI11_3/XI0/XI0_23/d_0_ DECAP_INV_G11
XG9850 XI11_3/XI0/XI0_23/d_15_ XI11_3/XI0/XI0_23/d__15_ DECAP_INV_G11
XG9851 XI11_3/XI0/XI0_23/d_14_ XI11_3/XI0/XI0_23/d__14_ DECAP_INV_G11
XG9852 XI11_3/XI0/XI0_23/d_13_ XI11_3/XI0/XI0_23/d__13_ DECAP_INV_G11
XG9853 XI11_3/XI0/XI0_23/d_12_ XI11_3/XI0/XI0_23/d__12_ DECAP_INV_G11
XG9854 XI11_3/XI0/XI0_23/d_11_ XI11_3/XI0/XI0_23/d__11_ DECAP_INV_G11
XG9855 XI11_3/XI0/XI0_23/d_10_ XI11_3/XI0/XI0_23/d__10_ DECAP_INV_G11
XG9856 XI11_3/XI0/XI0_23/d_9_ XI11_3/XI0/XI0_23/d__9_ DECAP_INV_G11
XG9857 XI11_3/XI0/XI0_23/d_8_ XI11_3/XI0/XI0_23/d__8_ DECAP_INV_G11
XG9858 XI11_3/XI0/XI0_23/d_7_ XI11_3/XI0/XI0_23/d__7_ DECAP_INV_G11
XG9859 XI11_3/XI0/XI0_23/d_6_ XI11_3/XI0/XI0_23/d__6_ DECAP_INV_G11
XG9860 XI11_3/XI0/XI0_23/d_5_ XI11_3/XI0/XI0_23/d__5_ DECAP_INV_G11
XG9861 XI11_3/XI0/XI0_23/d_4_ XI11_3/XI0/XI0_23/d__4_ DECAP_INV_G11
XG9862 XI11_3/XI0/XI0_23/d_3_ XI11_3/XI0/XI0_23/d__3_ DECAP_INV_G11
XG9863 XI11_3/XI0/XI0_23/d_2_ XI11_3/XI0/XI0_23/d__2_ DECAP_INV_G11
XG9864 XI11_3/XI0/XI0_23/d_1_ XI11_3/XI0/XI0_23/d__1_ DECAP_INV_G11
XG9865 XI11_3/XI0/XI0_23/d_0_ XI11_3/XI0/XI0_23/d__0_ DECAP_INV_G11
XG9866 XI11_3/XI0/XI0_22/d__15_ XI11_3/XI0/XI0_22/d_15_ DECAP_INV_G11
XG9867 XI11_3/XI0/XI0_22/d__14_ XI11_3/XI0/XI0_22/d_14_ DECAP_INV_G11
XG9868 XI11_3/XI0/XI0_22/d__13_ XI11_3/XI0/XI0_22/d_13_ DECAP_INV_G11
XG9869 XI11_3/XI0/XI0_22/d__12_ XI11_3/XI0/XI0_22/d_12_ DECAP_INV_G11
XG9870 XI11_3/XI0/XI0_22/d__11_ XI11_3/XI0/XI0_22/d_11_ DECAP_INV_G11
XG9871 XI11_3/XI0/XI0_22/d__10_ XI11_3/XI0/XI0_22/d_10_ DECAP_INV_G11
XG9872 XI11_3/XI0/XI0_22/d__9_ XI11_3/XI0/XI0_22/d_9_ DECAP_INV_G11
XG9873 XI11_3/XI0/XI0_22/d__8_ XI11_3/XI0/XI0_22/d_8_ DECAP_INV_G11
XG9874 XI11_3/XI0/XI0_22/d__7_ XI11_3/XI0/XI0_22/d_7_ DECAP_INV_G11
XG9875 XI11_3/XI0/XI0_22/d__6_ XI11_3/XI0/XI0_22/d_6_ DECAP_INV_G11
XG9876 XI11_3/XI0/XI0_22/d__5_ XI11_3/XI0/XI0_22/d_5_ DECAP_INV_G11
XG9877 XI11_3/XI0/XI0_22/d__4_ XI11_3/XI0/XI0_22/d_4_ DECAP_INV_G11
XG9878 XI11_3/XI0/XI0_22/d__3_ XI11_3/XI0/XI0_22/d_3_ DECAP_INV_G11
XG9879 XI11_3/XI0/XI0_22/d__2_ XI11_3/XI0/XI0_22/d_2_ DECAP_INV_G11
XG9880 XI11_3/XI0/XI0_22/d__1_ XI11_3/XI0/XI0_22/d_1_ DECAP_INV_G11
XG9881 XI11_3/XI0/XI0_22/d__0_ XI11_3/XI0/XI0_22/d_0_ DECAP_INV_G11
XG9882 XI11_3/XI0/XI0_22/d_15_ XI11_3/XI0/XI0_22/d__15_ DECAP_INV_G11
XG9883 XI11_3/XI0/XI0_22/d_14_ XI11_3/XI0/XI0_22/d__14_ DECAP_INV_G11
XG9884 XI11_3/XI0/XI0_22/d_13_ XI11_3/XI0/XI0_22/d__13_ DECAP_INV_G11
XG9885 XI11_3/XI0/XI0_22/d_12_ XI11_3/XI0/XI0_22/d__12_ DECAP_INV_G11
XG9886 XI11_3/XI0/XI0_22/d_11_ XI11_3/XI0/XI0_22/d__11_ DECAP_INV_G11
XG9887 XI11_3/XI0/XI0_22/d_10_ XI11_3/XI0/XI0_22/d__10_ DECAP_INV_G11
XG9888 XI11_3/XI0/XI0_22/d_9_ XI11_3/XI0/XI0_22/d__9_ DECAP_INV_G11
XG9889 XI11_3/XI0/XI0_22/d_8_ XI11_3/XI0/XI0_22/d__8_ DECAP_INV_G11
XG9890 XI11_3/XI0/XI0_22/d_7_ XI11_3/XI0/XI0_22/d__7_ DECAP_INV_G11
XG9891 XI11_3/XI0/XI0_22/d_6_ XI11_3/XI0/XI0_22/d__6_ DECAP_INV_G11
XG9892 XI11_3/XI0/XI0_22/d_5_ XI11_3/XI0/XI0_22/d__5_ DECAP_INV_G11
XG9893 XI11_3/XI0/XI0_22/d_4_ XI11_3/XI0/XI0_22/d__4_ DECAP_INV_G11
XG9894 XI11_3/XI0/XI0_22/d_3_ XI11_3/XI0/XI0_22/d__3_ DECAP_INV_G11
XG9895 XI11_3/XI0/XI0_22/d_2_ XI11_3/XI0/XI0_22/d__2_ DECAP_INV_G11
XG9896 XI11_3/XI0/XI0_22/d_1_ XI11_3/XI0/XI0_22/d__1_ DECAP_INV_G11
XG9897 XI11_3/XI0/XI0_22/d_0_ XI11_3/XI0/XI0_22/d__0_ DECAP_INV_G11
XG9898 XI11_3/XI0/XI0_21/d__15_ XI11_3/XI0/XI0_21/d_15_ DECAP_INV_G11
XG9899 XI11_3/XI0/XI0_21/d__14_ XI11_3/XI0/XI0_21/d_14_ DECAP_INV_G11
XG9900 XI11_3/XI0/XI0_21/d__13_ XI11_3/XI0/XI0_21/d_13_ DECAP_INV_G11
XG9901 XI11_3/XI0/XI0_21/d__12_ XI11_3/XI0/XI0_21/d_12_ DECAP_INV_G11
XG9902 XI11_3/XI0/XI0_21/d__11_ XI11_3/XI0/XI0_21/d_11_ DECAP_INV_G11
XG9903 XI11_3/XI0/XI0_21/d__10_ XI11_3/XI0/XI0_21/d_10_ DECAP_INV_G11
XG9904 XI11_3/XI0/XI0_21/d__9_ XI11_3/XI0/XI0_21/d_9_ DECAP_INV_G11
XG9905 XI11_3/XI0/XI0_21/d__8_ XI11_3/XI0/XI0_21/d_8_ DECAP_INV_G11
XG9906 XI11_3/XI0/XI0_21/d__7_ XI11_3/XI0/XI0_21/d_7_ DECAP_INV_G11
XG9907 XI11_3/XI0/XI0_21/d__6_ XI11_3/XI0/XI0_21/d_6_ DECAP_INV_G11
XG9908 XI11_3/XI0/XI0_21/d__5_ XI11_3/XI0/XI0_21/d_5_ DECAP_INV_G11
XG9909 XI11_3/XI0/XI0_21/d__4_ XI11_3/XI0/XI0_21/d_4_ DECAP_INV_G11
XG9910 XI11_3/XI0/XI0_21/d__3_ XI11_3/XI0/XI0_21/d_3_ DECAP_INV_G11
XG9911 XI11_3/XI0/XI0_21/d__2_ XI11_3/XI0/XI0_21/d_2_ DECAP_INV_G11
XG9912 XI11_3/XI0/XI0_21/d__1_ XI11_3/XI0/XI0_21/d_1_ DECAP_INV_G11
XG9913 XI11_3/XI0/XI0_21/d__0_ XI11_3/XI0/XI0_21/d_0_ DECAP_INV_G11
XG9914 XI11_3/XI0/XI0_21/d_15_ XI11_3/XI0/XI0_21/d__15_ DECAP_INV_G11
XG9915 XI11_3/XI0/XI0_21/d_14_ XI11_3/XI0/XI0_21/d__14_ DECAP_INV_G11
XG9916 XI11_3/XI0/XI0_21/d_13_ XI11_3/XI0/XI0_21/d__13_ DECAP_INV_G11
XG9917 XI11_3/XI0/XI0_21/d_12_ XI11_3/XI0/XI0_21/d__12_ DECAP_INV_G11
XG9918 XI11_3/XI0/XI0_21/d_11_ XI11_3/XI0/XI0_21/d__11_ DECAP_INV_G11
XG9919 XI11_3/XI0/XI0_21/d_10_ XI11_3/XI0/XI0_21/d__10_ DECAP_INV_G11
XG9920 XI11_3/XI0/XI0_21/d_9_ XI11_3/XI0/XI0_21/d__9_ DECAP_INV_G11
XG9921 XI11_3/XI0/XI0_21/d_8_ XI11_3/XI0/XI0_21/d__8_ DECAP_INV_G11
XG9922 XI11_3/XI0/XI0_21/d_7_ XI11_3/XI0/XI0_21/d__7_ DECAP_INV_G11
XG9923 XI11_3/XI0/XI0_21/d_6_ XI11_3/XI0/XI0_21/d__6_ DECAP_INV_G11
XG9924 XI11_3/XI0/XI0_21/d_5_ XI11_3/XI0/XI0_21/d__5_ DECAP_INV_G11
XG9925 XI11_3/XI0/XI0_21/d_4_ XI11_3/XI0/XI0_21/d__4_ DECAP_INV_G11
XG9926 XI11_3/XI0/XI0_21/d_3_ XI11_3/XI0/XI0_21/d__3_ DECAP_INV_G11
XG9927 XI11_3/XI0/XI0_21/d_2_ XI11_3/XI0/XI0_21/d__2_ DECAP_INV_G11
XG9928 XI11_3/XI0/XI0_21/d_1_ XI11_3/XI0/XI0_21/d__1_ DECAP_INV_G11
XG9929 XI11_3/XI0/XI0_21/d_0_ XI11_3/XI0/XI0_21/d__0_ DECAP_INV_G11
XG9930 XI11_3/XI0/XI0_20/d__15_ XI11_3/XI0/XI0_20/d_15_ DECAP_INV_G11
XG9931 XI11_3/XI0/XI0_20/d__14_ XI11_3/XI0/XI0_20/d_14_ DECAP_INV_G11
XG9932 XI11_3/XI0/XI0_20/d__13_ XI11_3/XI0/XI0_20/d_13_ DECAP_INV_G11
XG9933 XI11_3/XI0/XI0_20/d__12_ XI11_3/XI0/XI0_20/d_12_ DECAP_INV_G11
XG9934 XI11_3/XI0/XI0_20/d__11_ XI11_3/XI0/XI0_20/d_11_ DECAP_INV_G11
XG9935 XI11_3/XI0/XI0_20/d__10_ XI11_3/XI0/XI0_20/d_10_ DECAP_INV_G11
XG9936 XI11_3/XI0/XI0_20/d__9_ XI11_3/XI0/XI0_20/d_9_ DECAP_INV_G11
XG9937 XI11_3/XI0/XI0_20/d__8_ XI11_3/XI0/XI0_20/d_8_ DECAP_INV_G11
XG9938 XI11_3/XI0/XI0_20/d__7_ XI11_3/XI0/XI0_20/d_7_ DECAP_INV_G11
XG9939 XI11_3/XI0/XI0_20/d__6_ XI11_3/XI0/XI0_20/d_6_ DECAP_INV_G11
XG9940 XI11_3/XI0/XI0_20/d__5_ XI11_3/XI0/XI0_20/d_5_ DECAP_INV_G11
XG9941 XI11_3/XI0/XI0_20/d__4_ XI11_3/XI0/XI0_20/d_4_ DECAP_INV_G11
XG9942 XI11_3/XI0/XI0_20/d__3_ XI11_3/XI0/XI0_20/d_3_ DECAP_INV_G11
XG9943 XI11_3/XI0/XI0_20/d__2_ XI11_3/XI0/XI0_20/d_2_ DECAP_INV_G11
XG9944 XI11_3/XI0/XI0_20/d__1_ XI11_3/XI0/XI0_20/d_1_ DECAP_INV_G11
XG9945 XI11_3/XI0/XI0_20/d__0_ XI11_3/XI0/XI0_20/d_0_ DECAP_INV_G11
XG9946 XI11_3/XI0/XI0_20/d_15_ XI11_3/XI0/XI0_20/d__15_ DECAP_INV_G11
XG9947 XI11_3/XI0/XI0_20/d_14_ XI11_3/XI0/XI0_20/d__14_ DECAP_INV_G11
XG9948 XI11_3/XI0/XI0_20/d_13_ XI11_3/XI0/XI0_20/d__13_ DECAP_INV_G11
XG9949 XI11_3/XI0/XI0_20/d_12_ XI11_3/XI0/XI0_20/d__12_ DECAP_INV_G11
XG9950 XI11_3/XI0/XI0_20/d_11_ XI11_3/XI0/XI0_20/d__11_ DECAP_INV_G11
XG9951 XI11_3/XI0/XI0_20/d_10_ XI11_3/XI0/XI0_20/d__10_ DECAP_INV_G11
XG9952 XI11_3/XI0/XI0_20/d_9_ XI11_3/XI0/XI0_20/d__9_ DECAP_INV_G11
XG9953 XI11_3/XI0/XI0_20/d_8_ XI11_3/XI0/XI0_20/d__8_ DECAP_INV_G11
XG9954 XI11_3/XI0/XI0_20/d_7_ XI11_3/XI0/XI0_20/d__7_ DECAP_INV_G11
XG9955 XI11_3/XI0/XI0_20/d_6_ XI11_3/XI0/XI0_20/d__6_ DECAP_INV_G11
XG9956 XI11_3/XI0/XI0_20/d_5_ XI11_3/XI0/XI0_20/d__5_ DECAP_INV_G11
XG9957 XI11_3/XI0/XI0_20/d_4_ XI11_3/XI0/XI0_20/d__4_ DECAP_INV_G11
XG9958 XI11_3/XI0/XI0_20/d_3_ XI11_3/XI0/XI0_20/d__3_ DECAP_INV_G11
XG9959 XI11_3/XI0/XI0_20/d_2_ XI11_3/XI0/XI0_20/d__2_ DECAP_INV_G11
XG9960 XI11_3/XI0/XI0_20/d_1_ XI11_3/XI0/XI0_20/d__1_ DECAP_INV_G11
XG9961 XI11_3/XI0/XI0_20/d_0_ XI11_3/XI0/XI0_20/d__0_ DECAP_INV_G11
XG9962 XI11_3/XI0/XI0_19/d__15_ XI11_3/XI0/XI0_19/d_15_ DECAP_INV_G11
XG9963 XI11_3/XI0/XI0_19/d__14_ XI11_3/XI0/XI0_19/d_14_ DECAP_INV_G11
XG9964 XI11_3/XI0/XI0_19/d__13_ XI11_3/XI0/XI0_19/d_13_ DECAP_INV_G11
XG9965 XI11_3/XI0/XI0_19/d__12_ XI11_3/XI0/XI0_19/d_12_ DECAP_INV_G11
XG9966 XI11_3/XI0/XI0_19/d__11_ XI11_3/XI0/XI0_19/d_11_ DECAP_INV_G11
XG9967 XI11_3/XI0/XI0_19/d__10_ XI11_3/XI0/XI0_19/d_10_ DECAP_INV_G11
XG9968 XI11_3/XI0/XI0_19/d__9_ XI11_3/XI0/XI0_19/d_9_ DECAP_INV_G11
XG9969 XI11_3/XI0/XI0_19/d__8_ XI11_3/XI0/XI0_19/d_8_ DECAP_INV_G11
XG9970 XI11_3/XI0/XI0_19/d__7_ XI11_3/XI0/XI0_19/d_7_ DECAP_INV_G11
XG9971 XI11_3/XI0/XI0_19/d__6_ XI11_3/XI0/XI0_19/d_6_ DECAP_INV_G11
XG9972 XI11_3/XI0/XI0_19/d__5_ XI11_3/XI0/XI0_19/d_5_ DECAP_INV_G11
XG9973 XI11_3/XI0/XI0_19/d__4_ XI11_3/XI0/XI0_19/d_4_ DECAP_INV_G11
XG9974 XI11_3/XI0/XI0_19/d__3_ XI11_3/XI0/XI0_19/d_3_ DECAP_INV_G11
XG9975 XI11_3/XI0/XI0_19/d__2_ XI11_3/XI0/XI0_19/d_2_ DECAP_INV_G11
XG9976 XI11_3/XI0/XI0_19/d__1_ XI11_3/XI0/XI0_19/d_1_ DECAP_INV_G11
XG9977 XI11_3/XI0/XI0_19/d__0_ XI11_3/XI0/XI0_19/d_0_ DECAP_INV_G11
XG9978 XI11_3/XI0/XI0_19/d_15_ XI11_3/XI0/XI0_19/d__15_ DECAP_INV_G11
XG9979 XI11_3/XI0/XI0_19/d_14_ XI11_3/XI0/XI0_19/d__14_ DECAP_INV_G11
XG9980 XI11_3/XI0/XI0_19/d_13_ XI11_3/XI0/XI0_19/d__13_ DECAP_INV_G11
XG9981 XI11_3/XI0/XI0_19/d_12_ XI11_3/XI0/XI0_19/d__12_ DECAP_INV_G11
XG9982 XI11_3/XI0/XI0_19/d_11_ XI11_3/XI0/XI0_19/d__11_ DECAP_INV_G11
XG9983 XI11_3/XI0/XI0_19/d_10_ XI11_3/XI0/XI0_19/d__10_ DECAP_INV_G11
XG9984 XI11_3/XI0/XI0_19/d_9_ XI11_3/XI0/XI0_19/d__9_ DECAP_INV_G11
XG9985 XI11_3/XI0/XI0_19/d_8_ XI11_3/XI0/XI0_19/d__8_ DECAP_INV_G11
XG9986 XI11_3/XI0/XI0_19/d_7_ XI11_3/XI0/XI0_19/d__7_ DECAP_INV_G11
XG9987 XI11_3/XI0/XI0_19/d_6_ XI11_3/XI0/XI0_19/d__6_ DECAP_INV_G11
XG9988 XI11_3/XI0/XI0_19/d_5_ XI11_3/XI0/XI0_19/d__5_ DECAP_INV_G11
XG9989 XI11_3/XI0/XI0_19/d_4_ XI11_3/XI0/XI0_19/d__4_ DECAP_INV_G11
XG9990 XI11_3/XI0/XI0_19/d_3_ XI11_3/XI0/XI0_19/d__3_ DECAP_INV_G11
XG9991 XI11_3/XI0/XI0_19/d_2_ XI11_3/XI0/XI0_19/d__2_ DECAP_INV_G11
XG9992 XI11_3/XI0/XI0_19/d_1_ XI11_3/XI0/XI0_19/d__1_ DECAP_INV_G11
XG9993 XI11_3/XI0/XI0_19/d_0_ XI11_3/XI0/XI0_19/d__0_ DECAP_INV_G11
XG9994 XI11_3/XI0/XI0_18/d__15_ XI11_3/XI0/XI0_18/d_15_ DECAP_INV_G11
XG9995 XI11_3/XI0/XI0_18/d__14_ XI11_3/XI0/XI0_18/d_14_ DECAP_INV_G11
XG9996 XI11_3/XI0/XI0_18/d__13_ XI11_3/XI0/XI0_18/d_13_ DECAP_INV_G11
XG9997 XI11_3/XI0/XI0_18/d__12_ XI11_3/XI0/XI0_18/d_12_ DECAP_INV_G11
XG9998 XI11_3/XI0/XI0_18/d__11_ XI11_3/XI0/XI0_18/d_11_ DECAP_INV_G11
XG9999 XI11_3/XI0/XI0_18/d__10_ XI11_3/XI0/XI0_18/d_10_ DECAP_INV_G11
XG10000 XI11_3/XI0/XI0_18/d__9_ XI11_3/XI0/XI0_18/d_9_ DECAP_INV_G11
XG10001 XI11_3/XI0/XI0_18/d__8_ XI11_3/XI0/XI0_18/d_8_ DECAP_INV_G11
XG10002 XI11_3/XI0/XI0_18/d__7_ XI11_3/XI0/XI0_18/d_7_ DECAP_INV_G11
XG10003 XI11_3/XI0/XI0_18/d__6_ XI11_3/XI0/XI0_18/d_6_ DECAP_INV_G11
XG10004 XI11_3/XI0/XI0_18/d__5_ XI11_3/XI0/XI0_18/d_5_ DECAP_INV_G11
XG10005 XI11_3/XI0/XI0_18/d__4_ XI11_3/XI0/XI0_18/d_4_ DECAP_INV_G11
XG10006 XI11_3/XI0/XI0_18/d__3_ XI11_3/XI0/XI0_18/d_3_ DECAP_INV_G11
XG10007 XI11_3/XI0/XI0_18/d__2_ XI11_3/XI0/XI0_18/d_2_ DECAP_INV_G11
XG10008 XI11_3/XI0/XI0_18/d__1_ XI11_3/XI0/XI0_18/d_1_ DECAP_INV_G11
XG10009 XI11_3/XI0/XI0_18/d__0_ XI11_3/XI0/XI0_18/d_0_ DECAP_INV_G11
XG10010 XI11_3/XI0/XI0_18/d_15_ XI11_3/XI0/XI0_18/d__15_ DECAP_INV_G11
XG10011 XI11_3/XI0/XI0_18/d_14_ XI11_3/XI0/XI0_18/d__14_ DECAP_INV_G11
XG10012 XI11_3/XI0/XI0_18/d_13_ XI11_3/XI0/XI0_18/d__13_ DECAP_INV_G11
XG10013 XI11_3/XI0/XI0_18/d_12_ XI11_3/XI0/XI0_18/d__12_ DECAP_INV_G11
XG10014 XI11_3/XI0/XI0_18/d_11_ XI11_3/XI0/XI0_18/d__11_ DECAP_INV_G11
XG10015 XI11_3/XI0/XI0_18/d_10_ XI11_3/XI0/XI0_18/d__10_ DECAP_INV_G11
XG10016 XI11_3/XI0/XI0_18/d_9_ XI11_3/XI0/XI0_18/d__9_ DECAP_INV_G11
XG10017 XI11_3/XI0/XI0_18/d_8_ XI11_3/XI0/XI0_18/d__8_ DECAP_INV_G11
XG10018 XI11_3/XI0/XI0_18/d_7_ XI11_3/XI0/XI0_18/d__7_ DECAP_INV_G11
XG10019 XI11_3/XI0/XI0_18/d_6_ XI11_3/XI0/XI0_18/d__6_ DECAP_INV_G11
XG10020 XI11_3/XI0/XI0_18/d_5_ XI11_3/XI0/XI0_18/d__5_ DECAP_INV_G11
XG10021 XI11_3/XI0/XI0_18/d_4_ XI11_3/XI0/XI0_18/d__4_ DECAP_INV_G11
XG10022 XI11_3/XI0/XI0_18/d_3_ XI11_3/XI0/XI0_18/d__3_ DECAP_INV_G11
XG10023 XI11_3/XI0/XI0_18/d_2_ XI11_3/XI0/XI0_18/d__2_ DECAP_INV_G11
XG10024 XI11_3/XI0/XI0_18/d_1_ XI11_3/XI0/XI0_18/d__1_ DECAP_INV_G11
XG10025 XI11_3/XI0/XI0_18/d_0_ XI11_3/XI0/XI0_18/d__0_ DECAP_INV_G11
XG10026 XI11_3/XI0/XI0_17/d__15_ XI11_3/XI0/XI0_17/d_15_ DECAP_INV_G11
XG10027 XI11_3/XI0/XI0_17/d__14_ XI11_3/XI0/XI0_17/d_14_ DECAP_INV_G11
XG10028 XI11_3/XI0/XI0_17/d__13_ XI11_3/XI0/XI0_17/d_13_ DECAP_INV_G11
XG10029 XI11_3/XI0/XI0_17/d__12_ XI11_3/XI0/XI0_17/d_12_ DECAP_INV_G11
XG10030 XI11_3/XI0/XI0_17/d__11_ XI11_3/XI0/XI0_17/d_11_ DECAP_INV_G11
XG10031 XI11_3/XI0/XI0_17/d__10_ XI11_3/XI0/XI0_17/d_10_ DECAP_INV_G11
XG10032 XI11_3/XI0/XI0_17/d__9_ XI11_3/XI0/XI0_17/d_9_ DECAP_INV_G11
XG10033 XI11_3/XI0/XI0_17/d__8_ XI11_3/XI0/XI0_17/d_8_ DECAP_INV_G11
XG10034 XI11_3/XI0/XI0_17/d__7_ XI11_3/XI0/XI0_17/d_7_ DECAP_INV_G11
XG10035 XI11_3/XI0/XI0_17/d__6_ XI11_3/XI0/XI0_17/d_6_ DECAP_INV_G11
XG10036 XI11_3/XI0/XI0_17/d__5_ XI11_3/XI0/XI0_17/d_5_ DECAP_INV_G11
XG10037 XI11_3/XI0/XI0_17/d__4_ XI11_3/XI0/XI0_17/d_4_ DECAP_INV_G11
XG10038 XI11_3/XI0/XI0_17/d__3_ XI11_3/XI0/XI0_17/d_3_ DECAP_INV_G11
XG10039 XI11_3/XI0/XI0_17/d__2_ XI11_3/XI0/XI0_17/d_2_ DECAP_INV_G11
XG10040 XI11_3/XI0/XI0_17/d__1_ XI11_3/XI0/XI0_17/d_1_ DECAP_INV_G11
XG10041 XI11_3/XI0/XI0_17/d__0_ XI11_3/XI0/XI0_17/d_0_ DECAP_INV_G11
XG10042 XI11_3/XI0/XI0_17/d_15_ XI11_3/XI0/XI0_17/d__15_ DECAP_INV_G11
XG10043 XI11_3/XI0/XI0_17/d_14_ XI11_3/XI0/XI0_17/d__14_ DECAP_INV_G11
XG10044 XI11_3/XI0/XI0_17/d_13_ XI11_3/XI0/XI0_17/d__13_ DECAP_INV_G11
XG10045 XI11_3/XI0/XI0_17/d_12_ XI11_3/XI0/XI0_17/d__12_ DECAP_INV_G11
XG10046 XI11_3/XI0/XI0_17/d_11_ XI11_3/XI0/XI0_17/d__11_ DECAP_INV_G11
XG10047 XI11_3/XI0/XI0_17/d_10_ XI11_3/XI0/XI0_17/d__10_ DECAP_INV_G11
XG10048 XI11_3/XI0/XI0_17/d_9_ XI11_3/XI0/XI0_17/d__9_ DECAP_INV_G11
XG10049 XI11_3/XI0/XI0_17/d_8_ XI11_3/XI0/XI0_17/d__8_ DECAP_INV_G11
XG10050 XI11_3/XI0/XI0_17/d_7_ XI11_3/XI0/XI0_17/d__7_ DECAP_INV_G11
XG10051 XI11_3/XI0/XI0_17/d_6_ XI11_3/XI0/XI0_17/d__6_ DECAP_INV_G11
XG10052 XI11_3/XI0/XI0_17/d_5_ XI11_3/XI0/XI0_17/d__5_ DECAP_INV_G11
XG10053 XI11_3/XI0/XI0_17/d_4_ XI11_3/XI0/XI0_17/d__4_ DECAP_INV_G11
XG10054 XI11_3/XI0/XI0_17/d_3_ XI11_3/XI0/XI0_17/d__3_ DECAP_INV_G11
XG10055 XI11_3/XI0/XI0_17/d_2_ XI11_3/XI0/XI0_17/d__2_ DECAP_INV_G11
XG10056 XI11_3/XI0/XI0_17/d_1_ XI11_3/XI0/XI0_17/d__1_ DECAP_INV_G11
XG10057 XI11_3/XI0/XI0_17/d_0_ XI11_3/XI0/XI0_17/d__0_ DECAP_INV_G11
XG10058 XI11_3/XI0/XI0_16/d__15_ XI11_3/XI0/XI0_16/d_15_ DECAP_INV_G11
XG10059 XI11_3/XI0/XI0_16/d__14_ XI11_3/XI0/XI0_16/d_14_ DECAP_INV_G11
XG10060 XI11_3/XI0/XI0_16/d__13_ XI11_3/XI0/XI0_16/d_13_ DECAP_INV_G11
XG10061 XI11_3/XI0/XI0_16/d__12_ XI11_3/XI0/XI0_16/d_12_ DECAP_INV_G11
XG10062 XI11_3/XI0/XI0_16/d__11_ XI11_3/XI0/XI0_16/d_11_ DECAP_INV_G11
XG10063 XI11_3/XI0/XI0_16/d__10_ XI11_3/XI0/XI0_16/d_10_ DECAP_INV_G11
XG10064 XI11_3/XI0/XI0_16/d__9_ XI11_3/XI0/XI0_16/d_9_ DECAP_INV_G11
XG10065 XI11_3/XI0/XI0_16/d__8_ XI11_3/XI0/XI0_16/d_8_ DECAP_INV_G11
XG10066 XI11_3/XI0/XI0_16/d__7_ XI11_3/XI0/XI0_16/d_7_ DECAP_INV_G11
XG10067 XI11_3/XI0/XI0_16/d__6_ XI11_3/XI0/XI0_16/d_6_ DECAP_INV_G11
XG10068 XI11_3/XI0/XI0_16/d__5_ XI11_3/XI0/XI0_16/d_5_ DECAP_INV_G11
XG10069 XI11_3/XI0/XI0_16/d__4_ XI11_3/XI0/XI0_16/d_4_ DECAP_INV_G11
XG10070 XI11_3/XI0/XI0_16/d__3_ XI11_3/XI0/XI0_16/d_3_ DECAP_INV_G11
XG10071 XI11_3/XI0/XI0_16/d__2_ XI11_3/XI0/XI0_16/d_2_ DECAP_INV_G11
XG10072 XI11_3/XI0/XI0_16/d__1_ XI11_3/XI0/XI0_16/d_1_ DECAP_INV_G11
XG10073 XI11_3/XI0/XI0_16/d__0_ XI11_3/XI0/XI0_16/d_0_ DECAP_INV_G11
XG10074 XI11_3/XI0/XI0_16/d_15_ XI11_3/XI0/XI0_16/d__15_ DECAP_INV_G11
XG10075 XI11_3/XI0/XI0_16/d_14_ XI11_3/XI0/XI0_16/d__14_ DECAP_INV_G11
XG10076 XI11_3/XI0/XI0_16/d_13_ XI11_3/XI0/XI0_16/d__13_ DECAP_INV_G11
XG10077 XI11_3/XI0/XI0_16/d_12_ XI11_3/XI0/XI0_16/d__12_ DECAP_INV_G11
XG10078 XI11_3/XI0/XI0_16/d_11_ XI11_3/XI0/XI0_16/d__11_ DECAP_INV_G11
XG10079 XI11_3/XI0/XI0_16/d_10_ XI11_3/XI0/XI0_16/d__10_ DECAP_INV_G11
XG10080 XI11_3/XI0/XI0_16/d_9_ XI11_3/XI0/XI0_16/d__9_ DECAP_INV_G11
XG10081 XI11_3/XI0/XI0_16/d_8_ XI11_3/XI0/XI0_16/d__8_ DECAP_INV_G11
XG10082 XI11_3/XI0/XI0_16/d_7_ XI11_3/XI0/XI0_16/d__7_ DECAP_INV_G11
XG10083 XI11_3/XI0/XI0_16/d_6_ XI11_3/XI0/XI0_16/d__6_ DECAP_INV_G11
XG10084 XI11_3/XI0/XI0_16/d_5_ XI11_3/XI0/XI0_16/d__5_ DECAP_INV_G11
XG10085 XI11_3/XI0/XI0_16/d_4_ XI11_3/XI0/XI0_16/d__4_ DECAP_INV_G11
XG10086 XI11_3/XI0/XI0_16/d_3_ XI11_3/XI0/XI0_16/d__3_ DECAP_INV_G11
XG10087 XI11_3/XI0/XI0_16/d_2_ XI11_3/XI0/XI0_16/d__2_ DECAP_INV_G11
XG10088 XI11_3/XI0/XI0_16/d_1_ XI11_3/XI0/XI0_16/d__1_ DECAP_INV_G11
XG10089 XI11_3/XI0/XI0_16/d_0_ XI11_3/XI0/XI0_16/d__0_ DECAP_INV_G11
XG10090 XI11_3/XI0/XI0_15/d__15_ XI11_3/XI0/XI0_15/d_15_ DECAP_INV_G11
XG10091 XI11_3/XI0/XI0_15/d__14_ XI11_3/XI0/XI0_15/d_14_ DECAP_INV_G11
XG10092 XI11_3/XI0/XI0_15/d__13_ XI11_3/XI0/XI0_15/d_13_ DECAP_INV_G11
XG10093 XI11_3/XI0/XI0_15/d__12_ XI11_3/XI0/XI0_15/d_12_ DECAP_INV_G11
XG10094 XI11_3/XI0/XI0_15/d__11_ XI11_3/XI0/XI0_15/d_11_ DECAP_INV_G11
XG10095 XI11_3/XI0/XI0_15/d__10_ XI11_3/XI0/XI0_15/d_10_ DECAP_INV_G11
XG10096 XI11_3/XI0/XI0_15/d__9_ XI11_3/XI0/XI0_15/d_9_ DECAP_INV_G11
XG10097 XI11_3/XI0/XI0_15/d__8_ XI11_3/XI0/XI0_15/d_8_ DECAP_INV_G11
XG10098 XI11_3/XI0/XI0_15/d__7_ XI11_3/XI0/XI0_15/d_7_ DECAP_INV_G11
XG10099 XI11_3/XI0/XI0_15/d__6_ XI11_3/XI0/XI0_15/d_6_ DECAP_INV_G11
XG10100 XI11_3/XI0/XI0_15/d__5_ XI11_3/XI0/XI0_15/d_5_ DECAP_INV_G11
XG10101 XI11_3/XI0/XI0_15/d__4_ XI11_3/XI0/XI0_15/d_4_ DECAP_INV_G11
XG10102 XI11_3/XI0/XI0_15/d__3_ XI11_3/XI0/XI0_15/d_3_ DECAP_INV_G11
XG10103 XI11_3/XI0/XI0_15/d__2_ XI11_3/XI0/XI0_15/d_2_ DECAP_INV_G11
XG10104 XI11_3/XI0/XI0_15/d__1_ XI11_3/XI0/XI0_15/d_1_ DECAP_INV_G11
XG10105 XI11_3/XI0/XI0_15/d__0_ XI11_3/XI0/XI0_15/d_0_ DECAP_INV_G11
XG10106 XI11_3/XI0/XI0_15/d_15_ XI11_3/XI0/XI0_15/d__15_ DECAP_INV_G11
XG10107 XI11_3/XI0/XI0_15/d_14_ XI11_3/XI0/XI0_15/d__14_ DECAP_INV_G11
XG10108 XI11_3/XI0/XI0_15/d_13_ XI11_3/XI0/XI0_15/d__13_ DECAP_INV_G11
XG10109 XI11_3/XI0/XI0_15/d_12_ XI11_3/XI0/XI0_15/d__12_ DECAP_INV_G11
XG10110 XI11_3/XI0/XI0_15/d_11_ XI11_3/XI0/XI0_15/d__11_ DECAP_INV_G11
XG10111 XI11_3/XI0/XI0_15/d_10_ XI11_3/XI0/XI0_15/d__10_ DECAP_INV_G11
XG10112 XI11_3/XI0/XI0_15/d_9_ XI11_3/XI0/XI0_15/d__9_ DECAP_INV_G11
XG10113 XI11_3/XI0/XI0_15/d_8_ XI11_3/XI0/XI0_15/d__8_ DECAP_INV_G11
XG10114 XI11_3/XI0/XI0_15/d_7_ XI11_3/XI0/XI0_15/d__7_ DECAP_INV_G11
XG10115 XI11_3/XI0/XI0_15/d_6_ XI11_3/XI0/XI0_15/d__6_ DECAP_INV_G11
XG10116 XI11_3/XI0/XI0_15/d_5_ XI11_3/XI0/XI0_15/d__5_ DECAP_INV_G11
XG10117 XI11_3/XI0/XI0_15/d_4_ XI11_3/XI0/XI0_15/d__4_ DECAP_INV_G11
XG10118 XI11_3/XI0/XI0_15/d_3_ XI11_3/XI0/XI0_15/d__3_ DECAP_INV_G11
XG10119 XI11_3/XI0/XI0_15/d_2_ XI11_3/XI0/XI0_15/d__2_ DECAP_INV_G11
XG10120 XI11_3/XI0/XI0_15/d_1_ XI11_3/XI0/XI0_15/d__1_ DECAP_INV_G11
XG10121 XI11_3/XI0/XI0_15/d_0_ XI11_3/XI0/XI0_15/d__0_ DECAP_INV_G11
XG10122 XI11_3/XI0/XI0_14/d__15_ XI11_3/XI0/XI0_14/d_15_ DECAP_INV_G11
XG10123 XI11_3/XI0/XI0_14/d__14_ XI11_3/XI0/XI0_14/d_14_ DECAP_INV_G11
XG10124 XI11_3/XI0/XI0_14/d__13_ XI11_3/XI0/XI0_14/d_13_ DECAP_INV_G11
XG10125 XI11_3/XI0/XI0_14/d__12_ XI11_3/XI0/XI0_14/d_12_ DECAP_INV_G11
XG10126 XI11_3/XI0/XI0_14/d__11_ XI11_3/XI0/XI0_14/d_11_ DECAP_INV_G11
XG10127 XI11_3/XI0/XI0_14/d__10_ XI11_3/XI0/XI0_14/d_10_ DECAP_INV_G11
XG10128 XI11_3/XI0/XI0_14/d__9_ XI11_3/XI0/XI0_14/d_9_ DECAP_INV_G11
XG10129 XI11_3/XI0/XI0_14/d__8_ XI11_3/XI0/XI0_14/d_8_ DECAP_INV_G11
XG10130 XI11_3/XI0/XI0_14/d__7_ XI11_3/XI0/XI0_14/d_7_ DECAP_INV_G11
XG10131 XI11_3/XI0/XI0_14/d__6_ XI11_3/XI0/XI0_14/d_6_ DECAP_INV_G11
XG10132 XI11_3/XI0/XI0_14/d__5_ XI11_3/XI0/XI0_14/d_5_ DECAP_INV_G11
XG10133 XI11_3/XI0/XI0_14/d__4_ XI11_3/XI0/XI0_14/d_4_ DECAP_INV_G11
XG10134 XI11_3/XI0/XI0_14/d__3_ XI11_3/XI0/XI0_14/d_3_ DECAP_INV_G11
XG10135 XI11_3/XI0/XI0_14/d__2_ XI11_3/XI0/XI0_14/d_2_ DECAP_INV_G11
XG10136 XI11_3/XI0/XI0_14/d__1_ XI11_3/XI0/XI0_14/d_1_ DECAP_INV_G11
XG10137 XI11_3/XI0/XI0_14/d__0_ XI11_3/XI0/XI0_14/d_0_ DECAP_INV_G11
XG10138 XI11_3/XI0/XI0_14/d_15_ XI11_3/XI0/XI0_14/d__15_ DECAP_INV_G11
XG10139 XI11_3/XI0/XI0_14/d_14_ XI11_3/XI0/XI0_14/d__14_ DECAP_INV_G11
XG10140 XI11_3/XI0/XI0_14/d_13_ XI11_3/XI0/XI0_14/d__13_ DECAP_INV_G11
XG10141 XI11_3/XI0/XI0_14/d_12_ XI11_3/XI0/XI0_14/d__12_ DECAP_INV_G11
XG10142 XI11_3/XI0/XI0_14/d_11_ XI11_3/XI0/XI0_14/d__11_ DECAP_INV_G11
XG10143 XI11_3/XI0/XI0_14/d_10_ XI11_3/XI0/XI0_14/d__10_ DECAP_INV_G11
XG10144 XI11_3/XI0/XI0_14/d_9_ XI11_3/XI0/XI0_14/d__9_ DECAP_INV_G11
XG10145 XI11_3/XI0/XI0_14/d_8_ XI11_3/XI0/XI0_14/d__8_ DECAP_INV_G11
XG10146 XI11_3/XI0/XI0_14/d_7_ XI11_3/XI0/XI0_14/d__7_ DECAP_INV_G11
XG10147 XI11_3/XI0/XI0_14/d_6_ XI11_3/XI0/XI0_14/d__6_ DECAP_INV_G11
XG10148 XI11_3/XI0/XI0_14/d_5_ XI11_3/XI0/XI0_14/d__5_ DECAP_INV_G11
XG10149 XI11_3/XI0/XI0_14/d_4_ XI11_3/XI0/XI0_14/d__4_ DECAP_INV_G11
XG10150 XI11_3/XI0/XI0_14/d_3_ XI11_3/XI0/XI0_14/d__3_ DECAP_INV_G11
XG10151 XI11_3/XI0/XI0_14/d_2_ XI11_3/XI0/XI0_14/d__2_ DECAP_INV_G11
XG10152 XI11_3/XI0/XI0_14/d_1_ XI11_3/XI0/XI0_14/d__1_ DECAP_INV_G11
XG10153 XI11_3/XI0/XI0_14/d_0_ XI11_3/XI0/XI0_14/d__0_ DECAP_INV_G11
XG10154 XI11_3/XI0/XI0_13/d__15_ XI11_3/XI0/XI0_13/d_15_ DECAP_INV_G11
XG10155 XI11_3/XI0/XI0_13/d__14_ XI11_3/XI0/XI0_13/d_14_ DECAP_INV_G11
XG10156 XI11_3/XI0/XI0_13/d__13_ XI11_3/XI0/XI0_13/d_13_ DECAP_INV_G11
XG10157 XI11_3/XI0/XI0_13/d__12_ XI11_3/XI0/XI0_13/d_12_ DECAP_INV_G11
XG10158 XI11_3/XI0/XI0_13/d__11_ XI11_3/XI0/XI0_13/d_11_ DECAP_INV_G11
XG10159 XI11_3/XI0/XI0_13/d__10_ XI11_3/XI0/XI0_13/d_10_ DECAP_INV_G11
XG10160 XI11_3/XI0/XI0_13/d__9_ XI11_3/XI0/XI0_13/d_9_ DECAP_INV_G11
XG10161 XI11_3/XI0/XI0_13/d__8_ XI11_3/XI0/XI0_13/d_8_ DECAP_INV_G11
XG10162 XI11_3/XI0/XI0_13/d__7_ XI11_3/XI0/XI0_13/d_7_ DECAP_INV_G11
XG10163 XI11_3/XI0/XI0_13/d__6_ XI11_3/XI0/XI0_13/d_6_ DECAP_INV_G11
XG10164 XI11_3/XI0/XI0_13/d__5_ XI11_3/XI0/XI0_13/d_5_ DECAP_INV_G11
XG10165 XI11_3/XI0/XI0_13/d__4_ XI11_3/XI0/XI0_13/d_4_ DECAP_INV_G11
XG10166 XI11_3/XI0/XI0_13/d__3_ XI11_3/XI0/XI0_13/d_3_ DECAP_INV_G11
XG10167 XI11_3/XI0/XI0_13/d__2_ XI11_3/XI0/XI0_13/d_2_ DECAP_INV_G11
XG10168 XI11_3/XI0/XI0_13/d__1_ XI11_3/XI0/XI0_13/d_1_ DECAP_INV_G11
XG10169 XI11_3/XI0/XI0_13/d__0_ XI11_3/XI0/XI0_13/d_0_ DECAP_INV_G11
XG10170 XI11_3/XI0/XI0_13/d_15_ XI11_3/XI0/XI0_13/d__15_ DECAP_INV_G11
XG10171 XI11_3/XI0/XI0_13/d_14_ XI11_3/XI0/XI0_13/d__14_ DECAP_INV_G11
XG10172 XI11_3/XI0/XI0_13/d_13_ XI11_3/XI0/XI0_13/d__13_ DECAP_INV_G11
XG10173 XI11_3/XI0/XI0_13/d_12_ XI11_3/XI0/XI0_13/d__12_ DECAP_INV_G11
XG10174 XI11_3/XI0/XI0_13/d_11_ XI11_3/XI0/XI0_13/d__11_ DECAP_INV_G11
XG10175 XI11_3/XI0/XI0_13/d_10_ XI11_3/XI0/XI0_13/d__10_ DECAP_INV_G11
XG10176 XI11_3/XI0/XI0_13/d_9_ XI11_3/XI0/XI0_13/d__9_ DECAP_INV_G11
XG10177 XI11_3/XI0/XI0_13/d_8_ XI11_3/XI0/XI0_13/d__8_ DECAP_INV_G11
XG10178 XI11_3/XI0/XI0_13/d_7_ XI11_3/XI0/XI0_13/d__7_ DECAP_INV_G11
XG10179 XI11_3/XI0/XI0_13/d_6_ XI11_3/XI0/XI0_13/d__6_ DECAP_INV_G11
XG10180 XI11_3/XI0/XI0_13/d_5_ XI11_3/XI0/XI0_13/d__5_ DECAP_INV_G11
XG10181 XI11_3/XI0/XI0_13/d_4_ XI11_3/XI0/XI0_13/d__4_ DECAP_INV_G11
XG10182 XI11_3/XI0/XI0_13/d_3_ XI11_3/XI0/XI0_13/d__3_ DECAP_INV_G11
XG10183 XI11_3/XI0/XI0_13/d_2_ XI11_3/XI0/XI0_13/d__2_ DECAP_INV_G11
XG10184 XI11_3/XI0/XI0_13/d_1_ XI11_3/XI0/XI0_13/d__1_ DECAP_INV_G11
XG10185 XI11_3/XI0/XI0_13/d_0_ XI11_3/XI0/XI0_13/d__0_ DECAP_INV_G11
XG10186 XI11_3/XI0/XI0_12/d__15_ XI11_3/XI0/XI0_12/d_15_ DECAP_INV_G11
XG10187 XI11_3/XI0/XI0_12/d__14_ XI11_3/XI0/XI0_12/d_14_ DECAP_INV_G11
XG10188 XI11_3/XI0/XI0_12/d__13_ XI11_3/XI0/XI0_12/d_13_ DECAP_INV_G11
XG10189 XI11_3/XI0/XI0_12/d__12_ XI11_3/XI0/XI0_12/d_12_ DECAP_INV_G11
XG10190 XI11_3/XI0/XI0_12/d__11_ XI11_3/XI0/XI0_12/d_11_ DECAP_INV_G11
XG10191 XI11_3/XI0/XI0_12/d__10_ XI11_3/XI0/XI0_12/d_10_ DECAP_INV_G11
XG10192 XI11_3/XI0/XI0_12/d__9_ XI11_3/XI0/XI0_12/d_9_ DECAP_INV_G11
XG10193 XI11_3/XI0/XI0_12/d__8_ XI11_3/XI0/XI0_12/d_8_ DECAP_INV_G11
XG10194 XI11_3/XI0/XI0_12/d__7_ XI11_3/XI0/XI0_12/d_7_ DECAP_INV_G11
XG10195 XI11_3/XI0/XI0_12/d__6_ XI11_3/XI0/XI0_12/d_6_ DECAP_INV_G11
XG10196 XI11_3/XI0/XI0_12/d__5_ XI11_3/XI0/XI0_12/d_5_ DECAP_INV_G11
XG10197 XI11_3/XI0/XI0_12/d__4_ XI11_3/XI0/XI0_12/d_4_ DECAP_INV_G11
XG10198 XI11_3/XI0/XI0_12/d__3_ XI11_3/XI0/XI0_12/d_3_ DECAP_INV_G11
XG10199 XI11_3/XI0/XI0_12/d__2_ XI11_3/XI0/XI0_12/d_2_ DECAP_INV_G11
XG10200 XI11_3/XI0/XI0_12/d__1_ XI11_3/XI0/XI0_12/d_1_ DECAP_INV_G11
XG10201 XI11_3/XI0/XI0_12/d__0_ XI11_3/XI0/XI0_12/d_0_ DECAP_INV_G11
XG10202 XI11_3/XI0/XI0_12/d_15_ XI11_3/XI0/XI0_12/d__15_ DECAP_INV_G11
XG10203 XI11_3/XI0/XI0_12/d_14_ XI11_3/XI0/XI0_12/d__14_ DECAP_INV_G11
XG10204 XI11_3/XI0/XI0_12/d_13_ XI11_3/XI0/XI0_12/d__13_ DECAP_INV_G11
XG10205 XI11_3/XI0/XI0_12/d_12_ XI11_3/XI0/XI0_12/d__12_ DECAP_INV_G11
XG10206 XI11_3/XI0/XI0_12/d_11_ XI11_3/XI0/XI0_12/d__11_ DECAP_INV_G11
XG10207 XI11_3/XI0/XI0_12/d_10_ XI11_3/XI0/XI0_12/d__10_ DECAP_INV_G11
XG10208 XI11_3/XI0/XI0_12/d_9_ XI11_3/XI0/XI0_12/d__9_ DECAP_INV_G11
XG10209 XI11_3/XI0/XI0_12/d_8_ XI11_3/XI0/XI0_12/d__8_ DECAP_INV_G11
XG10210 XI11_3/XI0/XI0_12/d_7_ XI11_3/XI0/XI0_12/d__7_ DECAP_INV_G11
XG10211 XI11_3/XI0/XI0_12/d_6_ XI11_3/XI0/XI0_12/d__6_ DECAP_INV_G11
XG10212 XI11_3/XI0/XI0_12/d_5_ XI11_3/XI0/XI0_12/d__5_ DECAP_INV_G11
XG10213 XI11_3/XI0/XI0_12/d_4_ XI11_3/XI0/XI0_12/d__4_ DECAP_INV_G11
XG10214 XI11_3/XI0/XI0_12/d_3_ XI11_3/XI0/XI0_12/d__3_ DECAP_INV_G11
XG10215 XI11_3/XI0/XI0_12/d_2_ XI11_3/XI0/XI0_12/d__2_ DECAP_INV_G11
XG10216 XI11_3/XI0/XI0_12/d_1_ XI11_3/XI0/XI0_12/d__1_ DECAP_INV_G11
XG10217 XI11_3/XI0/XI0_12/d_0_ XI11_3/XI0/XI0_12/d__0_ DECAP_INV_G11
XG10218 XI11_3/XI0/XI0_11/d__15_ XI11_3/XI0/XI0_11/d_15_ DECAP_INV_G11
XG10219 XI11_3/XI0/XI0_11/d__14_ XI11_3/XI0/XI0_11/d_14_ DECAP_INV_G11
XG10220 XI11_3/XI0/XI0_11/d__13_ XI11_3/XI0/XI0_11/d_13_ DECAP_INV_G11
XG10221 XI11_3/XI0/XI0_11/d__12_ XI11_3/XI0/XI0_11/d_12_ DECAP_INV_G11
XG10222 XI11_3/XI0/XI0_11/d__11_ XI11_3/XI0/XI0_11/d_11_ DECAP_INV_G11
XG10223 XI11_3/XI0/XI0_11/d__10_ XI11_3/XI0/XI0_11/d_10_ DECAP_INV_G11
XG10224 XI11_3/XI0/XI0_11/d__9_ XI11_3/XI0/XI0_11/d_9_ DECAP_INV_G11
XG10225 XI11_3/XI0/XI0_11/d__8_ XI11_3/XI0/XI0_11/d_8_ DECAP_INV_G11
XG10226 XI11_3/XI0/XI0_11/d__7_ XI11_3/XI0/XI0_11/d_7_ DECAP_INV_G11
XG10227 XI11_3/XI0/XI0_11/d__6_ XI11_3/XI0/XI0_11/d_6_ DECAP_INV_G11
XG10228 XI11_3/XI0/XI0_11/d__5_ XI11_3/XI0/XI0_11/d_5_ DECAP_INV_G11
XG10229 XI11_3/XI0/XI0_11/d__4_ XI11_3/XI0/XI0_11/d_4_ DECAP_INV_G11
XG10230 XI11_3/XI0/XI0_11/d__3_ XI11_3/XI0/XI0_11/d_3_ DECAP_INV_G11
XG10231 XI11_3/XI0/XI0_11/d__2_ XI11_3/XI0/XI0_11/d_2_ DECAP_INV_G11
XG10232 XI11_3/XI0/XI0_11/d__1_ XI11_3/XI0/XI0_11/d_1_ DECAP_INV_G11
XG10233 XI11_3/XI0/XI0_11/d__0_ XI11_3/XI0/XI0_11/d_0_ DECAP_INV_G11
XG10234 XI11_3/XI0/XI0_11/d_15_ XI11_3/XI0/XI0_11/d__15_ DECAP_INV_G11
XG10235 XI11_3/XI0/XI0_11/d_14_ XI11_3/XI0/XI0_11/d__14_ DECAP_INV_G11
XG10236 XI11_3/XI0/XI0_11/d_13_ XI11_3/XI0/XI0_11/d__13_ DECAP_INV_G11
XG10237 XI11_3/XI0/XI0_11/d_12_ XI11_3/XI0/XI0_11/d__12_ DECAP_INV_G11
XG10238 XI11_3/XI0/XI0_11/d_11_ XI11_3/XI0/XI0_11/d__11_ DECAP_INV_G11
XG10239 XI11_3/XI0/XI0_11/d_10_ XI11_3/XI0/XI0_11/d__10_ DECAP_INV_G11
XG10240 XI11_3/XI0/XI0_11/d_9_ XI11_3/XI0/XI0_11/d__9_ DECAP_INV_G11
XG10241 XI11_3/XI0/XI0_11/d_8_ XI11_3/XI0/XI0_11/d__8_ DECAP_INV_G11
XG10242 XI11_3/XI0/XI0_11/d_7_ XI11_3/XI0/XI0_11/d__7_ DECAP_INV_G11
XG10243 XI11_3/XI0/XI0_11/d_6_ XI11_3/XI0/XI0_11/d__6_ DECAP_INV_G11
XG10244 XI11_3/XI0/XI0_11/d_5_ XI11_3/XI0/XI0_11/d__5_ DECAP_INV_G11
XG10245 XI11_3/XI0/XI0_11/d_4_ XI11_3/XI0/XI0_11/d__4_ DECAP_INV_G11
XG10246 XI11_3/XI0/XI0_11/d_3_ XI11_3/XI0/XI0_11/d__3_ DECAP_INV_G11
XG10247 XI11_3/XI0/XI0_11/d_2_ XI11_3/XI0/XI0_11/d__2_ DECAP_INV_G11
XG10248 XI11_3/XI0/XI0_11/d_1_ XI11_3/XI0/XI0_11/d__1_ DECAP_INV_G11
XG10249 XI11_3/XI0/XI0_11/d_0_ XI11_3/XI0/XI0_11/d__0_ DECAP_INV_G11
XG10250 XI11_3/XI0/XI0_10/d__15_ XI11_3/XI0/XI0_10/d_15_ DECAP_INV_G11
XG10251 XI11_3/XI0/XI0_10/d__14_ XI11_3/XI0/XI0_10/d_14_ DECAP_INV_G11
XG10252 XI11_3/XI0/XI0_10/d__13_ XI11_3/XI0/XI0_10/d_13_ DECAP_INV_G11
XG10253 XI11_3/XI0/XI0_10/d__12_ XI11_3/XI0/XI0_10/d_12_ DECAP_INV_G11
XG10254 XI11_3/XI0/XI0_10/d__11_ XI11_3/XI0/XI0_10/d_11_ DECAP_INV_G11
XG10255 XI11_3/XI0/XI0_10/d__10_ XI11_3/XI0/XI0_10/d_10_ DECAP_INV_G11
XG10256 XI11_3/XI0/XI0_10/d__9_ XI11_3/XI0/XI0_10/d_9_ DECAP_INV_G11
XG10257 XI11_3/XI0/XI0_10/d__8_ XI11_3/XI0/XI0_10/d_8_ DECAP_INV_G11
XG10258 XI11_3/XI0/XI0_10/d__7_ XI11_3/XI0/XI0_10/d_7_ DECAP_INV_G11
XG10259 XI11_3/XI0/XI0_10/d__6_ XI11_3/XI0/XI0_10/d_6_ DECAP_INV_G11
XG10260 XI11_3/XI0/XI0_10/d__5_ XI11_3/XI0/XI0_10/d_5_ DECAP_INV_G11
XG10261 XI11_3/XI0/XI0_10/d__4_ XI11_3/XI0/XI0_10/d_4_ DECAP_INV_G11
XG10262 XI11_3/XI0/XI0_10/d__3_ XI11_3/XI0/XI0_10/d_3_ DECAP_INV_G11
XG10263 XI11_3/XI0/XI0_10/d__2_ XI11_3/XI0/XI0_10/d_2_ DECAP_INV_G11
XG10264 XI11_3/XI0/XI0_10/d__1_ XI11_3/XI0/XI0_10/d_1_ DECAP_INV_G11
XG10265 XI11_3/XI0/XI0_10/d__0_ XI11_3/XI0/XI0_10/d_0_ DECAP_INV_G11
XG10266 XI11_3/XI0/XI0_10/d_15_ XI11_3/XI0/XI0_10/d__15_ DECAP_INV_G11
XG10267 XI11_3/XI0/XI0_10/d_14_ XI11_3/XI0/XI0_10/d__14_ DECAP_INV_G11
XG10268 XI11_3/XI0/XI0_10/d_13_ XI11_3/XI0/XI0_10/d__13_ DECAP_INV_G11
XG10269 XI11_3/XI0/XI0_10/d_12_ XI11_3/XI0/XI0_10/d__12_ DECAP_INV_G11
XG10270 XI11_3/XI0/XI0_10/d_11_ XI11_3/XI0/XI0_10/d__11_ DECAP_INV_G11
XG10271 XI11_3/XI0/XI0_10/d_10_ XI11_3/XI0/XI0_10/d__10_ DECAP_INV_G11
XG10272 XI11_3/XI0/XI0_10/d_9_ XI11_3/XI0/XI0_10/d__9_ DECAP_INV_G11
XG10273 XI11_3/XI0/XI0_10/d_8_ XI11_3/XI0/XI0_10/d__8_ DECAP_INV_G11
XG10274 XI11_3/XI0/XI0_10/d_7_ XI11_3/XI0/XI0_10/d__7_ DECAP_INV_G11
XG10275 XI11_3/XI0/XI0_10/d_6_ XI11_3/XI0/XI0_10/d__6_ DECAP_INV_G11
XG10276 XI11_3/XI0/XI0_10/d_5_ XI11_3/XI0/XI0_10/d__5_ DECAP_INV_G11
XG10277 XI11_3/XI0/XI0_10/d_4_ XI11_3/XI0/XI0_10/d__4_ DECAP_INV_G11
XG10278 XI11_3/XI0/XI0_10/d_3_ XI11_3/XI0/XI0_10/d__3_ DECAP_INV_G11
XG10279 XI11_3/XI0/XI0_10/d_2_ XI11_3/XI0/XI0_10/d__2_ DECAP_INV_G11
XG10280 XI11_3/XI0/XI0_10/d_1_ XI11_3/XI0/XI0_10/d__1_ DECAP_INV_G11
XG10281 XI11_3/XI0/XI0_10/d_0_ XI11_3/XI0/XI0_10/d__0_ DECAP_INV_G11
XG10282 XI11_3/XI0/XI0_9/d__15_ XI11_3/XI0/XI0_9/d_15_ DECAP_INV_G11
XG10283 XI11_3/XI0/XI0_9/d__14_ XI11_3/XI0/XI0_9/d_14_ DECAP_INV_G11
XG10284 XI11_3/XI0/XI0_9/d__13_ XI11_3/XI0/XI0_9/d_13_ DECAP_INV_G11
XG10285 XI11_3/XI0/XI0_9/d__12_ XI11_3/XI0/XI0_9/d_12_ DECAP_INV_G11
XG10286 XI11_3/XI0/XI0_9/d__11_ XI11_3/XI0/XI0_9/d_11_ DECAP_INV_G11
XG10287 XI11_3/XI0/XI0_9/d__10_ XI11_3/XI0/XI0_9/d_10_ DECAP_INV_G11
XG10288 XI11_3/XI0/XI0_9/d__9_ XI11_3/XI0/XI0_9/d_9_ DECAP_INV_G11
XG10289 XI11_3/XI0/XI0_9/d__8_ XI11_3/XI0/XI0_9/d_8_ DECAP_INV_G11
XG10290 XI11_3/XI0/XI0_9/d__7_ XI11_3/XI0/XI0_9/d_7_ DECAP_INV_G11
XG10291 XI11_3/XI0/XI0_9/d__6_ XI11_3/XI0/XI0_9/d_6_ DECAP_INV_G11
XG10292 XI11_3/XI0/XI0_9/d__5_ XI11_3/XI0/XI0_9/d_5_ DECAP_INV_G11
XG10293 XI11_3/XI0/XI0_9/d__4_ XI11_3/XI0/XI0_9/d_4_ DECAP_INV_G11
XG10294 XI11_3/XI0/XI0_9/d__3_ XI11_3/XI0/XI0_9/d_3_ DECAP_INV_G11
XG10295 XI11_3/XI0/XI0_9/d__2_ XI11_3/XI0/XI0_9/d_2_ DECAP_INV_G11
XG10296 XI11_3/XI0/XI0_9/d__1_ XI11_3/XI0/XI0_9/d_1_ DECAP_INV_G11
XG10297 XI11_3/XI0/XI0_9/d__0_ XI11_3/XI0/XI0_9/d_0_ DECAP_INV_G11
XG10298 XI11_3/XI0/XI0_9/d_15_ XI11_3/XI0/XI0_9/d__15_ DECAP_INV_G11
XG10299 XI11_3/XI0/XI0_9/d_14_ XI11_3/XI0/XI0_9/d__14_ DECAP_INV_G11
XG10300 XI11_3/XI0/XI0_9/d_13_ XI11_3/XI0/XI0_9/d__13_ DECAP_INV_G11
XG10301 XI11_3/XI0/XI0_9/d_12_ XI11_3/XI0/XI0_9/d__12_ DECAP_INV_G11
XG10302 XI11_3/XI0/XI0_9/d_11_ XI11_3/XI0/XI0_9/d__11_ DECAP_INV_G11
XG10303 XI11_3/XI0/XI0_9/d_10_ XI11_3/XI0/XI0_9/d__10_ DECAP_INV_G11
XG10304 XI11_3/XI0/XI0_9/d_9_ XI11_3/XI0/XI0_9/d__9_ DECAP_INV_G11
XG10305 XI11_3/XI0/XI0_9/d_8_ XI11_3/XI0/XI0_9/d__8_ DECAP_INV_G11
XG10306 XI11_3/XI0/XI0_9/d_7_ XI11_3/XI0/XI0_9/d__7_ DECAP_INV_G11
XG10307 XI11_3/XI0/XI0_9/d_6_ XI11_3/XI0/XI0_9/d__6_ DECAP_INV_G11
XG10308 XI11_3/XI0/XI0_9/d_5_ XI11_3/XI0/XI0_9/d__5_ DECAP_INV_G11
XG10309 XI11_3/XI0/XI0_9/d_4_ XI11_3/XI0/XI0_9/d__4_ DECAP_INV_G11
XG10310 XI11_3/XI0/XI0_9/d_3_ XI11_3/XI0/XI0_9/d__3_ DECAP_INV_G11
XG10311 XI11_3/XI0/XI0_9/d_2_ XI11_3/XI0/XI0_9/d__2_ DECAP_INV_G11
XG10312 XI11_3/XI0/XI0_9/d_1_ XI11_3/XI0/XI0_9/d__1_ DECAP_INV_G11
XG10313 XI11_3/XI0/XI0_9/d_0_ XI11_3/XI0/XI0_9/d__0_ DECAP_INV_G11
XG10314 XI11_3/XI0/XI0_8/d__15_ XI11_3/XI0/XI0_8/d_15_ DECAP_INV_G11
XG10315 XI11_3/XI0/XI0_8/d__14_ XI11_3/XI0/XI0_8/d_14_ DECAP_INV_G11
XG10316 XI11_3/XI0/XI0_8/d__13_ XI11_3/XI0/XI0_8/d_13_ DECAP_INV_G11
XG10317 XI11_3/XI0/XI0_8/d__12_ XI11_3/XI0/XI0_8/d_12_ DECAP_INV_G11
XG10318 XI11_3/XI0/XI0_8/d__11_ XI11_3/XI0/XI0_8/d_11_ DECAP_INV_G11
XG10319 XI11_3/XI0/XI0_8/d__10_ XI11_3/XI0/XI0_8/d_10_ DECAP_INV_G11
XG10320 XI11_3/XI0/XI0_8/d__9_ XI11_3/XI0/XI0_8/d_9_ DECAP_INV_G11
XG10321 XI11_3/XI0/XI0_8/d__8_ XI11_3/XI0/XI0_8/d_8_ DECAP_INV_G11
XG10322 XI11_3/XI0/XI0_8/d__7_ XI11_3/XI0/XI0_8/d_7_ DECAP_INV_G11
XG10323 XI11_3/XI0/XI0_8/d__6_ XI11_3/XI0/XI0_8/d_6_ DECAP_INV_G11
XG10324 XI11_3/XI0/XI0_8/d__5_ XI11_3/XI0/XI0_8/d_5_ DECAP_INV_G11
XG10325 XI11_3/XI0/XI0_8/d__4_ XI11_3/XI0/XI0_8/d_4_ DECAP_INV_G11
XG10326 XI11_3/XI0/XI0_8/d__3_ XI11_3/XI0/XI0_8/d_3_ DECAP_INV_G11
XG10327 XI11_3/XI0/XI0_8/d__2_ XI11_3/XI0/XI0_8/d_2_ DECAP_INV_G11
XG10328 XI11_3/XI0/XI0_8/d__1_ XI11_3/XI0/XI0_8/d_1_ DECAP_INV_G11
XG10329 XI11_3/XI0/XI0_8/d__0_ XI11_3/XI0/XI0_8/d_0_ DECAP_INV_G11
XG10330 XI11_3/XI0/XI0_8/d_15_ XI11_3/XI0/XI0_8/d__15_ DECAP_INV_G11
XG10331 XI11_3/XI0/XI0_8/d_14_ XI11_3/XI0/XI0_8/d__14_ DECAP_INV_G11
XG10332 XI11_3/XI0/XI0_8/d_13_ XI11_3/XI0/XI0_8/d__13_ DECAP_INV_G11
XG10333 XI11_3/XI0/XI0_8/d_12_ XI11_3/XI0/XI0_8/d__12_ DECAP_INV_G11
XG10334 XI11_3/XI0/XI0_8/d_11_ XI11_3/XI0/XI0_8/d__11_ DECAP_INV_G11
XG10335 XI11_3/XI0/XI0_8/d_10_ XI11_3/XI0/XI0_8/d__10_ DECAP_INV_G11
XG10336 XI11_3/XI0/XI0_8/d_9_ XI11_3/XI0/XI0_8/d__9_ DECAP_INV_G11
XG10337 XI11_3/XI0/XI0_8/d_8_ XI11_3/XI0/XI0_8/d__8_ DECAP_INV_G11
XG10338 XI11_3/XI0/XI0_8/d_7_ XI11_3/XI0/XI0_8/d__7_ DECAP_INV_G11
XG10339 XI11_3/XI0/XI0_8/d_6_ XI11_3/XI0/XI0_8/d__6_ DECAP_INV_G11
XG10340 XI11_3/XI0/XI0_8/d_5_ XI11_3/XI0/XI0_8/d__5_ DECAP_INV_G11
XG10341 XI11_3/XI0/XI0_8/d_4_ XI11_3/XI0/XI0_8/d__4_ DECAP_INV_G11
XG10342 XI11_3/XI0/XI0_8/d_3_ XI11_3/XI0/XI0_8/d__3_ DECAP_INV_G11
XG10343 XI11_3/XI0/XI0_8/d_2_ XI11_3/XI0/XI0_8/d__2_ DECAP_INV_G11
XG10344 XI11_3/XI0/XI0_8/d_1_ XI11_3/XI0/XI0_8/d__1_ DECAP_INV_G11
XG10345 XI11_3/XI0/XI0_8/d_0_ XI11_3/XI0/XI0_8/d__0_ DECAP_INV_G11
XG10346 XI11_3/XI0/XI0_7/d__15_ XI11_3/XI0/XI0_7/d_15_ DECAP_INV_G11
XG10347 XI11_3/XI0/XI0_7/d__14_ XI11_3/XI0/XI0_7/d_14_ DECAP_INV_G11
XG10348 XI11_3/XI0/XI0_7/d__13_ XI11_3/XI0/XI0_7/d_13_ DECAP_INV_G11
XG10349 XI11_3/XI0/XI0_7/d__12_ XI11_3/XI0/XI0_7/d_12_ DECAP_INV_G11
XG10350 XI11_3/XI0/XI0_7/d__11_ XI11_3/XI0/XI0_7/d_11_ DECAP_INV_G11
XG10351 XI11_3/XI0/XI0_7/d__10_ XI11_3/XI0/XI0_7/d_10_ DECAP_INV_G11
XG10352 XI11_3/XI0/XI0_7/d__9_ XI11_3/XI0/XI0_7/d_9_ DECAP_INV_G11
XG10353 XI11_3/XI0/XI0_7/d__8_ XI11_3/XI0/XI0_7/d_8_ DECAP_INV_G11
XG10354 XI11_3/XI0/XI0_7/d__7_ XI11_3/XI0/XI0_7/d_7_ DECAP_INV_G11
XG10355 XI11_3/XI0/XI0_7/d__6_ XI11_3/XI0/XI0_7/d_6_ DECAP_INV_G11
XG10356 XI11_3/XI0/XI0_7/d__5_ XI11_3/XI0/XI0_7/d_5_ DECAP_INV_G11
XG10357 XI11_3/XI0/XI0_7/d__4_ XI11_3/XI0/XI0_7/d_4_ DECAP_INV_G11
XG10358 XI11_3/XI0/XI0_7/d__3_ XI11_3/XI0/XI0_7/d_3_ DECAP_INV_G11
XG10359 XI11_3/XI0/XI0_7/d__2_ XI11_3/XI0/XI0_7/d_2_ DECAP_INV_G11
XG10360 XI11_3/XI0/XI0_7/d__1_ XI11_3/XI0/XI0_7/d_1_ DECAP_INV_G11
XG10361 XI11_3/XI0/XI0_7/d__0_ XI11_3/XI0/XI0_7/d_0_ DECAP_INV_G11
XG10362 XI11_3/XI0/XI0_7/d_15_ XI11_3/XI0/XI0_7/d__15_ DECAP_INV_G11
XG10363 XI11_3/XI0/XI0_7/d_14_ XI11_3/XI0/XI0_7/d__14_ DECAP_INV_G11
XG10364 XI11_3/XI0/XI0_7/d_13_ XI11_3/XI0/XI0_7/d__13_ DECAP_INV_G11
XG10365 XI11_3/XI0/XI0_7/d_12_ XI11_3/XI0/XI0_7/d__12_ DECAP_INV_G11
XG10366 XI11_3/XI0/XI0_7/d_11_ XI11_3/XI0/XI0_7/d__11_ DECAP_INV_G11
XG10367 XI11_3/XI0/XI0_7/d_10_ XI11_3/XI0/XI0_7/d__10_ DECAP_INV_G11
XG10368 XI11_3/XI0/XI0_7/d_9_ XI11_3/XI0/XI0_7/d__9_ DECAP_INV_G11
XG10369 XI11_3/XI0/XI0_7/d_8_ XI11_3/XI0/XI0_7/d__8_ DECAP_INV_G11
XG10370 XI11_3/XI0/XI0_7/d_7_ XI11_3/XI0/XI0_7/d__7_ DECAP_INV_G11
XG10371 XI11_3/XI0/XI0_7/d_6_ XI11_3/XI0/XI0_7/d__6_ DECAP_INV_G11
XG10372 XI11_3/XI0/XI0_7/d_5_ XI11_3/XI0/XI0_7/d__5_ DECAP_INV_G11
XG10373 XI11_3/XI0/XI0_7/d_4_ XI11_3/XI0/XI0_7/d__4_ DECAP_INV_G11
XG10374 XI11_3/XI0/XI0_7/d_3_ XI11_3/XI0/XI0_7/d__3_ DECAP_INV_G11
XG10375 XI11_3/XI0/XI0_7/d_2_ XI11_3/XI0/XI0_7/d__2_ DECAP_INV_G11
XG10376 XI11_3/XI0/XI0_7/d_1_ XI11_3/XI0/XI0_7/d__1_ DECAP_INV_G11
XG10377 XI11_3/XI0/XI0_7/d_0_ XI11_3/XI0/XI0_7/d__0_ DECAP_INV_G11
XG10378 XI11_3/XI0/XI0_6/d__15_ XI11_3/XI0/XI0_6/d_15_ DECAP_INV_G11
XG10379 XI11_3/XI0/XI0_6/d__14_ XI11_3/XI0/XI0_6/d_14_ DECAP_INV_G11
XG10380 XI11_3/XI0/XI0_6/d__13_ XI11_3/XI0/XI0_6/d_13_ DECAP_INV_G11
XG10381 XI11_3/XI0/XI0_6/d__12_ XI11_3/XI0/XI0_6/d_12_ DECAP_INV_G11
XG10382 XI11_3/XI0/XI0_6/d__11_ XI11_3/XI0/XI0_6/d_11_ DECAP_INV_G11
XG10383 XI11_3/XI0/XI0_6/d__10_ XI11_3/XI0/XI0_6/d_10_ DECAP_INV_G11
XG10384 XI11_3/XI0/XI0_6/d__9_ XI11_3/XI0/XI0_6/d_9_ DECAP_INV_G11
XG10385 XI11_3/XI0/XI0_6/d__8_ XI11_3/XI0/XI0_6/d_8_ DECAP_INV_G11
XG10386 XI11_3/XI0/XI0_6/d__7_ XI11_3/XI0/XI0_6/d_7_ DECAP_INV_G11
XG10387 XI11_3/XI0/XI0_6/d__6_ XI11_3/XI0/XI0_6/d_6_ DECAP_INV_G11
XG10388 XI11_3/XI0/XI0_6/d__5_ XI11_3/XI0/XI0_6/d_5_ DECAP_INV_G11
XG10389 XI11_3/XI0/XI0_6/d__4_ XI11_3/XI0/XI0_6/d_4_ DECAP_INV_G11
XG10390 XI11_3/XI0/XI0_6/d__3_ XI11_3/XI0/XI0_6/d_3_ DECAP_INV_G11
XG10391 XI11_3/XI0/XI0_6/d__2_ XI11_3/XI0/XI0_6/d_2_ DECAP_INV_G11
XG10392 XI11_3/XI0/XI0_6/d__1_ XI11_3/XI0/XI0_6/d_1_ DECAP_INV_G11
XG10393 XI11_3/XI0/XI0_6/d__0_ XI11_3/XI0/XI0_6/d_0_ DECAP_INV_G11
XG10394 XI11_3/XI0/XI0_6/d_15_ XI11_3/XI0/XI0_6/d__15_ DECAP_INV_G11
XG10395 XI11_3/XI0/XI0_6/d_14_ XI11_3/XI0/XI0_6/d__14_ DECAP_INV_G11
XG10396 XI11_3/XI0/XI0_6/d_13_ XI11_3/XI0/XI0_6/d__13_ DECAP_INV_G11
XG10397 XI11_3/XI0/XI0_6/d_12_ XI11_3/XI0/XI0_6/d__12_ DECAP_INV_G11
XG10398 XI11_3/XI0/XI0_6/d_11_ XI11_3/XI0/XI0_6/d__11_ DECAP_INV_G11
XG10399 XI11_3/XI0/XI0_6/d_10_ XI11_3/XI0/XI0_6/d__10_ DECAP_INV_G11
XG10400 XI11_3/XI0/XI0_6/d_9_ XI11_3/XI0/XI0_6/d__9_ DECAP_INV_G11
XG10401 XI11_3/XI0/XI0_6/d_8_ XI11_3/XI0/XI0_6/d__8_ DECAP_INV_G11
XG10402 XI11_3/XI0/XI0_6/d_7_ XI11_3/XI0/XI0_6/d__7_ DECAP_INV_G11
XG10403 XI11_3/XI0/XI0_6/d_6_ XI11_3/XI0/XI0_6/d__6_ DECAP_INV_G11
XG10404 XI11_3/XI0/XI0_6/d_5_ XI11_3/XI0/XI0_6/d__5_ DECAP_INV_G11
XG10405 XI11_3/XI0/XI0_6/d_4_ XI11_3/XI0/XI0_6/d__4_ DECAP_INV_G11
XG10406 XI11_3/XI0/XI0_6/d_3_ XI11_3/XI0/XI0_6/d__3_ DECAP_INV_G11
XG10407 XI11_3/XI0/XI0_6/d_2_ XI11_3/XI0/XI0_6/d__2_ DECAP_INV_G11
XG10408 XI11_3/XI0/XI0_6/d_1_ XI11_3/XI0/XI0_6/d__1_ DECAP_INV_G11
XG10409 XI11_3/XI0/XI0_6/d_0_ XI11_3/XI0/XI0_6/d__0_ DECAP_INV_G11
XG10410 XI11_3/XI0/XI0_5/d__15_ XI11_3/XI0/XI0_5/d_15_ DECAP_INV_G11
XG10411 XI11_3/XI0/XI0_5/d__14_ XI11_3/XI0/XI0_5/d_14_ DECAP_INV_G11
XG10412 XI11_3/XI0/XI0_5/d__13_ XI11_3/XI0/XI0_5/d_13_ DECAP_INV_G11
XG10413 XI11_3/XI0/XI0_5/d__12_ XI11_3/XI0/XI0_5/d_12_ DECAP_INV_G11
XG10414 XI11_3/XI0/XI0_5/d__11_ XI11_3/XI0/XI0_5/d_11_ DECAP_INV_G11
XG10415 XI11_3/XI0/XI0_5/d__10_ XI11_3/XI0/XI0_5/d_10_ DECAP_INV_G11
XG10416 XI11_3/XI0/XI0_5/d__9_ XI11_3/XI0/XI0_5/d_9_ DECAP_INV_G11
XG10417 XI11_3/XI0/XI0_5/d__8_ XI11_3/XI0/XI0_5/d_8_ DECAP_INV_G11
XG10418 XI11_3/XI0/XI0_5/d__7_ XI11_3/XI0/XI0_5/d_7_ DECAP_INV_G11
XG10419 XI11_3/XI0/XI0_5/d__6_ XI11_3/XI0/XI0_5/d_6_ DECAP_INV_G11
XG10420 XI11_3/XI0/XI0_5/d__5_ XI11_3/XI0/XI0_5/d_5_ DECAP_INV_G11
XG10421 XI11_3/XI0/XI0_5/d__4_ XI11_3/XI0/XI0_5/d_4_ DECAP_INV_G11
XG10422 XI11_3/XI0/XI0_5/d__3_ XI11_3/XI0/XI0_5/d_3_ DECAP_INV_G11
XG10423 XI11_3/XI0/XI0_5/d__2_ XI11_3/XI0/XI0_5/d_2_ DECAP_INV_G11
XG10424 XI11_3/XI0/XI0_5/d__1_ XI11_3/XI0/XI0_5/d_1_ DECAP_INV_G11
XG10425 XI11_3/XI0/XI0_5/d__0_ XI11_3/XI0/XI0_5/d_0_ DECAP_INV_G11
XG10426 XI11_3/XI0/XI0_5/d_15_ XI11_3/XI0/XI0_5/d__15_ DECAP_INV_G11
XG10427 XI11_3/XI0/XI0_5/d_14_ XI11_3/XI0/XI0_5/d__14_ DECAP_INV_G11
XG10428 XI11_3/XI0/XI0_5/d_13_ XI11_3/XI0/XI0_5/d__13_ DECAP_INV_G11
XG10429 XI11_3/XI0/XI0_5/d_12_ XI11_3/XI0/XI0_5/d__12_ DECAP_INV_G11
XG10430 XI11_3/XI0/XI0_5/d_11_ XI11_3/XI0/XI0_5/d__11_ DECAP_INV_G11
XG10431 XI11_3/XI0/XI0_5/d_10_ XI11_3/XI0/XI0_5/d__10_ DECAP_INV_G11
XG10432 XI11_3/XI0/XI0_5/d_9_ XI11_3/XI0/XI0_5/d__9_ DECAP_INV_G11
XG10433 XI11_3/XI0/XI0_5/d_8_ XI11_3/XI0/XI0_5/d__8_ DECAP_INV_G11
XG10434 XI11_3/XI0/XI0_5/d_7_ XI11_3/XI0/XI0_5/d__7_ DECAP_INV_G11
XG10435 XI11_3/XI0/XI0_5/d_6_ XI11_3/XI0/XI0_5/d__6_ DECAP_INV_G11
XG10436 XI11_3/XI0/XI0_5/d_5_ XI11_3/XI0/XI0_5/d__5_ DECAP_INV_G11
XG10437 XI11_3/XI0/XI0_5/d_4_ XI11_3/XI0/XI0_5/d__4_ DECAP_INV_G11
XG10438 XI11_3/XI0/XI0_5/d_3_ XI11_3/XI0/XI0_5/d__3_ DECAP_INV_G11
XG10439 XI11_3/XI0/XI0_5/d_2_ XI11_3/XI0/XI0_5/d__2_ DECAP_INV_G11
XG10440 XI11_3/XI0/XI0_5/d_1_ XI11_3/XI0/XI0_5/d__1_ DECAP_INV_G11
XG10441 XI11_3/XI0/XI0_5/d_0_ XI11_3/XI0/XI0_5/d__0_ DECAP_INV_G11
XG10442 XI11_3/XI0/XI0_4/d__15_ XI11_3/XI0/XI0_4/d_15_ DECAP_INV_G11
XG10443 XI11_3/XI0/XI0_4/d__14_ XI11_3/XI0/XI0_4/d_14_ DECAP_INV_G11
XG10444 XI11_3/XI0/XI0_4/d__13_ XI11_3/XI0/XI0_4/d_13_ DECAP_INV_G11
XG10445 XI11_3/XI0/XI0_4/d__12_ XI11_3/XI0/XI0_4/d_12_ DECAP_INV_G11
XG10446 XI11_3/XI0/XI0_4/d__11_ XI11_3/XI0/XI0_4/d_11_ DECAP_INV_G11
XG10447 XI11_3/XI0/XI0_4/d__10_ XI11_3/XI0/XI0_4/d_10_ DECAP_INV_G11
XG10448 XI11_3/XI0/XI0_4/d__9_ XI11_3/XI0/XI0_4/d_9_ DECAP_INV_G11
XG10449 XI11_3/XI0/XI0_4/d__8_ XI11_3/XI0/XI0_4/d_8_ DECAP_INV_G11
XG10450 XI11_3/XI0/XI0_4/d__7_ XI11_3/XI0/XI0_4/d_7_ DECAP_INV_G11
XG10451 XI11_3/XI0/XI0_4/d__6_ XI11_3/XI0/XI0_4/d_6_ DECAP_INV_G11
XG10452 XI11_3/XI0/XI0_4/d__5_ XI11_3/XI0/XI0_4/d_5_ DECAP_INV_G11
XG10453 XI11_3/XI0/XI0_4/d__4_ XI11_3/XI0/XI0_4/d_4_ DECAP_INV_G11
XG10454 XI11_3/XI0/XI0_4/d__3_ XI11_3/XI0/XI0_4/d_3_ DECAP_INV_G11
XG10455 XI11_3/XI0/XI0_4/d__2_ XI11_3/XI0/XI0_4/d_2_ DECAP_INV_G11
XG10456 XI11_3/XI0/XI0_4/d__1_ XI11_3/XI0/XI0_4/d_1_ DECAP_INV_G11
XG10457 XI11_3/XI0/XI0_4/d__0_ XI11_3/XI0/XI0_4/d_0_ DECAP_INV_G11
XG10458 XI11_3/XI0/XI0_4/d_15_ XI11_3/XI0/XI0_4/d__15_ DECAP_INV_G11
XG10459 XI11_3/XI0/XI0_4/d_14_ XI11_3/XI0/XI0_4/d__14_ DECAP_INV_G11
XG10460 XI11_3/XI0/XI0_4/d_13_ XI11_3/XI0/XI0_4/d__13_ DECAP_INV_G11
XG10461 XI11_3/XI0/XI0_4/d_12_ XI11_3/XI0/XI0_4/d__12_ DECAP_INV_G11
XG10462 XI11_3/XI0/XI0_4/d_11_ XI11_3/XI0/XI0_4/d__11_ DECAP_INV_G11
XG10463 XI11_3/XI0/XI0_4/d_10_ XI11_3/XI0/XI0_4/d__10_ DECAP_INV_G11
XG10464 XI11_3/XI0/XI0_4/d_9_ XI11_3/XI0/XI0_4/d__9_ DECAP_INV_G11
XG10465 XI11_3/XI0/XI0_4/d_8_ XI11_3/XI0/XI0_4/d__8_ DECAP_INV_G11
XG10466 XI11_3/XI0/XI0_4/d_7_ XI11_3/XI0/XI0_4/d__7_ DECAP_INV_G11
XG10467 XI11_3/XI0/XI0_4/d_6_ XI11_3/XI0/XI0_4/d__6_ DECAP_INV_G11
XG10468 XI11_3/XI0/XI0_4/d_5_ XI11_3/XI0/XI0_4/d__5_ DECAP_INV_G11
XG10469 XI11_3/XI0/XI0_4/d_4_ XI11_3/XI0/XI0_4/d__4_ DECAP_INV_G11
XG10470 XI11_3/XI0/XI0_4/d_3_ XI11_3/XI0/XI0_4/d__3_ DECAP_INV_G11
XG10471 XI11_3/XI0/XI0_4/d_2_ XI11_3/XI0/XI0_4/d__2_ DECAP_INV_G11
XG10472 XI11_3/XI0/XI0_4/d_1_ XI11_3/XI0/XI0_4/d__1_ DECAP_INV_G11
XG10473 XI11_3/XI0/XI0_4/d_0_ XI11_3/XI0/XI0_4/d__0_ DECAP_INV_G11
XG10474 XI11_3/XI0/XI0_3/d__15_ XI11_3/XI0/XI0_3/d_15_ DECAP_INV_G11
XG10475 XI11_3/XI0/XI0_3/d__14_ XI11_3/XI0/XI0_3/d_14_ DECAP_INV_G11
XG10476 XI11_3/XI0/XI0_3/d__13_ XI11_3/XI0/XI0_3/d_13_ DECAP_INV_G11
XG10477 XI11_3/XI0/XI0_3/d__12_ XI11_3/XI0/XI0_3/d_12_ DECAP_INV_G11
XG10478 XI11_3/XI0/XI0_3/d__11_ XI11_3/XI0/XI0_3/d_11_ DECAP_INV_G11
XG10479 XI11_3/XI0/XI0_3/d__10_ XI11_3/XI0/XI0_3/d_10_ DECAP_INV_G11
XG10480 XI11_3/XI0/XI0_3/d__9_ XI11_3/XI0/XI0_3/d_9_ DECAP_INV_G11
XG10481 XI11_3/XI0/XI0_3/d__8_ XI11_3/XI0/XI0_3/d_8_ DECAP_INV_G11
XG10482 XI11_3/XI0/XI0_3/d__7_ XI11_3/XI0/XI0_3/d_7_ DECAP_INV_G11
XG10483 XI11_3/XI0/XI0_3/d__6_ XI11_3/XI0/XI0_3/d_6_ DECAP_INV_G11
XG10484 XI11_3/XI0/XI0_3/d__5_ XI11_3/XI0/XI0_3/d_5_ DECAP_INV_G11
XG10485 XI11_3/XI0/XI0_3/d__4_ XI11_3/XI0/XI0_3/d_4_ DECAP_INV_G11
XG10486 XI11_3/XI0/XI0_3/d__3_ XI11_3/XI0/XI0_3/d_3_ DECAP_INV_G11
XG10487 XI11_3/XI0/XI0_3/d__2_ XI11_3/XI0/XI0_3/d_2_ DECAP_INV_G11
XG10488 XI11_3/XI0/XI0_3/d__1_ XI11_3/XI0/XI0_3/d_1_ DECAP_INV_G11
XG10489 XI11_3/XI0/XI0_3/d__0_ XI11_3/XI0/XI0_3/d_0_ DECAP_INV_G11
XG10490 XI11_3/XI0/XI0_3/d_15_ XI11_3/XI0/XI0_3/d__15_ DECAP_INV_G11
XG10491 XI11_3/XI0/XI0_3/d_14_ XI11_3/XI0/XI0_3/d__14_ DECAP_INV_G11
XG10492 XI11_3/XI0/XI0_3/d_13_ XI11_3/XI0/XI0_3/d__13_ DECAP_INV_G11
XG10493 XI11_3/XI0/XI0_3/d_12_ XI11_3/XI0/XI0_3/d__12_ DECAP_INV_G11
XG10494 XI11_3/XI0/XI0_3/d_11_ XI11_3/XI0/XI0_3/d__11_ DECAP_INV_G11
XG10495 XI11_3/XI0/XI0_3/d_10_ XI11_3/XI0/XI0_3/d__10_ DECAP_INV_G11
XG10496 XI11_3/XI0/XI0_3/d_9_ XI11_3/XI0/XI0_3/d__9_ DECAP_INV_G11
XG10497 XI11_3/XI0/XI0_3/d_8_ XI11_3/XI0/XI0_3/d__8_ DECAP_INV_G11
XG10498 XI11_3/XI0/XI0_3/d_7_ XI11_3/XI0/XI0_3/d__7_ DECAP_INV_G11
XG10499 XI11_3/XI0/XI0_3/d_6_ XI11_3/XI0/XI0_3/d__6_ DECAP_INV_G11
XG10500 XI11_3/XI0/XI0_3/d_5_ XI11_3/XI0/XI0_3/d__5_ DECAP_INV_G11
XG10501 XI11_3/XI0/XI0_3/d_4_ XI11_3/XI0/XI0_3/d__4_ DECAP_INV_G11
XG10502 XI11_3/XI0/XI0_3/d_3_ XI11_3/XI0/XI0_3/d__3_ DECAP_INV_G11
XG10503 XI11_3/XI0/XI0_3/d_2_ XI11_3/XI0/XI0_3/d__2_ DECAP_INV_G11
XG10504 XI11_3/XI0/XI0_3/d_1_ XI11_3/XI0/XI0_3/d__1_ DECAP_INV_G11
XG10505 XI11_3/XI0/XI0_3/d_0_ XI11_3/XI0/XI0_3/d__0_ DECAP_INV_G11
XG10506 XI11_3/XI0/XI0_2/d__15_ XI11_3/XI0/XI0_2/d_15_ DECAP_INV_G11
XG10507 XI11_3/XI0/XI0_2/d__14_ XI11_3/XI0/XI0_2/d_14_ DECAP_INV_G11
XG10508 XI11_3/XI0/XI0_2/d__13_ XI11_3/XI0/XI0_2/d_13_ DECAP_INV_G11
XG10509 XI11_3/XI0/XI0_2/d__12_ XI11_3/XI0/XI0_2/d_12_ DECAP_INV_G11
XG10510 XI11_3/XI0/XI0_2/d__11_ XI11_3/XI0/XI0_2/d_11_ DECAP_INV_G11
XG10511 XI11_3/XI0/XI0_2/d__10_ XI11_3/XI0/XI0_2/d_10_ DECAP_INV_G11
XG10512 XI11_3/XI0/XI0_2/d__9_ XI11_3/XI0/XI0_2/d_9_ DECAP_INV_G11
XG10513 XI11_3/XI0/XI0_2/d__8_ XI11_3/XI0/XI0_2/d_8_ DECAP_INV_G11
XG10514 XI11_3/XI0/XI0_2/d__7_ XI11_3/XI0/XI0_2/d_7_ DECAP_INV_G11
XG10515 XI11_3/XI0/XI0_2/d__6_ XI11_3/XI0/XI0_2/d_6_ DECAP_INV_G11
XG10516 XI11_3/XI0/XI0_2/d__5_ XI11_3/XI0/XI0_2/d_5_ DECAP_INV_G11
XG10517 XI11_3/XI0/XI0_2/d__4_ XI11_3/XI0/XI0_2/d_4_ DECAP_INV_G11
XG10518 XI11_3/XI0/XI0_2/d__3_ XI11_3/XI0/XI0_2/d_3_ DECAP_INV_G11
XG10519 XI11_3/XI0/XI0_2/d__2_ XI11_3/XI0/XI0_2/d_2_ DECAP_INV_G11
XG10520 XI11_3/XI0/XI0_2/d__1_ XI11_3/XI0/XI0_2/d_1_ DECAP_INV_G11
XG10521 XI11_3/XI0/XI0_2/d__0_ XI11_3/XI0/XI0_2/d_0_ DECAP_INV_G11
XG10522 XI11_3/XI0/XI0_2/d_15_ XI11_3/XI0/XI0_2/d__15_ DECAP_INV_G11
XG10523 XI11_3/XI0/XI0_2/d_14_ XI11_3/XI0/XI0_2/d__14_ DECAP_INV_G11
XG10524 XI11_3/XI0/XI0_2/d_13_ XI11_3/XI0/XI0_2/d__13_ DECAP_INV_G11
XG10525 XI11_3/XI0/XI0_2/d_12_ XI11_3/XI0/XI0_2/d__12_ DECAP_INV_G11
XG10526 XI11_3/XI0/XI0_2/d_11_ XI11_3/XI0/XI0_2/d__11_ DECAP_INV_G11
XG10527 XI11_3/XI0/XI0_2/d_10_ XI11_3/XI0/XI0_2/d__10_ DECAP_INV_G11
XG10528 XI11_3/XI0/XI0_2/d_9_ XI11_3/XI0/XI0_2/d__9_ DECAP_INV_G11
XG10529 XI11_3/XI0/XI0_2/d_8_ XI11_3/XI0/XI0_2/d__8_ DECAP_INV_G11
XG10530 XI11_3/XI0/XI0_2/d_7_ XI11_3/XI0/XI0_2/d__7_ DECAP_INV_G11
XG10531 XI11_3/XI0/XI0_2/d_6_ XI11_3/XI0/XI0_2/d__6_ DECAP_INV_G11
XG10532 XI11_3/XI0/XI0_2/d_5_ XI11_3/XI0/XI0_2/d__5_ DECAP_INV_G11
XG10533 XI11_3/XI0/XI0_2/d_4_ XI11_3/XI0/XI0_2/d__4_ DECAP_INV_G11
XG10534 XI11_3/XI0/XI0_2/d_3_ XI11_3/XI0/XI0_2/d__3_ DECAP_INV_G11
XG10535 XI11_3/XI0/XI0_2/d_2_ XI11_3/XI0/XI0_2/d__2_ DECAP_INV_G11
XG10536 XI11_3/XI0/XI0_2/d_1_ XI11_3/XI0/XI0_2/d__1_ DECAP_INV_G11
XG10537 XI11_3/XI0/XI0_2/d_0_ XI11_3/XI0/XI0_2/d__0_ DECAP_INV_G11
XG10538 XI11_3/XI0/XI0_1/d__15_ XI11_3/XI0/XI0_1/d_15_ DECAP_INV_G11
XG10539 XI11_3/XI0/XI0_1/d__14_ XI11_3/XI0/XI0_1/d_14_ DECAP_INV_G11
XG10540 XI11_3/XI0/XI0_1/d__13_ XI11_3/XI0/XI0_1/d_13_ DECAP_INV_G11
XG10541 XI11_3/XI0/XI0_1/d__12_ XI11_3/XI0/XI0_1/d_12_ DECAP_INV_G11
XG10542 XI11_3/XI0/XI0_1/d__11_ XI11_3/XI0/XI0_1/d_11_ DECAP_INV_G11
XG10543 XI11_3/XI0/XI0_1/d__10_ XI11_3/XI0/XI0_1/d_10_ DECAP_INV_G11
XG10544 XI11_3/XI0/XI0_1/d__9_ XI11_3/XI0/XI0_1/d_9_ DECAP_INV_G11
XG10545 XI11_3/XI0/XI0_1/d__8_ XI11_3/XI0/XI0_1/d_8_ DECAP_INV_G11
XG10546 XI11_3/XI0/XI0_1/d__7_ XI11_3/XI0/XI0_1/d_7_ DECAP_INV_G11
XG10547 XI11_3/XI0/XI0_1/d__6_ XI11_3/XI0/XI0_1/d_6_ DECAP_INV_G11
XG10548 XI11_3/XI0/XI0_1/d__5_ XI11_3/XI0/XI0_1/d_5_ DECAP_INV_G11
XG10549 XI11_3/XI0/XI0_1/d__4_ XI11_3/XI0/XI0_1/d_4_ DECAP_INV_G11
XG10550 XI11_3/XI0/XI0_1/d__3_ XI11_3/XI0/XI0_1/d_3_ DECAP_INV_G11
XG10551 XI11_3/XI0/XI0_1/d__2_ XI11_3/XI0/XI0_1/d_2_ DECAP_INV_G11
XG10552 XI11_3/XI0/XI0_1/d__1_ XI11_3/XI0/XI0_1/d_1_ DECAP_INV_G11
XG10553 XI11_3/XI0/XI0_1/d__0_ XI11_3/XI0/XI0_1/d_0_ DECAP_INV_G11
XG10554 XI11_3/XI0/XI0_1/d_15_ XI11_3/XI0/XI0_1/d__15_ DECAP_INV_G11
XG10555 XI11_3/XI0/XI0_1/d_14_ XI11_3/XI0/XI0_1/d__14_ DECAP_INV_G11
XG10556 XI11_3/XI0/XI0_1/d_13_ XI11_3/XI0/XI0_1/d__13_ DECAP_INV_G11
XG10557 XI11_3/XI0/XI0_1/d_12_ XI11_3/XI0/XI0_1/d__12_ DECAP_INV_G11
XG10558 XI11_3/XI0/XI0_1/d_11_ XI11_3/XI0/XI0_1/d__11_ DECAP_INV_G11
XG10559 XI11_3/XI0/XI0_1/d_10_ XI11_3/XI0/XI0_1/d__10_ DECAP_INV_G11
XG10560 XI11_3/XI0/XI0_1/d_9_ XI11_3/XI0/XI0_1/d__9_ DECAP_INV_G11
XG10561 XI11_3/XI0/XI0_1/d_8_ XI11_3/XI0/XI0_1/d__8_ DECAP_INV_G11
XG10562 XI11_3/XI0/XI0_1/d_7_ XI11_3/XI0/XI0_1/d__7_ DECAP_INV_G11
XG10563 XI11_3/XI0/XI0_1/d_6_ XI11_3/XI0/XI0_1/d__6_ DECAP_INV_G11
XG10564 XI11_3/XI0/XI0_1/d_5_ XI11_3/XI0/XI0_1/d__5_ DECAP_INV_G11
XG10565 XI11_3/XI0/XI0_1/d_4_ XI11_3/XI0/XI0_1/d__4_ DECAP_INV_G11
XG10566 XI11_3/XI0/XI0_1/d_3_ XI11_3/XI0/XI0_1/d__3_ DECAP_INV_G11
XG10567 XI11_3/XI0/XI0_1/d_2_ XI11_3/XI0/XI0_1/d__2_ DECAP_INV_G11
XG10568 XI11_3/XI0/XI0_1/d_1_ XI11_3/XI0/XI0_1/d__1_ DECAP_INV_G11
XG10569 XI11_3/XI0/XI0_1/d_0_ XI11_3/XI0/XI0_1/d__0_ DECAP_INV_G11
XG10570 XI11_3/XI0/XI0_0/d__15_ XI11_3/XI0/XI0_0/d_15_ DECAP_INV_G11
XG10571 XI11_3/XI0/XI0_0/d__14_ XI11_3/XI0/XI0_0/d_14_ DECAP_INV_G11
XG10572 XI11_3/XI0/XI0_0/d__13_ XI11_3/XI0/XI0_0/d_13_ DECAP_INV_G11
XG10573 XI11_3/XI0/XI0_0/d__12_ XI11_3/XI0/XI0_0/d_12_ DECAP_INV_G11
XG10574 XI11_3/XI0/XI0_0/d__11_ XI11_3/XI0/XI0_0/d_11_ DECAP_INV_G11
XG10575 XI11_3/XI0/XI0_0/d__10_ XI11_3/XI0/XI0_0/d_10_ DECAP_INV_G11
XG10576 XI11_3/XI0/XI0_0/d__9_ XI11_3/XI0/XI0_0/d_9_ DECAP_INV_G11
XG10577 XI11_3/XI0/XI0_0/d__8_ XI11_3/XI0/XI0_0/d_8_ DECAP_INV_G11
XG10578 XI11_3/XI0/XI0_0/d__7_ XI11_3/XI0/XI0_0/d_7_ DECAP_INV_G11
XG10579 XI11_3/XI0/XI0_0/d__6_ XI11_3/XI0/XI0_0/d_6_ DECAP_INV_G11
XG10580 XI11_3/XI0/XI0_0/d__5_ XI11_3/XI0/XI0_0/d_5_ DECAP_INV_G11
XG10581 XI11_3/XI0/XI0_0/d__4_ XI11_3/XI0/XI0_0/d_4_ DECAP_INV_G11
XG10582 XI11_3/XI0/XI0_0/d__3_ XI11_3/XI0/XI0_0/d_3_ DECAP_INV_G11
XG10583 XI11_3/XI0/XI0_0/d__2_ XI11_3/XI0/XI0_0/d_2_ DECAP_INV_G11
XG10584 XI11_3/XI0/XI0_0/d__1_ XI11_3/XI0/XI0_0/d_1_ DECAP_INV_G11
XG10585 XI11_3/XI0/XI0_0/d__0_ XI11_3/XI0/XI0_0/d_0_ DECAP_INV_G11
XG10586 XI11_3/XI0/XI0_0/d_15_ XI11_3/XI0/XI0_0/d__15_ DECAP_INV_G11
XG10587 XI11_3/XI0/XI0_0/d_14_ XI11_3/XI0/XI0_0/d__14_ DECAP_INV_G11
XG10588 XI11_3/XI0/XI0_0/d_13_ XI11_3/XI0/XI0_0/d__13_ DECAP_INV_G11
XG10589 XI11_3/XI0/XI0_0/d_12_ XI11_3/XI0/XI0_0/d__12_ DECAP_INV_G11
XG10590 XI11_3/XI0/XI0_0/d_11_ XI11_3/XI0/XI0_0/d__11_ DECAP_INV_G11
XG10591 XI11_3/XI0/XI0_0/d_10_ XI11_3/XI0/XI0_0/d__10_ DECAP_INV_G11
XG10592 XI11_3/XI0/XI0_0/d_9_ XI11_3/XI0/XI0_0/d__9_ DECAP_INV_G11
XG10593 XI11_3/XI0/XI0_0/d_8_ XI11_3/XI0/XI0_0/d__8_ DECAP_INV_G11
XG10594 XI11_3/XI0/XI0_0/d_7_ XI11_3/XI0/XI0_0/d__7_ DECAP_INV_G11
XG10595 XI11_3/XI0/XI0_0/d_6_ XI11_3/XI0/XI0_0/d__6_ DECAP_INV_G11
XG10596 XI11_3/XI0/XI0_0/d_5_ XI11_3/XI0/XI0_0/d__5_ DECAP_INV_G11
XG10597 XI11_3/XI0/XI0_0/d_4_ XI11_3/XI0/XI0_0/d__4_ DECAP_INV_G11
XG10598 XI11_3/XI0/XI0_0/d_3_ XI11_3/XI0/XI0_0/d__3_ DECAP_INV_G11
XG10599 XI11_3/XI0/XI0_0/d_2_ XI11_3/XI0/XI0_0/d__2_ DECAP_INV_G11
XG10600 XI11_3/XI0/XI0_0/d_1_ XI11_3/XI0/XI0_0/d__1_ DECAP_INV_G11
XG10601 XI11_3/XI0/XI0_0/d_0_ XI11_3/XI0/XI0_0/d__0_ DECAP_INV_G11
XG10602 XI11_2/XI3/net17 XI11_2/XI3/net5 DECAP_INV_G7
XG10603 XI11_2/XI3/net5 XI11_2/preck DECAP_INV_G8
XG10604 sck_bar XI11_2/XI3/net018 DECAP_INV_G9
XG10605 XI11_2/XI3/net018 XI11_2/XI3/net012 DECAP_INV_G9
XG10606 XI11_2/XI3/net014 XI11_2/XI3/net7 DECAP_INV_G9
XG10607 XI11_2/XI3/net012 XI11_2/XI3/net014 DECAP_INV_G9
XG10608 XI11_2/XI4/net063 XI11_2/XI4/net0112 DECAP_INV_G10
XG10609 XI11_2/XI4/net26 XI11_2/XI4/net089 DECAP_INV_G10
XG10610 XI11_2/XI4/data_out XI11_2/XI4/data_out_ DECAP_INV_G10
XG10611 XI11_2/XI4/net20 XI11_2/XI4/net0103 DECAP_INV_G10
XG10612 XI11_2/net12 XI11_2/XI4/net32 DECAP_INV_G7
XG10613 XI11_2/net9 XI11_2/XI4/net52 DECAP_INV_G7
XG10614 XI11_2/XI4/data_out_ XI11_2/XI4/data_out DECAP_INV_G10
XG10615 XI11_2/XI0/XI0_63/d__15_ XI11_2/XI0/XI0_63/d_15_ DECAP_INV_G11
XG10616 XI11_2/XI0/XI0_63/d__14_ XI11_2/XI0/XI0_63/d_14_ DECAP_INV_G11
XG10617 XI11_2/XI0/XI0_63/d__13_ XI11_2/XI0/XI0_63/d_13_ DECAP_INV_G11
XG10618 XI11_2/XI0/XI0_63/d__12_ XI11_2/XI0/XI0_63/d_12_ DECAP_INV_G11
XG10619 XI11_2/XI0/XI0_63/d__11_ XI11_2/XI0/XI0_63/d_11_ DECAP_INV_G11
XG10620 XI11_2/XI0/XI0_63/d__10_ XI11_2/XI0/XI0_63/d_10_ DECAP_INV_G11
XG10621 XI11_2/XI0/XI0_63/d__9_ XI11_2/XI0/XI0_63/d_9_ DECAP_INV_G11
XG10622 XI11_2/XI0/XI0_63/d__8_ XI11_2/XI0/XI0_63/d_8_ DECAP_INV_G11
XG10623 XI11_2/XI0/XI0_63/d__7_ XI11_2/XI0/XI0_63/d_7_ DECAP_INV_G11
XG10624 XI11_2/XI0/XI0_63/d__6_ XI11_2/XI0/XI0_63/d_6_ DECAP_INV_G11
XG10625 XI11_2/XI0/XI0_63/d__5_ XI11_2/XI0/XI0_63/d_5_ DECAP_INV_G11
XG10626 XI11_2/XI0/XI0_63/d__4_ XI11_2/XI0/XI0_63/d_4_ DECAP_INV_G11
XG10627 XI11_2/XI0/XI0_63/d__3_ XI11_2/XI0/XI0_63/d_3_ DECAP_INV_G11
XG10628 XI11_2/XI0/XI0_63/d__2_ XI11_2/XI0/XI0_63/d_2_ DECAP_INV_G11
XG10629 XI11_2/XI0/XI0_63/d__1_ XI11_2/XI0/XI0_63/d_1_ DECAP_INV_G11
XG10630 XI11_2/XI0/XI0_63/d__0_ XI11_2/XI0/XI0_63/d_0_ DECAP_INV_G11
XG10631 XI11_2/XI0/XI0_63/d_15_ XI11_2/XI0/XI0_63/d__15_ DECAP_INV_G11
XG10632 XI11_2/XI0/XI0_63/d_14_ XI11_2/XI0/XI0_63/d__14_ DECAP_INV_G11
XG10633 XI11_2/XI0/XI0_63/d_13_ XI11_2/XI0/XI0_63/d__13_ DECAP_INV_G11
XG10634 XI11_2/XI0/XI0_63/d_12_ XI11_2/XI0/XI0_63/d__12_ DECAP_INV_G11
XG10635 XI11_2/XI0/XI0_63/d_11_ XI11_2/XI0/XI0_63/d__11_ DECAP_INV_G11
XG10636 XI11_2/XI0/XI0_63/d_10_ XI11_2/XI0/XI0_63/d__10_ DECAP_INV_G11
XG10637 XI11_2/XI0/XI0_63/d_9_ XI11_2/XI0/XI0_63/d__9_ DECAP_INV_G11
XG10638 XI11_2/XI0/XI0_63/d_8_ XI11_2/XI0/XI0_63/d__8_ DECAP_INV_G11
XG10639 XI11_2/XI0/XI0_63/d_7_ XI11_2/XI0/XI0_63/d__7_ DECAP_INV_G11
XG10640 XI11_2/XI0/XI0_63/d_6_ XI11_2/XI0/XI0_63/d__6_ DECAP_INV_G11
XG10641 XI11_2/XI0/XI0_63/d_5_ XI11_2/XI0/XI0_63/d__5_ DECAP_INV_G11
XG10642 XI11_2/XI0/XI0_63/d_4_ XI11_2/XI0/XI0_63/d__4_ DECAP_INV_G11
XG10643 XI11_2/XI0/XI0_63/d_3_ XI11_2/XI0/XI0_63/d__3_ DECAP_INV_G11
XG10644 XI11_2/XI0/XI0_63/d_2_ XI11_2/XI0/XI0_63/d__2_ DECAP_INV_G11
XG10645 XI11_2/XI0/XI0_63/d_1_ XI11_2/XI0/XI0_63/d__1_ DECAP_INV_G11
XG10646 XI11_2/XI0/XI0_63/d_0_ XI11_2/XI0/XI0_63/d__0_ DECAP_INV_G11
XG10647 XI11_2/XI0/XI0_62/d__15_ XI11_2/XI0/XI0_62/d_15_ DECAP_INV_G11
XG10648 XI11_2/XI0/XI0_62/d__14_ XI11_2/XI0/XI0_62/d_14_ DECAP_INV_G11
XG10649 XI11_2/XI0/XI0_62/d__13_ XI11_2/XI0/XI0_62/d_13_ DECAP_INV_G11
XG10650 XI11_2/XI0/XI0_62/d__12_ XI11_2/XI0/XI0_62/d_12_ DECAP_INV_G11
XG10651 XI11_2/XI0/XI0_62/d__11_ XI11_2/XI0/XI0_62/d_11_ DECAP_INV_G11
XG10652 XI11_2/XI0/XI0_62/d__10_ XI11_2/XI0/XI0_62/d_10_ DECAP_INV_G11
XG10653 XI11_2/XI0/XI0_62/d__9_ XI11_2/XI0/XI0_62/d_9_ DECAP_INV_G11
XG10654 XI11_2/XI0/XI0_62/d__8_ XI11_2/XI0/XI0_62/d_8_ DECAP_INV_G11
XG10655 XI11_2/XI0/XI0_62/d__7_ XI11_2/XI0/XI0_62/d_7_ DECAP_INV_G11
XG10656 XI11_2/XI0/XI0_62/d__6_ XI11_2/XI0/XI0_62/d_6_ DECAP_INV_G11
XG10657 XI11_2/XI0/XI0_62/d__5_ XI11_2/XI0/XI0_62/d_5_ DECAP_INV_G11
XG10658 XI11_2/XI0/XI0_62/d__4_ XI11_2/XI0/XI0_62/d_4_ DECAP_INV_G11
XG10659 XI11_2/XI0/XI0_62/d__3_ XI11_2/XI0/XI0_62/d_3_ DECAP_INV_G11
XG10660 XI11_2/XI0/XI0_62/d__2_ XI11_2/XI0/XI0_62/d_2_ DECAP_INV_G11
XG10661 XI11_2/XI0/XI0_62/d__1_ XI11_2/XI0/XI0_62/d_1_ DECAP_INV_G11
XG10662 XI11_2/XI0/XI0_62/d__0_ XI11_2/XI0/XI0_62/d_0_ DECAP_INV_G11
XG10663 XI11_2/XI0/XI0_62/d_15_ XI11_2/XI0/XI0_62/d__15_ DECAP_INV_G11
XG10664 XI11_2/XI0/XI0_62/d_14_ XI11_2/XI0/XI0_62/d__14_ DECAP_INV_G11
XG10665 XI11_2/XI0/XI0_62/d_13_ XI11_2/XI0/XI0_62/d__13_ DECAP_INV_G11
XG10666 XI11_2/XI0/XI0_62/d_12_ XI11_2/XI0/XI0_62/d__12_ DECAP_INV_G11
XG10667 XI11_2/XI0/XI0_62/d_11_ XI11_2/XI0/XI0_62/d__11_ DECAP_INV_G11
XG10668 XI11_2/XI0/XI0_62/d_10_ XI11_2/XI0/XI0_62/d__10_ DECAP_INV_G11
XG10669 XI11_2/XI0/XI0_62/d_9_ XI11_2/XI0/XI0_62/d__9_ DECAP_INV_G11
XG10670 XI11_2/XI0/XI0_62/d_8_ XI11_2/XI0/XI0_62/d__8_ DECAP_INV_G11
XG10671 XI11_2/XI0/XI0_62/d_7_ XI11_2/XI0/XI0_62/d__7_ DECAP_INV_G11
XG10672 XI11_2/XI0/XI0_62/d_6_ XI11_2/XI0/XI0_62/d__6_ DECAP_INV_G11
XG10673 XI11_2/XI0/XI0_62/d_5_ XI11_2/XI0/XI0_62/d__5_ DECAP_INV_G11
XG10674 XI11_2/XI0/XI0_62/d_4_ XI11_2/XI0/XI0_62/d__4_ DECAP_INV_G11
XG10675 XI11_2/XI0/XI0_62/d_3_ XI11_2/XI0/XI0_62/d__3_ DECAP_INV_G11
XG10676 XI11_2/XI0/XI0_62/d_2_ XI11_2/XI0/XI0_62/d__2_ DECAP_INV_G11
XG10677 XI11_2/XI0/XI0_62/d_1_ XI11_2/XI0/XI0_62/d__1_ DECAP_INV_G11
XG10678 XI11_2/XI0/XI0_62/d_0_ XI11_2/XI0/XI0_62/d__0_ DECAP_INV_G11
XG10679 XI11_2/XI0/XI0_61/d__15_ XI11_2/XI0/XI0_61/d_15_ DECAP_INV_G11
XG10680 XI11_2/XI0/XI0_61/d__14_ XI11_2/XI0/XI0_61/d_14_ DECAP_INV_G11
XG10681 XI11_2/XI0/XI0_61/d__13_ XI11_2/XI0/XI0_61/d_13_ DECAP_INV_G11
XG10682 XI11_2/XI0/XI0_61/d__12_ XI11_2/XI0/XI0_61/d_12_ DECAP_INV_G11
XG10683 XI11_2/XI0/XI0_61/d__11_ XI11_2/XI0/XI0_61/d_11_ DECAP_INV_G11
XG10684 XI11_2/XI0/XI0_61/d__10_ XI11_2/XI0/XI0_61/d_10_ DECAP_INV_G11
XG10685 XI11_2/XI0/XI0_61/d__9_ XI11_2/XI0/XI0_61/d_9_ DECAP_INV_G11
XG10686 XI11_2/XI0/XI0_61/d__8_ XI11_2/XI0/XI0_61/d_8_ DECAP_INV_G11
XG10687 XI11_2/XI0/XI0_61/d__7_ XI11_2/XI0/XI0_61/d_7_ DECAP_INV_G11
XG10688 XI11_2/XI0/XI0_61/d__6_ XI11_2/XI0/XI0_61/d_6_ DECAP_INV_G11
XG10689 XI11_2/XI0/XI0_61/d__5_ XI11_2/XI0/XI0_61/d_5_ DECAP_INV_G11
XG10690 XI11_2/XI0/XI0_61/d__4_ XI11_2/XI0/XI0_61/d_4_ DECAP_INV_G11
XG10691 XI11_2/XI0/XI0_61/d__3_ XI11_2/XI0/XI0_61/d_3_ DECAP_INV_G11
XG10692 XI11_2/XI0/XI0_61/d__2_ XI11_2/XI0/XI0_61/d_2_ DECAP_INV_G11
XG10693 XI11_2/XI0/XI0_61/d__1_ XI11_2/XI0/XI0_61/d_1_ DECAP_INV_G11
XG10694 XI11_2/XI0/XI0_61/d__0_ XI11_2/XI0/XI0_61/d_0_ DECAP_INV_G11
XG10695 XI11_2/XI0/XI0_61/d_15_ XI11_2/XI0/XI0_61/d__15_ DECAP_INV_G11
XG10696 XI11_2/XI0/XI0_61/d_14_ XI11_2/XI0/XI0_61/d__14_ DECAP_INV_G11
XG10697 XI11_2/XI0/XI0_61/d_13_ XI11_2/XI0/XI0_61/d__13_ DECAP_INV_G11
XG10698 XI11_2/XI0/XI0_61/d_12_ XI11_2/XI0/XI0_61/d__12_ DECAP_INV_G11
XG10699 XI11_2/XI0/XI0_61/d_11_ XI11_2/XI0/XI0_61/d__11_ DECAP_INV_G11
XG10700 XI11_2/XI0/XI0_61/d_10_ XI11_2/XI0/XI0_61/d__10_ DECAP_INV_G11
XG10701 XI11_2/XI0/XI0_61/d_9_ XI11_2/XI0/XI0_61/d__9_ DECAP_INV_G11
XG10702 XI11_2/XI0/XI0_61/d_8_ XI11_2/XI0/XI0_61/d__8_ DECAP_INV_G11
XG10703 XI11_2/XI0/XI0_61/d_7_ XI11_2/XI0/XI0_61/d__7_ DECAP_INV_G11
XG10704 XI11_2/XI0/XI0_61/d_6_ XI11_2/XI0/XI0_61/d__6_ DECAP_INV_G11
XG10705 XI11_2/XI0/XI0_61/d_5_ XI11_2/XI0/XI0_61/d__5_ DECAP_INV_G11
XG10706 XI11_2/XI0/XI0_61/d_4_ XI11_2/XI0/XI0_61/d__4_ DECAP_INV_G11
XG10707 XI11_2/XI0/XI0_61/d_3_ XI11_2/XI0/XI0_61/d__3_ DECAP_INV_G11
XG10708 XI11_2/XI0/XI0_61/d_2_ XI11_2/XI0/XI0_61/d__2_ DECAP_INV_G11
XG10709 XI11_2/XI0/XI0_61/d_1_ XI11_2/XI0/XI0_61/d__1_ DECAP_INV_G11
XG10710 XI11_2/XI0/XI0_61/d_0_ XI11_2/XI0/XI0_61/d__0_ DECAP_INV_G11
XG10711 XI11_2/XI0/XI0_60/d__15_ XI11_2/XI0/XI0_60/d_15_ DECAP_INV_G11
XG10712 XI11_2/XI0/XI0_60/d__14_ XI11_2/XI0/XI0_60/d_14_ DECAP_INV_G11
XG10713 XI11_2/XI0/XI0_60/d__13_ XI11_2/XI0/XI0_60/d_13_ DECAP_INV_G11
XG10714 XI11_2/XI0/XI0_60/d__12_ XI11_2/XI0/XI0_60/d_12_ DECAP_INV_G11
XG10715 XI11_2/XI0/XI0_60/d__11_ XI11_2/XI0/XI0_60/d_11_ DECAP_INV_G11
XG10716 XI11_2/XI0/XI0_60/d__10_ XI11_2/XI0/XI0_60/d_10_ DECAP_INV_G11
XG10717 XI11_2/XI0/XI0_60/d__9_ XI11_2/XI0/XI0_60/d_9_ DECAP_INV_G11
XG10718 XI11_2/XI0/XI0_60/d__8_ XI11_2/XI0/XI0_60/d_8_ DECAP_INV_G11
XG10719 XI11_2/XI0/XI0_60/d__7_ XI11_2/XI0/XI0_60/d_7_ DECAP_INV_G11
XG10720 XI11_2/XI0/XI0_60/d__6_ XI11_2/XI0/XI0_60/d_6_ DECAP_INV_G11
XG10721 XI11_2/XI0/XI0_60/d__5_ XI11_2/XI0/XI0_60/d_5_ DECAP_INV_G11
XG10722 XI11_2/XI0/XI0_60/d__4_ XI11_2/XI0/XI0_60/d_4_ DECAP_INV_G11
XG10723 XI11_2/XI0/XI0_60/d__3_ XI11_2/XI0/XI0_60/d_3_ DECAP_INV_G11
XG10724 XI11_2/XI0/XI0_60/d__2_ XI11_2/XI0/XI0_60/d_2_ DECAP_INV_G11
XG10725 XI11_2/XI0/XI0_60/d__1_ XI11_2/XI0/XI0_60/d_1_ DECAP_INV_G11
XG10726 XI11_2/XI0/XI0_60/d__0_ XI11_2/XI0/XI0_60/d_0_ DECAP_INV_G11
XG10727 XI11_2/XI0/XI0_60/d_15_ XI11_2/XI0/XI0_60/d__15_ DECAP_INV_G11
XG10728 XI11_2/XI0/XI0_60/d_14_ XI11_2/XI0/XI0_60/d__14_ DECAP_INV_G11
XG10729 XI11_2/XI0/XI0_60/d_13_ XI11_2/XI0/XI0_60/d__13_ DECAP_INV_G11
XG10730 XI11_2/XI0/XI0_60/d_12_ XI11_2/XI0/XI0_60/d__12_ DECAP_INV_G11
XG10731 XI11_2/XI0/XI0_60/d_11_ XI11_2/XI0/XI0_60/d__11_ DECAP_INV_G11
XG10732 XI11_2/XI0/XI0_60/d_10_ XI11_2/XI0/XI0_60/d__10_ DECAP_INV_G11
XG10733 XI11_2/XI0/XI0_60/d_9_ XI11_2/XI0/XI0_60/d__9_ DECAP_INV_G11
XG10734 XI11_2/XI0/XI0_60/d_8_ XI11_2/XI0/XI0_60/d__8_ DECAP_INV_G11
XG10735 XI11_2/XI0/XI0_60/d_7_ XI11_2/XI0/XI0_60/d__7_ DECAP_INV_G11
XG10736 XI11_2/XI0/XI0_60/d_6_ XI11_2/XI0/XI0_60/d__6_ DECAP_INV_G11
XG10737 XI11_2/XI0/XI0_60/d_5_ XI11_2/XI0/XI0_60/d__5_ DECAP_INV_G11
XG10738 XI11_2/XI0/XI0_60/d_4_ XI11_2/XI0/XI0_60/d__4_ DECAP_INV_G11
XG10739 XI11_2/XI0/XI0_60/d_3_ XI11_2/XI0/XI0_60/d__3_ DECAP_INV_G11
XG10740 XI11_2/XI0/XI0_60/d_2_ XI11_2/XI0/XI0_60/d__2_ DECAP_INV_G11
XG10741 XI11_2/XI0/XI0_60/d_1_ XI11_2/XI0/XI0_60/d__1_ DECAP_INV_G11
XG10742 XI11_2/XI0/XI0_60/d_0_ XI11_2/XI0/XI0_60/d__0_ DECAP_INV_G11
XG10743 XI11_2/XI0/XI0_59/d__15_ XI11_2/XI0/XI0_59/d_15_ DECAP_INV_G11
XG10744 XI11_2/XI0/XI0_59/d__14_ XI11_2/XI0/XI0_59/d_14_ DECAP_INV_G11
XG10745 XI11_2/XI0/XI0_59/d__13_ XI11_2/XI0/XI0_59/d_13_ DECAP_INV_G11
XG10746 XI11_2/XI0/XI0_59/d__12_ XI11_2/XI0/XI0_59/d_12_ DECAP_INV_G11
XG10747 XI11_2/XI0/XI0_59/d__11_ XI11_2/XI0/XI0_59/d_11_ DECAP_INV_G11
XG10748 XI11_2/XI0/XI0_59/d__10_ XI11_2/XI0/XI0_59/d_10_ DECAP_INV_G11
XG10749 XI11_2/XI0/XI0_59/d__9_ XI11_2/XI0/XI0_59/d_9_ DECAP_INV_G11
XG10750 XI11_2/XI0/XI0_59/d__8_ XI11_2/XI0/XI0_59/d_8_ DECAP_INV_G11
XG10751 XI11_2/XI0/XI0_59/d__7_ XI11_2/XI0/XI0_59/d_7_ DECAP_INV_G11
XG10752 XI11_2/XI0/XI0_59/d__6_ XI11_2/XI0/XI0_59/d_6_ DECAP_INV_G11
XG10753 XI11_2/XI0/XI0_59/d__5_ XI11_2/XI0/XI0_59/d_5_ DECAP_INV_G11
XG10754 XI11_2/XI0/XI0_59/d__4_ XI11_2/XI0/XI0_59/d_4_ DECAP_INV_G11
XG10755 XI11_2/XI0/XI0_59/d__3_ XI11_2/XI0/XI0_59/d_3_ DECAP_INV_G11
XG10756 XI11_2/XI0/XI0_59/d__2_ XI11_2/XI0/XI0_59/d_2_ DECAP_INV_G11
XG10757 XI11_2/XI0/XI0_59/d__1_ XI11_2/XI0/XI0_59/d_1_ DECAP_INV_G11
XG10758 XI11_2/XI0/XI0_59/d__0_ XI11_2/XI0/XI0_59/d_0_ DECAP_INV_G11
XG10759 XI11_2/XI0/XI0_59/d_15_ XI11_2/XI0/XI0_59/d__15_ DECAP_INV_G11
XG10760 XI11_2/XI0/XI0_59/d_14_ XI11_2/XI0/XI0_59/d__14_ DECAP_INV_G11
XG10761 XI11_2/XI0/XI0_59/d_13_ XI11_2/XI0/XI0_59/d__13_ DECAP_INV_G11
XG10762 XI11_2/XI0/XI0_59/d_12_ XI11_2/XI0/XI0_59/d__12_ DECAP_INV_G11
XG10763 XI11_2/XI0/XI0_59/d_11_ XI11_2/XI0/XI0_59/d__11_ DECAP_INV_G11
XG10764 XI11_2/XI0/XI0_59/d_10_ XI11_2/XI0/XI0_59/d__10_ DECAP_INV_G11
XG10765 XI11_2/XI0/XI0_59/d_9_ XI11_2/XI0/XI0_59/d__9_ DECAP_INV_G11
XG10766 XI11_2/XI0/XI0_59/d_8_ XI11_2/XI0/XI0_59/d__8_ DECAP_INV_G11
XG10767 XI11_2/XI0/XI0_59/d_7_ XI11_2/XI0/XI0_59/d__7_ DECAP_INV_G11
XG10768 XI11_2/XI0/XI0_59/d_6_ XI11_2/XI0/XI0_59/d__6_ DECAP_INV_G11
XG10769 XI11_2/XI0/XI0_59/d_5_ XI11_2/XI0/XI0_59/d__5_ DECAP_INV_G11
XG10770 XI11_2/XI0/XI0_59/d_4_ XI11_2/XI0/XI0_59/d__4_ DECAP_INV_G11
XG10771 XI11_2/XI0/XI0_59/d_3_ XI11_2/XI0/XI0_59/d__3_ DECAP_INV_G11
XG10772 XI11_2/XI0/XI0_59/d_2_ XI11_2/XI0/XI0_59/d__2_ DECAP_INV_G11
XG10773 XI11_2/XI0/XI0_59/d_1_ XI11_2/XI0/XI0_59/d__1_ DECAP_INV_G11
XG10774 XI11_2/XI0/XI0_59/d_0_ XI11_2/XI0/XI0_59/d__0_ DECAP_INV_G11
XG10775 XI11_2/XI0/XI0_58/d__15_ XI11_2/XI0/XI0_58/d_15_ DECAP_INV_G11
XG10776 XI11_2/XI0/XI0_58/d__14_ XI11_2/XI0/XI0_58/d_14_ DECAP_INV_G11
XG10777 XI11_2/XI0/XI0_58/d__13_ XI11_2/XI0/XI0_58/d_13_ DECAP_INV_G11
XG10778 XI11_2/XI0/XI0_58/d__12_ XI11_2/XI0/XI0_58/d_12_ DECAP_INV_G11
XG10779 XI11_2/XI0/XI0_58/d__11_ XI11_2/XI0/XI0_58/d_11_ DECAP_INV_G11
XG10780 XI11_2/XI0/XI0_58/d__10_ XI11_2/XI0/XI0_58/d_10_ DECAP_INV_G11
XG10781 XI11_2/XI0/XI0_58/d__9_ XI11_2/XI0/XI0_58/d_9_ DECAP_INV_G11
XG10782 XI11_2/XI0/XI0_58/d__8_ XI11_2/XI0/XI0_58/d_8_ DECAP_INV_G11
XG10783 XI11_2/XI0/XI0_58/d__7_ XI11_2/XI0/XI0_58/d_7_ DECAP_INV_G11
XG10784 XI11_2/XI0/XI0_58/d__6_ XI11_2/XI0/XI0_58/d_6_ DECAP_INV_G11
XG10785 XI11_2/XI0/XI0_58/d__5_ XI11_2/XI0/XI0_58/d_5_ DECAP_INV_G11
XG10786 XI11_2/XI0/XI0_58/d__4_ XI11_2/XI0/XI0_58/d_4_ DECAP_INV_G11
XG10787 XI11_2/XI0/XI0_58/d__3_ XI11_2/XI0/XI0_58/d_3_ DECAP_INV_G11
XG10788 XI11_2/XI0/XI0_58/d__2_ XI11_2/XI0/XI0_58/d_2_ DECAP_INV_G11
XG10789 XI11_2/XI0/XI0_58/d__1_ XI11_2/XI0/XI0_58/d_1_ DECAP_INV_G11
XG10790 XI11_2/XI0/XI0_58/d__0_ XI11_2/XI0/XI0_58/d_0_ DECAP_INV_G11
XG10791 XI11_2/XI0/XI0_58/d_15_ XI11_2/XI0/XI0_58/d__15_ DECAP_INV_G11
XG10792 XI11_2/XI0/XI0_58/d_14_ XI11_2/XI0/XI0_58/d__14_ DECAP_INV_G11
XG10793 XI11_2/XI0/XI0_58/d_13_ XI11_2/XI0/XI0_58/d__13_ DECAP_INV_G11
XG10794 XI11_2/XI0/XI0_58/d_12_ XI11_2/XI0/XI0_58/d__12_ DECAP_INV_G11
XG10795 XI11_2/XI0/XI0_58/d_11_ XI11_2/XI0/XI0_58/d__11_ DECAP_INV_G11
XG10796 XI11_2/XI0/XI0_58/d_10_ XI11_2/XI0/XI0_58/d__10_ DECAP_INV_G11
XG10797 XI11_2/XI0/XI0_58/d_9_ XI11_2/XI0/XI0_58/d__9_ DECAP_INV_G11
XG10798 XI11_2/XI0/XI0_58/d_8_ XI11_2/XI0/XI0_58/d__8_ DECAP_INV_G11
XG10799 XI11_2/XI0/XI0_58/d_7_ XI11_2/XI0/XI0_58/d__7_ DECAP_INV_G11
XG10800 XI11_2/XI0/XI0_58/d_6_ XI11_2/XI0/XI0_58/d__6_ DECAP_INV_G11
XG10801 XI11_2/XI0/XI0_58/d_5_ XI11_2/XI0/XI0_58/d__5_ DECAP_INV_G11
XG10802 XI11_2/XI0/XI0_58/d_4_ XI11_2/XI0/XI0_58/d__4_ DECAP_INV_G11
XG10803 XI11_2/XI0/XI0_58/d_3_ XI11_2/XI0/XI0_58/d__3_ DECAP_INV_G11
XG10804 XI11_2/XI0/XI0_58/d_2_ XI11_2/XI0/XI0_58/d__2_ DECAP_INV_G11
XG10805 XI11_2/XI0/XI0_58/d_1_ XI11_2/XI0/XI0_58/d__1_ DECAP_INV_G11
XG10806 XI11_2/XI0/XI0_58/d_0_ XI11_2/XI0/XI0_58/d__0_ DECAP_INV_G11
XG10807 XI11_2/XI0/XI0_57/d__15_ XI11_2/XI0/XI0_57/d_15_ DECAP_INV_G11
XG10808 XI11_2/XI0/XI0_57/d__14_ XI11_2/XI0/XI0_57/d_14_ DECAP_INV_G11
XG10809 XI11_2/XI0/XI0_57/d__13_ XI11_2/XI0/XI0_57/d_13_ DECAP_INV_G11
XG10810 XI11_2/XI0/XI0_57/d__12_ XI11_2/XI0/XI0_57/d_12_ DECAP_INV_G11
XG10811 XI11_2/XI0/XI0_57/d__11_ XI11_2/XI0/XI0_57/d_11_ DECAP_INV_G11
XG10812 XI11_2/XI0/XI0_57/d__10_ XI11_2/XI0/XI0_57/d_10_ DECAP_INV_G11
XG10813 XI11_2/XI0/XI0_57/d__9_ XI11_2/XI0/XI0_57/d_9_ DECAP_INV_G11
XG10814 XI11_2/XI0/XI0_57/d__8_ XI11_2/XI0/XI0_57/d_8_ DECAP_INV_G11
XG10815 XI11_2/XI0/XI0_57/d__7_ XI11_2/XI0/XI0_57/d_7_ DECAP_INV_G11
XG10816 XI11_2/XI0/XI0_57/d__6_ XI11_2/XI0/XI0_57/d_6_ DECAP_INV_G11
XG10817 XI11_2/XI0/XI0_57/d__5_ XI11_2/XI0/XI0_57/d_5_ DECAP_INV_G11
XG10818 XI11_2/XI0/XI0_57/d__4_ XI11_2/XI0/XI0_57/d_4_ DECAP_INV_G11
XG10819 XI11_2/XI0/XI0_57/d__3_ XI11_2/XI0/XI0_57/d_3_ DECAP_INV_G11
XG10820 XI11_2/XI0/XI0_57/d__2_ XI11_2/XI0/XI0_57/d_2_ DECAP_INV_G11
XG10821 XI11_2/XI0/XI0_57/d__1_ XI11_2/XI0/XI0_57/d_1_ DECAP_INV_G11
XG10822 XI11_2/XI0/XI0_57/d__0_ XI11_2/XI0/XI0_57/d_0_ DECAP_INV_G11
XG10823 XI11_2/XI0/XI0_57/d_15_ XI11_2/XI0/XI0_57/d__15_ DECAP_INV_G11
XG10824 XI11_2/XI0/XI0_57/d_14_ XI11_2/XI0/XI0_57/d__14_ DECAP_INV_G11
XG10825 XI11_2/XI0/XI0_57/d_13_ XI11_2/XI0/XI0_57/d__13_ DECAP_INV_G11
XG10826 XI11_2/XI0/XI0_57/d_12_ XI11_2/XI0/XI0_57/d__12_ DECAP_INV_G11
XG10827 XI11_2/XI0/XI0_57/d_11_ XI11_2/XI0/XI0_57/d__11_ DECAP_INV_G11
XG10828 XI11_2/XI0/XI0_57/d_10_ XI11_2/XI0/XI0_57/d__10_ DECAP_INV_G11
XG10829 XI11_2/XI0/XI0_57/d_9_ XI11_2/XI0/XI0_57/d__9_ DECAP_INV_G11
XG10830 XI11_2/XI0/XI0_57/d_8_ XI11_2/XI0/XI0_57/d__8_ DECAP_INV_G11
XG10831 XI11_2/XI0/XI0_57/d_7_ XI11_2/XI0/XI0_57/d__7_ DECAP_INV_G11
XG10832 XI11_2/XI0/XI0_57/d_6_ XI11_2/XI0/XI0_57/d__6_ DECAP_INV_G11
XG10833 XI11_2/XI0/XI0_57/d_5_ XI11_2/XI0/XI0_57/d__5_ DECAP_INV_G11
XG10834 XI11_2/XI0/XI0_57/d_4_ XI11_2/XI0/XI0_57/d__4_ DECAP_INV_G11
XG10835 XI11_2/XI0/XI0_57/d_3_ XI11_2/XI0/XI0_57/d__3_ DECAP_INV_G11
XG10836 XI11_2/XI0/XI0_57/d_2_ XI11_2/XI0/XI0_57/d__2_ DECAP_INV_G11
XG10837 XI11_2/XI0/XI0_57/d_1_ XI11_2/XI0/XI0_57/d__1_ DECAP_INV_G11
XG10838 XI11_2/XI0/XI0_57/d_0_ XI11_2/XI0/XI0_57/d__0_ DECAP_INV_G11
XG10839 XI11_2/XI0/XI0_56/d__15_ XI11_2/XI0/XI0_56/d_15_ DECAP_INV_G11
XG10840 XI11_2/XI0/XI0_56/d__14_ XI11_2/XI0/XI0_56/d_14_ DECAP_INV_G11
XG10841 XI11_2/XI0/XI0_56/d__13_ XI11_2/XI0/XI0_56/d_13_ DECAP_INV_G11
XG10842 XI11_2/XI0/XI0_56/d__12_ XI11_2/XI0/XI0_56/d_12_ DECAP_INV_G11
XG10843 XI11_2/XI0/XI0_56/d__11_ XI11_2/XI0/XI0_56/d_11_ DECAP_INV_G11
XG10844 XI11_2/XI0/XI0_56/d__10_ XI11_2/XI0/XI0_56/d_10_ DECAP_INV_G11
XG10845 XI11_2/XI0/XI0_56/d__9_ XI11_2/XI0/XI0_56/d_9_ DECAP_INV_G11
XG10846 XI11_2/XI0/XI0_56/d__8_ XI11_2/XI0/XI0_56/d_8_ DECAP_INV_G11
XG10847 XI11_2/XI0/XI0_56/d__7_ XI11_2/XI0/XI0_56/d_7_ DECAP_INV_G11
XG10848 XI11_2/XI0/XI0_56/d__6_ XI11_2/XI0/XI0_56/d_6_ DECAP_INV_G11
XG10849 XI11_2/XI0/XI0_56/d__5_ XI11_2/XI0/XI0_56/d_5_ DECAP_INV_G11
XG10850 XI11_2/XI0/XI0_56/d__4_ XI11_2/XI0/XI0_56/d_4_ DECAP_INV_G11
XG10851 XI11_2/XI0/XI0_56/d__3_ XI11_2/XI0/XI0_56/d_3_ DECAP_INV_G11
XG10852 XI11_2/XI0/XI0_56/d__2_ XI11_2/XI0/XI0_56/d_2_ DECAP_INV_G11
XG10853 XI11_2/XI0/XI0_56/d__1_ XI11_2/XI0/XI0_56/d_1_ DECAP_INV_G11
XG10854 XI11_2/XI0/XI0_56/d__0_ XI11_2/XI0/XI0_56/d_0_ DECAP_INV_G11
XG10855 XI11_2/XI0/XI0_56/d_15_ XI11_2/XI0/XI0_56/d__15_ DECAP_INV_G11
XG10856 XI11_2/XI0/XI0_56/d_14_ XI11_2/XI0/XI0_56/d__14_ DECAP_INV_G11
XG10857 XI11_2/XI0/XI0_56/d_13_ XI11_2/XI0/XI0_56/d__13_ DECAP_INV_G11
XG10858 XI11_2/XI0/XI0_56/d_12_ XI11_2/XI0/XI0_56/d__12_ DECAP_INV_G11
XG10859 XI11_2/XI0/XI0_56/d_11_ XI11_2/XI0/XI0_56/d__11_ DECAP_INV_G11
XG10860 XI11_2/XI0/XI0_56/d_10_ XI11_2/XI0/XI0_56/d__10_ DECAP_INV_G11
XG10861 XI11_2/XI0/XI0_56/d_9_ XI11_2/XI0/XI0_56/d__9_ DECAP_INV_G11
XG10862 XI11_2/XI0/XI0_56/d_8_ XI11_2/XI0/XI0_56/d__8_ DECAP_INV_G11
XG10863 XI11_2/XI0/XI0_56/d_7_ XI11_2/XI0/XI0_56/d__7_ DECAP_INV_G11
XG10864 XI11_2/XI0/XI0_56/d_6_ XI11_2/XI0/XI0_56/d__6_ DECAP_INV_G11
XG10865 XI11_2/XI0/XI0_56/d_5_ XI11_2/XI0/XI0_56/d__5_ DECAP_INV_G11
XG10866 XI11_2/XI0/XI0_56/d_4_ XI11_2/XI0/XI0_56/d__4_ DECAP_INV_G11
XG10867 XI11_2/XI0/XI0_56/d_3_ XI11_2/XI0/XI0_56/d__3_ DECAP_INV_G11
XG10868 XI11_2/XI0/XI0_56/d_2_ XI11_2/XI0/XI0_56/d__2_ DECAP_INV_G11
XG10869 XI11_2/XI0/XI0_56/d_1_ XI11_2/XI0/XI0_56/d__1_ DECAP_INV_G11
XG10870 XI11_2/XI0/XI0_56/d_0_ XI11_2/XI0/XI0_56/d__0_ DECAP_INV_G11
XG10871 XI11_2/XI0/XI0_55/d__15_ XI11_2/XI0/XI0_55/d_15_ DECAP_INV_G11
XG10872 XI11_2/XI0/XI0_55/d__14_ XI11_2/XI0/XI0_55/d_14_ DECAP_INV_G11
XG10873 XI11_2/XI0/XI0_55/d__13_ XI11_2/XI0/XI0_55/d_13_ DECAP_INV_G11
XG10874 XI11_2/XI0/XI0_55/d__12_ XI11_2/XI0/XI0_55/d_12_ DECAP_INV_G11
XG10875 XI11_2/XI0/XI0_55/d__11_ XI11_2/XI0/XI0_55/d_11_ DECAP_INV_G11
XG10876 XI11_2/XI0/XI0_55/d__10_ XI11_2/XI0/XI0_55/d_10_ DECAP_INV_G11
XG10877 XI11_2/XI0/XI0_55/d__9_ XI11_2/XI0/XI0_55/d_9_ DECAP_INV_G11
XG10878 XI11_2/XI0/XI0_55/d__8_ XI11_2/XI0/XI0_55/d_8_ DECAP_INV_G11
XG10879 XI11_2/XI0/XI0_55/d__7_ XI11_2/XI0/XI0_55/d_7_ DECAP_INV_G11
XG10880 XI11_2/XI0/XI0_55/d__6_ XI11_2/XI0/XI0_55/d_6_ DECAP_INV_G11
XG10881 XI11_2/XI0/XI0_55/d__5_ XI11_2/XI0/XI0_55/d_5_ DECAP_INV_G11
XG10882 XI11_2/XI0/XI0_55/d__4_ XI11_2/XI0/XI0_55/d_4_ DECAP_INV_G11
XG10883 XI11_2/XI0/XI0_55/d__3_ XI11_2/XI0/XI0_55/d_3_ DECAP_INV_G11
XG10884 XI11_2/XI0/XI0_55/d__2_ XI11_2/XI0/XI0_55/d_2_ DECAP_INV_G11
XG10885 XI11_2/XI0/XI0_55/d__1_ XI11_2/XI0/XI0_55/d_1_ DECAP_INV_G11
XG10886 XI11_2/XI0/XI0_55/d__0_ XI11_2/XI0/XI0_55/d_0_ DECAP_INV_G11
XG10887 XI11_2/XI0/XI0_55/d_15_ XI11_2/XI0/XI0_55/d__15_ DECAP_INV_G11
XG10888 XI11_2/XI0/XI0_55/d_14_ XI11_2/XI0/XI0_55/d__14_ DECAP_INV_G11
XG10889 XI11_2/XI0/XI0_55/d_13_ XI11_2/XI0/XI0_55/d__13_ DECAP_INV_G11
XG10890 XI11_2/XI0/XI0_55/d_12_ XI11_2/XI0/XI0_55/d__12_ DECAP_INV_G11
XG10891 XI11_2/XI0/XI0_55/d_11_ XI11_2/XI0/XI0_55/d__11_ DECAP_INV_G11
XG10892 XI11_2/XI0/XI0_55/d_10_ XI11_2/XI0/XI0_55/d__10_ DECAP_INV_G11
XG10893 XI11_2/XI0/XI0_55/d_9_ XI11_2/XI0/XI0_55/d__9_ DECAP_INV_G11
XG10894 XI11_2/XI0/XI0_55/d_8_ XI11_2/XI0/XI0_55/d__8_ DECAP_INV_G11
XG10895 XI11_2/XI0/XI0_55/d_7_ XI11_2/XI0/XI0_55/d__7_ DECAP_INV_G11
XG10896 XI11_2/XI0/XI0_55/d_6_ XI11_2/XI0/XI0_55/d__6_ DECAP_INV_G11
XG10897 XI11_2/XI0/XI0_55/d_5_ XI11_2/XI0/XI0_55/d__5_ DECAP_INV_G11
XG10898 XI11_2/XI0/XI0_55/d_4_ XI11_2/XI0/XI0_55/d__4_ DECAP_INV_G11
XG10899 XI11_2/XI0/XI0_55/d_3_ XI11_2/XI0/XI0_55/d__3_ DECAP_INV_G11
XG10900 XI11_2/XI0/XI0_55/d_2_ XI11_2/XI0/XI0_55/d__2_ DECAP_INV_G11
XG10901 XI11_2/XI0/XI0_55/d_1_ XI11_2/XI0/XI0_55/d__1_ DECAP_INV_G11
XG10902 XI11_2/XI0/XI0_55/d_0_ XI11_2/XI0/XI0_55/d__0_ DECAP_INV_G11
XG10903 XI11_2/XI0/XI0_54/d__15_ XI11_2/XI0/XI0_54/d_15_ DECAP_INV_G11
XG10904 XI11_2/XI0/XI0_54/d__14_ XI11_2/XI0/XI0_54/d_14_ DECAP_INV_G11
XG10905 XI11_2/XI0/XI0_54/d__13_ XI11_2/XI0/XI0_54/d_13_ DECAP_INV_G11
XG10906 XI11_2/XI0/XI0_54/d__12_ XI11_2/XI0/XI0_54/d_12_ DECAP_INV_G11
XG10907 XI11_2/XI0/XI0_54/d__11_ XI11_2/XI0/XI0_54/d_11_ DECAP_INV_G11
XG10908 XI11_2/XI0/XI0_54/d__10_ XI11_2/XI0/XI0_54/d_10_ DECAP_INV_G11
XG10909 XI11_2/XI0/XI0_54/d__9_ XI11_2/XI0/XI0_54/d_9_ DECAP_INV_G11
XG10910 XI11_2/XI0/XI0_54/d__8_ XI11_2/XI0/XI0_54/d_8_ DECAP_INV_G11
XG10911 XI11_2/XI0/XI0_54/d__7_ XI11_2/XI0/XI0_54/d_7_ DECAP_INV_G11
XG10912 XI11_2/XI0/XI0_54/d__6_ XI11_2/XI0/XI0_54/d_6_ DECAP_INV_G11
XG10913 XI11_2/XI0/XI0_54/d__5_ XI11_2/XI0/XI0_54/d_5_ DECAP_INV_G11
XG10914 XI11_2/XI0/XI0_54/d__4_ XI11_2/XI0/XI0_54/d_4_ DECAP_INV_G11
XG10915 XI11_2/XI0/XI0_54/d__3_ XI11_2/XI0/XI0_54/d_3_ DECAP_INV_G11
XG10916 XI11_2/XI0/XI0_54/d__2_ XI11_2/XI0/XI0_54/d_2_ DECAP_INV_G11
XG10917 XI11_2/XI0/XI0_54/d__1_ XI11_2/XI0/XI0_54/d_1_ DECAP_INV_G11
XG10918 XI11_2/XI0/XI0_54/d__0_ XI11_2/XI0/XI0_54/d_0_ DECAP_INV_G11
XG10919 XI11_2/XI0/XI0_54/d_15_ XI11_2/XI0/XI0_54/d__15_ DECAP_INV_G11
XG10920 XI11_2/XI0/XI0_54/d_14_ XI11_2/XI0/XI0_54/d__14_ DECAP_INV_G11
XG10921 XI11_2/XI0/XI0_54/d_13_ XI11_2/XI0/XI0_54/d__13_ DECAP_INV_G11
XG10922 XI11_2/XI0/XI0_54/d_12_ XI11_2/XI0/XI0_54/d__12_ DECAP_INV_G11
XG10923 XI11_2/XI0/XI0_54/d_11_ XI11_2/XI0/XI0_54/d__11_ DECAP_INV_G11
XG10924 XI11_2/XI0/XI0_54/d_10_ XI11_2/XI0/XI0_54/d__10_ DECAP_INV_G11
XG10925 XI11_2/XI0/XI0_54/d_9_ XI11_2/XI0/XI0_54/d__9_ DECAP_INV_G11
XG10926 XI11_2/XI0/XI0_54/d_8_ XI11_2/XI0/XI0_54/d__8_ DECAP_INV_G11
XG10927 XI11_2/XI0/XI0_54/d_7_ XI11_2/XI0/XI0_54/d__7_ DECAP_INV_G11
XG10928 XI11_2/XI0/XI0_54/d_6_ XI11_2/XI0/XI0_54/d__6_ DECAP_INV_G11
XG10929 XI11_2/XI0/XI0_54/d_5_ XI11_2/XI0/XI0_54/d__5_ DECAP_INV_G11
XG10930 XI11_2/XI0/XI0_54/d_4_ XI11_2/XI0/XI0_54/d__4_ DECAP_INV_G11
XG10931 XI11_2/XI0/XI0_54/d_3_ XI11_2/XI0/XI0_54/d__3_ DECAP_INV_G11
XG10932 XI11_2/XI0/XI0_54/d_2_ XI11_2/XI0/XI0_54/d__2_ DECAP_INV_G11
XG10933 XI11_2/XI0/XI0_54/d_1_ XI11_2/XI0/XI0_54/d__1_ DECAP_INV_G11
XG10934 XI11_2/XI0/XI0_54/d_0_ XI11_2/XI0/XI0_54/d__0_ DECAP_INV_G11
XG10935 XI11_2/XI0/XI0_53/d__15_ XI11_2/XI0/XI0_53/d_15_ DECAP_INV_G11
XG10936 XI11_2/XI0/XI0_53/d__14_ XI11_2/XI0/XI0_53/d_14_ DECAP_INV_G11
XG10937 XI11_2/XI0/XI0_53/d__13_ XI11_2/XI0/XI0_53/d_13_ DECAP_INV_G11
XG10938 XI11_2/XI0/XI0_53/d__12_ XI11_2/XI0/XI0_53/d_12_ DECAP_INV_G11
XG10939 XI11_2/XI0/XI0_53/d__11_ XI11_2/XI0/XI0_53/d_11_ DECAP_INV_G11
XG10940 XI11_2/XI0/XI0_53/d__10_ XI11_2/XI0/XI0_53/d_10_ DECAP_INV_G11
XG10941 XI11_2/XI0/XI0_53/d__9_ XI11_2/XI0/XI0_53/d_9_ DECAP_INV_G11
XG10942 XI11_2/XI0/XI0_53/d__8_ XI11_2/XI0/XI0_53/d_8_ DECAP_INV_G11
XG10943 XI11_2/XI0/XI0_53/d__7_ XI11_2/XI0/XI0_53/d_7_ DECAP_INV_G11
XG10944 XI11_2/XI0/XI0_53/d__6_ XI11_2/XI0/XI0_53/d_6_ DECAP_INV_G11
XG10945 XI11_2/XI0/XI0_53/d__5_ XI11_2/XI0/XI0_53/d_5_ DECAP_INV_G11
XG10946 XI11_2/XI0/XI0_53/d__4_ XI11_2/XI0/XI0_53/d_4_ DECAP_INV_G11
XG10947 XI11_2/XI0/XI0_53/d__3_ XI11_2/XI0/XI0_53/d_3_ DECAP_INV_G11
XG10948 XI11_2/XI0/XI0_53/d__2_ XI11_2/XI0/XI0_53/d_2_ DECAP_INV_G11
XG10949 XI11_2/XI0/XI0_53/d__1_ XI11_2/XI0/XI0_53/d_1_ DECAP_INV_G11
XG10950 XI11_2/XI0/XI0_53/d__0_ XI11_2/XI0/XI0_53/d_0_ DECAP_INV_G11
XG10951 XI11_2/XI0/XI0_53/d_15_ XI11_2/XI0/XI0_53/d__15_ DECAP_INV_G11
XG10952 XI11_2/XI0/XI0_53/d_14_ XI11_2/XI0/XI0_53/d__14_ DECAP_INV_G11
XG10953 XI11_2/XI0/XI0_53/d_13_ XI11_2/XI0/XI0_53/d__13_ DECAP_INV_G11
XG10954 XI11_2/XI0/XI0_53/d_12_ XI11_2/XI0/XI0_53/d__12_ DECAP_INV_G11
XG10955 XI11_2/XI0/XI0_53/d_11_ XI11_2/XI0/XI0_53/d__11_ DECAP_INV_G11
XG10956 XI11_2/XI0/XI0_53/d_10_ XI11_2/XI0/XI0_53/d__10_ DECAP_INV_G11
XG10957 XI11_2/XI0/XI0_53/d_9_ XI11_2/XI0/XI0_53/d__9_ DECAP_INV_G11
XG10958 XI11_2/XI0/XI0_53/d_8_ XI11_2/XI0/XI0_53/d__8_ DECAP_INV_G11
XG10959 XI11_2/XI0/XI0_53/d_7_ XI11_2/XI0/XI0_53/d__7_ DECAP_INV_G11
XG10960 XI11_2/XI0/XI0_53/d_6_ XI11_2/XI0/XI0_53/d__6_ DECAP_INV_G11
XG10961 XI11_2/XI0/XI0_53/d_5_ XI11_2/XI0/XI0_53/d__5_ DECAP_INV_G11
XG10962 XI11_2/XI0/XI0_53/d_4_ XI11_2/XI0/XI0_53/d__4_ DECAP_INV_G11
XG10963 XI11_2/XI0/XI0_53/d_3_ XI11_2/XI0/XI0_53/d__3_ DECAP_INV_G11
XG10964 XI11_2/XI0/XI0_53/d_2_ XI11_2/XI0/XI0_53/d__2_ DECAP_INV_G11
XG10965 XI11_2/XI0/XI0_53/d_1_ XI11_2/XI0/XI0_53/d__1_ DECAP_INV_G11
XG10966 XI11_2/XI0/XI0_53/d_0_ XI11_2/XI0/XI0_53/d__0_ DECAP_INV_G11
XG10967 XI11_2/XI0/XI0_52/d__15_ XI11_2/XI0/XI0_52/d_15_ DECAP_INV_G11
XG10968 XI11_2/XI0/XI0_52/d__14_ XI11_2/XI0/XI0_52/d_14_ DECAP_INV_G11
XG10969 XI11_2/XI0/XI0_52/d__13_ XI11_2/XI0/XI0_52/d_13_ DECAP_INV_G11
XG10970 XI11_2/XI0/XI0_52/d__12_ XI11_2/XI0/XI0_52/d_12_ DECAP_INV_G11
XG10971 XI11_2/XI0/XI0_52/d__11_ XI11_2/XI0/XI0_52/d_11_ DECAP_INV_G11
XG10972 XI11_2/XI0/XI0_52/d__10_ XI11_2/XI0/XI0_52/d_10_ DECAP_INV_G11
XG10973 XI11_2/XI0/XI0_52/d__9_ XI11_2/XI0/XI0_52/d_9_ DECAP_INV_G11
XG10974 XI11_2/XI0/XI0_52/d__8_ XI11_2/XI0/XI0_52/d_8_ DECAP_INV_G11
XG10975 XI11_2/XI0/XI0_52/d__7_ XI11_2/XI0/XI0_52/d_7_ DECAP_INV_G11
XG10976 XI11_2/XI0/XI0_52/d__6_ XI11_2/XI0/XI0_52/d_6_ DECAP_INV_G11
XG10977 XI11_2/XI0/XI0_52/d__5_ XI11_2/XI0/XI0_52/d_5_ DECAP_INV_G11
XG10978 XI11_2/XI0/XI0_52/d__4_ XI11_2/XI0/XI0_52/d_4_ DECAP_INV_G11
XG10979 XI11_2/XI0/XI0_52/d__3_ XI11_2/XI0/XI0_52/d_3_ DECAP_INV_G11
XG10980 XI11_2/XI0/XI0_52/d__2_ XI11_2/XI0/XI0_52/d_2_ DECAP_INV_G11
XG10981 XI11_2/XI0/XI0_52/d__1_ XI11_2/XI0/XI0_52/d_1_ DECAP_INV_G11
XG10982 XI11_2/XI0/XI0_52/d__0_ XI11_2/XI0/XI0_52/d_0_ DECAP_INV_G11
XG10983 XI11_2/XI0/XI0_52/d_15_ XI11_2/XI0/XI0_52/d__15_ DECAP_INV_G11
XG10984 XI11_2/XI0/XI0_52/d_14_ XI11_2/XI0/XI0_52/d__14_ DECAP_INV_G11
XG10985 XI11_2/XI0/XI0_52/d_13_ XI11_2/XI0/XI0_52/d__13_ DECAP_INV_G11
XG10986 XI11_2/XI0/XI0_52/d_12_ XI11_2/XI0/XI0_52/d__12_ DECAP_INV_G11
XG10987 XI11_2/XI0/XI0_52/d_11_ XI11_2/XI0/XI0_52/d__11_ DECAP_INV_G11
XG10988 XI11_2/XI0/XI0_52/d_10_ XI11_2/XI0/XI0_52/d__10_ DECAP_INV_G11
XG10989 XI11_2/XI0/XI0_52/d_9_ XI11_2/XI0/XI0_52/d__9_ DECAP_INV_G11
XG10990 XI11_2/XI0/XI0_52/d_8_ XI11_2/XI0/XI0_52/d__8_ DECAP_INV_G11
XG10991 XI11_2/XI0/XI0_52/d_7_ XI11_2/XI0/XI0_52/d__7_ DECAP_INV_G11
XG10992 XI11_2/XI0/XI0_52/d_6_ XI11_2/XI0/XI0_52/d__6_ DECAP_INV_G11
XG10993 XI11_2/XI0/XI0_52/d_5_ XI11_2/XI0/XI0_52/d__5_ DECAP_INV_G11
XG10994 XI11_2/XI0/XI0_52/d_4_ XI11_2/XI0/XI0_52/d__4_ DECAP_INV_G11
XG10995 XI11_2/XI0/XI0_52/d_3_ XI11_2/XI0/XI0_52/d__3_ DECAP_INV_G11
XG10996 XI11_2/XI0/XI0_52/d_2_ XI11_2/XI0/XI0_52/d__2_ DECAP_INV_G11
XG10997 XI11_2/XI0/XI0_52/d_1_ XI11_2/XI0/XI0_52/d__1_ DECAP_INV_G11
XG10998 XI11_2/XI0/XI0_52/d_0_ XI11_2/XI0/XI0_52/d__0_ DECAP_INV_G11
XG10999 XI11_2/XI0/XI0_51/d__15_ XI11_2/XI0/XI0_51/d_15_ DECAP_INV_G11
XG11000 XI11_2/XI0/XI0_51/d__14_ XI11_2/XI0/XI0_51/d_14_ DECAP_INV_G11
XG11001 XI11_2/XI0/XI0_51/d__13_ XI11_2/XI0/XI0_51/d_13_ DECAP_INV_G11
XG11002 XI11_2/XI0/XI0_51/d__12_ XI11_2/XI0/XI0_51/d_12_ DECAP_INV_G11
XG11003 XI11_2/XI0/XI0_51/d__11_ XI11_2/XI0/XI0_51/d_11_ DECAP_INV_G11
XG11004 XI11_2/XI0/XI0_51/d__10_ XI11_2/XI0/XI0_51/d_10_ DECAP_INV_G11
XG11005 XI11_2/XI0/XI0_51/d__9_ XI11_2/XI0/XI0_51/d_9_ DECAP_INV_G11
XG11006 XI11_2/XI0/XI0_51/d__8_ XI11_2/XI0/XI0_51/d_8_ DECAP_INV_G11
XG11007 XI11_2/XI0/XI0_51/d__7_ XI11_2/XI0/XI0_51/d_7_ DECAP_INV_G11
XG11008 XI11_2/XI0/XI0_51/d__6_ XI11_2/XI0/XI0_51/d_6_ DECAP_INV_G11
XG11009 XI11_2/XI0/XI0_51/d__5_ XI11_2/XI0/XI0_51/d_5_ DECAP_INV_G11
XG11010 XI11_2/XI0/XI0_51/d__4_ XI11_2/XI0/XI0_51/d_4_ DECAP_INV_G11
XG11011 XI11_2/XI0/XI0_51/d__3_ XI11_2/XI0/XI0_51/d_3_ DECAP_INV_G11
XG11012 XI11_2/XI0/XI0_51/d__2_ XI11_2/XI0/XI0_51/d_2_ DECAP_INV_G11
XG11013 XI11_2/XI0/XI0_51/d__1_ XI11_2/XI0/XI0_51/d_1_ DECAP_INV_G11
XG11014 XI11_2/XI0/XI0_51/d__0_ XI11_2/XI0/XI0_51/d_0_ DECAP_INV_G11
XG11015 XI11_2/XI0/XI0_51/d_15_ XI11_2/XI0/XI0_51/d__15_ DECAP_INV_G11
XG11016 XI11_2/XI0/XI0_51/d_14_ XI11_2/XI0/XI0_51/d__14_ DECAP_INV_G11
XG11017 XI11_2/XI0/XI0_51/d_13_ XI11_2/XI0/XI0_51/d__13_ DECAP_INV_G11
XG11018 XI11_2/XI0/XI0_51/d_12_ XI11_2/XI0/XI0_51/d__12_ DECAP_INV_G11
XG11019 XI11_2/XI0/XI0_51/d_11_ XI11_2/XI0/XI0_51/d__11_ DECAP_INV_G11
XG11020 XI11_2/XI0/XI0_51/d_10_ XI11_2/XI0/XI0_51/d__10_ DECAP_INV_G11
XG11021 XI11_2/XI0/XI0_51/d_9_ XI11_2/XI0/XI0_51/d__9_ DECAP_INV_G11
XG11022 XI11_2/XI0/XI0_51/d_8_ XI11_2/XI0/XI0_51/d__8_ DECAP_INV_G11
XG11023 XI11_2/XI0/XI0_51/d_7_ XI11_2/XI0/XI0_51/d__7_ DECAP_INV_G11
XG11024 XI11_2/XI0/XI0_51/d_6_ XI11_2/XI0/XI0_51/d__6_ DECAP_INV_G11
XG11025 XI11_2/XI0/XI0_51/d_5_ XI11_2/XI0/XI0_51/d__5_ DECAP_INV_G11
XG11026 XI11_2/XI0/XI0_51/d_4_ XI11_2/XI0/XI0_51/d__4_ DECAP_INV_G11
XG11027 XI11_2/XI0/XI0_51/d_3_ XI11_2/XI0/XI0_51/d__3_ DECAP_INV_G11
XG11028 XI11_2/XI0/XI0_51/d_2_ XI11_2/XI0/XI0_51/d__2_ DECAP_INV_G11
XG11029 XI11_2/XI0/XI0_51/d_1_ XI11_2/XI0/XI0_51/d__1_ DECAP_INV_G11
XG11030 XI11_2/XI0/XI0_51/d_0_ XI11_2/XI0/XI0_51/d__0_ DECAP_INV_G11
XG11031 XI11_2/XI0/XI0_50/d__15_ XI11_2/XI0/XI0_50/d_15_ DECAP_INV_G11
XG11032 XI11_2/XI0/XI0_50/d__14_ XI11_2/XI0/XI0_50/d_14_ DECAP_INV_G11
XG11033 XI11_2/XI0/XI0_50/d__13_ XI11_2/XI0/XI0_50/d_13_ DECAP_INV_G11
XG11034 XI11_2/XI0/XI0_50/d__12_ XI11_2/XI0/XI0_50/d_12_ DECAP_INV_G11
XG11035 XI11_2/XI0/XI0_50/d__11_ XI11_2/XI0/XI0_50/d_11_ DECAP_INV_G11
XG11036 XI11_2/XI0/XI0_50/d__10_ XI11_2/XI0/XI0_50/d_10_ DECAP_INV_G11
XG11037 XI11_2/XI0/XI0_50/d__9_ XI11_2/XI0/XI0_50/d_9_ DECAP_INV_G11
XG11038 XI11_2/XI0/XI0_50/d__8_ XI11_2/XI0/XI0_50/d_8_ DECAP_INV_G11
XG11039 XI11_2/XI0/XI0_50/d__7_ XI11_2/XI0/XI0_50/d_7_ DECAP_INV_G11
XG11040 XI11_2/XI0/XI0_50/d__6_ XI11_2/XI0/XI0_50/d_6_ DECAP_INV_G11
XG11041 XI11_2/XI0/XI0_50/d__5_ XI11_2/XI0/XI0_50/d_5_ DECAP_INV_G11
XG11042 XI11_2/XI0/XI0_50/d__4_ XI11_2/XI0/XI0_50/d_4_ DECAP_INV_G11
XG11043 XI11_2/XI0/XI0_50/d__3_ XI11_2/XI0/XI0_50/d_3_ DECAP_INV_G11
XG11044 XI11_2/XI0/XI0_50/d__2_ XI11_2/XI0/XI0_50/d_2_ DECAP_INV_G11
XG11045 XI11_2/XI0/XI0_50/d__1_ XI11_2/XI0/XI0_50/d_1_ DECAP_INV_G11
XG11046 XI11_2/XI0/XI0_50/d__0_ XI11_2/XI0/XI0_50/d_0_ DECAP_INV_G11
XG11047 XI11_2/XI0/XI0_50/d_15_ XI11_2/XI0/XI0_50/d__15_ DECAP_INV_G11
XG11048 XI11_2/XI0/XI0_50/d_14_ XI11_2/XI0/XI0_50/d__14_ DECAP_INV_G11
XG11049 XI11_2/XI0/XI0_50/d_13_ XI11_2/XI0/XI0_50/d__13_ DECAP_INV_G11
XG11050 XI11_2/XI0/XI0_50/d_12_ XI11_2/XI0/XI0_50/d__12_ DECAP_INV_G11
XG11051 XI11_2/XI0/XI0_50/d_11_ XI11_2/XI0/XI0_50/d__11_ DECAP_INV_G11
XG11052 XI11_2/XI0/XI0_50/d_10_ XI11_2/XI0/XI0_50/d__10_ DECAP_INV_G11
XG11053 XI11_2/XI0/XI0_50/d_9_ XI11_2/XI0/XI0_50/d__9_ DECAP_INV_G11
XG11054 XI11_2/XI0/XI0_50/d_8_ XI11_2/XI0/XI0_50/d__8_ DECAP_INV_G11
XG11055 XI11_2/XI0/XI0_50/d_7_ XI11_2/XI0/XI0_50/d__7_ DECAP_INV_G11
XG11056 XI11_2/XI0/XI0_50/d_6_ XI11_2/XI0/XI0_50/d__6_ DECAP_INV_G11
XG11057 XI11_2/XI0/XI0_50/d_5_ XI11_2/XI0/XI0_50/d__5_ DECAP_INV_G11
XG11058 XI11_2/XI0/XI0_50/d_4_ XI11_2/XI0/XI0_50/d__4_ DECAP_INV_G11
XG11059 XI11_2/XI0/XI0_50/d_3_ XI11_2/XI0/XI0_50/d__3_ DECAP_INV_G11
XG11060 XI11_2/XI0/XI0_50/d_2_ XI11_2/XI0/XI0_50/d__2_ DECAP_INV_G11
XG11061 XI11_2/XI0/XI0_50/d_1_ XI11_2/XI0/XI0_50/d__1_ DECAP_INV_G11
XG11062 XI11_2/XI0/XI0_50/d_0_ XI11_2/XI0/XI0_50/d__0_ DECAP_INV_G11
XG11063 XI11_2/XI0/XI0_49/d__15_ XI11_2/XI0/XI0_49/d_15_ DECAP_INV_G11
XG11064 XI11_2/XI0/XI0_49/d__14_ XI11_2/XI0/XI0_49/d_14_ DECAP_INV_G11
XG11065 XI11_2/XI0/XI0_49/d__13_ XI11_2/XI0/XI0_49/d_13_ DECAP_INV_G11
XG11066 XI11_2/XI0/XI0_49/d__12_ XI11_2/XI0/XI0_49/d_12_ DECAP_INV_G11
XG11067 XI11_2/XI0/XI0_49/d__11_ XI11_2/XI0/XI0_49/d_11_ DECAP_INV_G11
XG11068 XI11_2/XI0/XI0_49/d__10_ XI11_2/XI0/XI0_49/d_10_ DECAP_INV_G11
XG11069 XI11_2/XI0/XI0_49/d__9_ XI11_2/XI0/XI0_49/d_9_ DECAP_INV_G11
XG11070 XI11_2/XI0/XI0_49/d__8_ XI11_2/XI0/XI0_49/d_8_ DECAP_INV_G11
XG11071 XI11_2/XI0/XI0_49/d__7_ XI11_2/XI0/XI0_49/d_7_ DECAP_INV_G11
XG11072 XI11_2/XI0/XI0_49/d__6_ XI11_2/XI0/XI0_49/d_6_ DECAP_INV_G11
XG11073 XI11_2/XI0/XI0_49/d__5_ XI11_2/XI0/XI0_49/d_5_ DECAP_INV_G11
XG11074 XI11_2/XI0/XI0_49/d__4_ XI11_2/XI0/XI0_49/d_4_ DECAP_INV_G11
XG11075 XI11_2/XI0/XI0_49/d__3_ XI11_2/XI0/XI0_49/d_3_ DECAP_INV_G11
XG11076 XI11_2/XI0/XI0_49/d__2_ XI11_2/XI0/XI0_49/d_2_ DECAP_INV_G11
XG11077 XI11_2/XI0/XI0_49/d__1_ XI11_2/XI0/XI0_49/d_1_ DECAP_INV_G11
XG11078 XI11_2/XI0/XI0_49/d__0_ XI11_2/XI0/XI0_49/d_0_ DECAP_INV_G11
XG11079 XI11_2/XI0/XI0_49/d_15_ XI11_2/XI0/XI0_49/d__15_ DECAP_INV_G11
XG11080 XI11_2/XI0/XI0_49/d_14_ XI11_2/XI0/XI0_49/d__14_ DECAP_INV_G11
XG11081 XI11_2/XI0/XI0_49/d_13_ XI11_2/XI0/XI0_49/d__13_ DECAP_INV_G11
XG11082 XI11_2/XI0/XI0_49/d_12_ XI11_2/XI0/XI0_49/d__12_ DECAP_INV_G11
XG11083 XI11_2/XI0/XI0_49/d_11_ XI11_2/XI0/XI0_49/d__11_ DECAP_INV_G11
XG11084 XI11_2/XI0/XI0_49/d_10_ XI11_2/XI0/XI0_49/d__10_ DECAP_INV_G11
XG11085 XI11_2/XI0/XI0_49/d_9_ XI11_2/XI0/XI0_49/d__9_ DECAP_INV_G11
XG11086 XI11_2/XI0/XI0_49/d_8_ XI11_2/XI0/XI0_49/d__8_ DECAP_INV_G11
XG11087 XI11_2/XI0/XI0_49/d_7_ XI11_2/XI0/XI0_49/d__7_ DECAP_INV_G11
XG11088 XI11_2/XI0/XI0_49/d_6_ XI11_2/XI0/XI0_49/d__6_ DECAP_INV_G11
XG11089 XI11_2/XI0/XI0_49/d_5_ XI11_2/XI0/XI0_49/d__5_ DECAP_INV_G11
XG11090 XI11_2/XI0/XI0_49/d_4_ XI11_2/XI0/XI0_49/d__4_ DECAP_INV_G11
XG11091 XI11_2/XI0/XI0_49/d_3_ XI11_2/XI0/XI0_49/d__3_ DECAP_INV_G11
XG11092 XI11_2/XI0/XI0_49/d_2_ XI11_2/XI0/XI0_49/d__2_ DECAP_INV_G11
XG11093 XI11_2/XI0/XI0_49/d_1_ XI11_2/XI0/XI0_49/d__1_ DECAP_INV_G11
XG11094 XI11_2/XI0/XI0_49/d_0_ XI11_2/XI0/XI0_49/d__0_ DECAP_INV_G11
XG11095 XI11_2/XI0/XI0_48/d__15_ XI11_2/XI0/XI0_48/d_15_ DECAP_INV_G11
XG11096 XI11_2/XI0/XI0_48/d__14_ XI11_2/XI0/XI0_48/d_14_ DECAP_INV_G11
XG11097 XI11_2/XI0/XI0_48/d__13_ XI11_2/XI0/XI0_48/d_13_ DECAP_INV_G11
XG11098 XI11_2/XI0/XI0_48/d__12_ XI11_2/XI0/XI0_48/d_12_ DECAP_INV_G11
XG11099 XI11_2/XI0/XI0_48/d__11_ XI11_2/XI0/XI0_48/d_11_ DECAP_INV_G11
XG11100 XI11_2/XI0/XI0_48/d__10_ XI11_2/XI0/XI0_48/d_10_ DECAP_INV_G11
XG11101 XI11_2/XI0/XI0_48/d__9_ XI11_2/XI0/XI0_48/d_9_ DECAP_INV_G11
XG11102 XI11_2/XI0/XI0_48/d__8_ XI11_2/XI0/XI0_48/d_8_ DECAP_INV_G11
XG11103 XI11_2/XI0/XI0_48/d__7_ XI11_2/XI0/XI0_48/d_7_ DECAP_INV_G11
XG11104 XI11_2/XI0/XI0_48/d__6_ XI11_2/XI0/XI0_48/d_6_ DECAP_INV_G11
XG11105 XI11_2/XI0/XI0_48/d__5_ XI11_2/XI0/XI0_48/d_5_ DECAP_INV_G11
XG11106 XI11_2/XI0/XI0_48/d__4_ XI11_2/XI0/XI0_48/d_4_ DECAP_INV_G11
XG11107 XI11_2/XI0/XI0_48/d__3_ XI11_2/XI0/XI0_48/d_3_ DECAP_INV_G11
XG11108 XI11_2/XI0/XI0_48/d__2_ XI11_2/XI0/XI0_48/d_2_ DECAP_INV_G11
XG11109 XI11_2/XI0/XI0_48/d__1_ XI11_2/XI0/XI0_48/d_1_ DECAP_INV_G11
XG11110 XI11_2/XI0/XI0_48/d__0_ XI11_2/XI0/XI0_48/d_0_ DECAP_INV_G11
XG11111 XI11_2/XI0/XI0_48/d_15_ XI11_2/XI0/XI0_48/d__15_ DECAP_INV_G11
XG11112 XI11_2/XI0/XI0_48/d_14_ XI11_2/XI0/XI0_48/d__14_ DECAP_INV_G11
XG11113 XI11_2/XI0/XI0_48/d_13_ XI11_2/XI0/XI0_48/d__13_ DECAP_INV_G11
XG11114 XI11_2/XI0/XI0_48/d_12_ XI11_2/XI0/XI0_48/d__12_ DECAP_INV_G11
XG11115 XI11_2/XI0/XI0_48/d_11_ XI11_2/XI0/XI0_48/d__11_ DECAP_INV_G11
XG11116 XI11_2/XI0/XI0_48/d_10_ XI11_2/XI0/XI0_48/d__10_ DECAP_INV_G11
XG11117 XI11_2/XI0/XI0_48/d_9_ XI11_2/XI0/XI0_48/d__9_ DECAP_INV_G11
XG11118 XI11_2/XI0/XI0_48/d_8_ XI11_2/XI0/XI0_48/d__8_ DECAP_INV_G11
XG11119 XI11_2/XI0/XI0_48/d_7_ XI11_2/XI0/XI0_48/d__7_ DECAP_INV_G11
XG11120 XI11_2/XI0/XI0_48/d_6_ XI11_2/XI0/XI0_48/d__6_ DECAP_INV_G11
XG11121 XI11_2/XI0/XI0_48/d_5_ XI11_2/XI0/XI0_48/d__5_ DECAP_INV_G11
XG11122 XI11_2/XI0/XI0_48/d_4_ XI11_2/XI0/XI0_48/d__4_ DECAP_INV_G11
XG11123 XI11_2/XI0/XI0_48/d_3_ XI11_2/XI0/XI0_48/d__3_ DECAP_INV_G11
XG11124 XI11_2/XI0/XI0_48/d_2_ XI11_2/XI0/XI0_48/d__2_ DECAP_INV_G11
XG11125 XI11_2/XI0/XI0_48/d_1_ XI11_2/XI0/XI0_48/d__1_ DECAP_INV_G11
XG11126 XI11_2/XI0/XI0_48/d_0_ XI11_2/XI0/XI0_48/d__0_ DECAP_INV_G11
XG11127 XI11_2/XI0/XI0_47/d__15_ XI11_2/XI0/XI0_47/d_15_ DECAP_INV_G11
XG11128 XI11_2/XI0/XI0_47/d__14_ XI11_2/XI0/XI0_47/d_14_ DECAP_INV_G11
XG11129 XI11_2/XI0/XI0_47/d__13_ XI11_2/XI0/XI0_47/d_13_ DECAP_INV_G11
XG11130 XI11_2/XI0/XI0_47/d__12_ XI11_2/XI0/XI0_47/d_12_ DECAP_INV_G11
XG11131 XI11_2/XI0/XI0_47/d__11_ XI11_2/XI0/XI0_47/d_11_ DECAP_INV_G11
XG11132 XI11_2/XI0/XI0_47/d__10_ XI11_2/XI0/XI0_47/d_10_ DECAP_INV_G11
XG11133 XI11_2/XI0/XI0_47/d__9_ XI11_2/XI0/XI0_47/d_9_ DECAP_INV_G11
XG11134 XI11_2/XI0/XI0_47/d__8_ XI11_2/XI0/XI0_47/d_8_ DECAP_INV_G11
XG11135 XI11_2/XI0/XI0_47/d__7_ XI11_2/XI0/XI0_47/d_7_ DECAP_INV_G11
XG11136 XI11_2/XI0/XI0_47/d__6_ XI11_2/XI0/XI0_47/d_6_ DECAP_INV_G11
XG11137 XI11_2/XI0/XI0_47/d__5_ XI11_2/XI0/XI0_47/d_5_ DECAP_INV_G11
XG11138 XI11_2/XI0/XI0_47/d__4_ XI11_2/XI0/XI0_47/d_4_ DECAP_INV_G11
XG11139 XI11_2/XI0/XI0_47/d__3_ XI11_2/XI0/XI0_47/d_3_ DECAP_INV_G11
XG11140 XI11_2/XI0/XI0_47/d__2_ XI11_2/XI0/XI0_47/d_2_ DECAP_INV_G11
XG11141 XI11_2/XI0/XI0_47/d__1_ XI11_2/XI0/XI0_47/d_1_ DECAP_INV_G11
XG11142 XI11_2/XI0/XI0_47/d__0_ XI11_2/XI0/XI0_47/d_0_ DECAP_INV_G11
XG11143 XI11_2/XI0/XI0_47/d_15_ XI11_2/XI0/XI0_47/d__15_ DECAP_INV_G11
XG11144 XI11_2/XI0/XI0_47/d_14_ XI11_2/XI0/XI0_47/d__14_ DECAP_INV_G11
XG11145 XI11_2/XI0/XI0_47/d_13_ XI11_2/XI0/XI0_47/d__13_ DECAP_INV_G11
XG11146 XI11_2/XI0/XI0_47/d_12_ XI11_2/XI0/XI0_47/d__12_ DECAP_INV_G11
XG11147 XI11_2/XI0/XI0_47/d_11_ XI11_2/XI0/XI0_47/d__11_ DECAP_INV_G11
XG11148 XI11_2/XI0/XI0_47/d_10_ XI11_2/XI0/XI0_47/d__10_ DECAP_INV_G11
XG11149 XI11_2/XI0/XI0_47/d_9_ XI11_2/XI0/XI0_47/d__9_ DECAP_INV_G11
XG11150 XI11_2/XI0/XI0_47/d_8_ XI11_2/XI0/XI0_47/d__8_ DECAP_INV_G11
XG11151 XI11_2/XI0/XI0_47/d_7_ XI11_2/XI0/XI0_47/d__7_ DECAP_INV_G11
XG11152 XI11_2/XI0/XI0_47/d_6_ XI11_2/XI0/XI0_47/d__6_ DECAP_INV_G11
XG11153 XI11_2/XI0/XI0_47/d_5_ XI11_2/XI0/XI0_47/d__5_ DECAP_INV_G11
XG11154 XI11_2/XI0/XI0_47/d_4_ XI11_2/XI0/XI0_47/d__4_ DECAP_INV_G11
XG11155 XI11_2/XI0/XI0_47/d_3_ XI11_2/XI0/XI0_47/d__3_ DECAP_INV_G11
XG11156 XI11_2/XI0/XI0_47/d_2_ XI11_2/XI0/XI0_47/d__2_ DECAP_INV_G11
XG11157 XI11_2/XI0/XI0_47/d_1_ XI11_2/XI0/XI0_47/d__1_ DECAP_INV_G11
XG11158 XI11_2/XI0/XI0_47/d_0_ XI11_2/XI0/XI0_47/d__0_ DECAP_INV_G11
XG11159 XI11_2/XI0/XI0_46/d__15_ XI11_2/XI0/XI0_46/d_15_ DECAP_INV_G11
XG11160 XI11_2/XI0/XI0_46/d__14_ XI11_2/XI0/XI0_46/d_14_ DECAP_INV_G11
XG11161 XI11_2/XI0/XI0_46/d__13_ XI11_2/XI0/XI0_46/d_13_ DECAP_INV_G11
XG11162 XI11_2/XI0/XI0_46/d__12_ XI11_2/XI0/XI0_46/d_12_ DECAP_INV_G11
XG11163 XI11_2/XI0/XI0_46/d__11_ XI11_2/XI0/XI0_46/d_11_ DECAP_INV_G11
XG11164 XI11_2/XI0/XI0_46/d__10_ XI11_2/XI0/XI0_46/d_10_ DECAP_INV_G11
XG11165 XI11_2/XI0/XI0_46/d__9_ XI11_2/XI0/XI0_46/d_9_ DECAP_INV_G11
XG11166 XI11_2/XI0/XI0_46/d__8_ XI11_2/XI0/XI0_46/d_8_ DECAP_INV_G11
XG11167 XI11_2/XI0/XI0_46/d__7_ XI11_2/XI0/XI0_46/d_7_ DECAP_INV_G11
XG11168 XI11_2/XI0/XI0_46/d__6_ XI11_2/XI0/XI0_46/d_6_ DECAP_INV_G11
XG11169 XI11_2/XI0/XI0_46/d__5_ XI11_2/XI0/XI0_46/d_5_ DECAP_INV_G11
XG11170 XI11_2/XI0/XI0_46/d__4_ XI11_2/XI0/XI0_46/d_4_ DECAP_INV_G11
XG11171 XI11_2/XI0/XI0_46/d__3_ XI11_2/XI0/XI0_46/d_3_ DECAP_INV_G11
XG11172 XI11_2/XI0/XI0_46/d__2_ XI11_2/XI0/XI0_46/d_2_ DECAP_INV_G11
XG11173 XI11_2/XI0/XI0_46/d__1_ XI11_2/XI0/XI0_46/d_1_ DECAP_INV_G11
XG11174 XI11_2/XI0/XI0_46/d__0_ XI11_2/XI0/XI0_46/d_0_ DECAP_INV_G11
XG11175 XI11_2/XI0/XI0_46/d_15_ XI11_2/XI0/XI0_46/d__15_ DECAP_INV_G11
XG11176 XI11_2/XI0/XI0_46/d_14_ XI11_2/XI0/XI0_46/d__14_ DECAP_INV_G11
XG11177 XI11_2/XI0/XI0_46/d_13_ XI11_2/XI0/XI0_46/d__13_ DECAP_INV_G11
XG11178 XI11_2/XI0/XI0_46/d_12_ XI11_2/XI0/XI0_46/d__12_ DECAP_INV_G11
XG11179 XI11_2/XI0/XI0_46/d_11_ XI11_2/XI0/XI0_46/d__11_ DECAP_INV_G11
XG11180 XI11_2/XI0/XI0_46/d_10_ XI11_2/XI0/XI0_46/d__10_ DECAP_INV_G11
XG11181 XI11_2/XI0/XI0_46/d_9_ XI11_2/XI0/XI0_46/d__9_ DECAP_INV_G11
XG11182 XI11_2/XI0/XI0_46/d_8_ XI11_2/XI0/XI0_46/d__8_ DECAP_INV_G11
XG11183 XI11_2/XI0/XI0_46/d_7_ XI11_2/XI0/XI0_46/d__7_ DECAP_INV_G11
XG11184 XI11_2/XI0/XI0_46/d_6_ XI11_2/XI0/XI0_46/d__6_ DECAP_INV_G11
XG11185 XI11_2/XI0/XI0_46/d_5_ XI11_2/XI0/XI0_46/d__5_ DECAP_INV_G11
XG11186 XI11_2/XI0/XI0_46/d_4_ XI11_2/XI0/XI0_46/d__4_ DECAP_INV_G11
XG11187 XI11_2/XI0/XI0_46/d_3_ XI11_2/XI0/XI0_46/d__3_ DECAP_INV_G11
XG11188 XI11_2/XI0/XI0_46/d_2_ XI11_2/XI0/XI0_46/d__2_ DECAP_INV_G11
XG11189 XI11_2/XI0/XI0_46/d_1_ XI11_2/XI0/XI0_46/d__1_ DECAP_INV_G11
XG11190 XI11_2/XI0/XI0_46/d_0_ XI11_2/XI0/XI0_46/d__0_ DECAP_INV_G11
XG11191 XI11_2/XI0/XI0_45/d__15_ XI11_2/XI0/XI0_45/d_15_ DECAP_INV_G11
XG11192 XI11_2/XI0/XI0_45/d__14_ XI11_2/XI0/XI0_45/d_14_ DECAP_INV_G11
XG11193 XI11_2/XI0/XI0_45/d__13_ XI11_2/XI0/XI0_45/d_13_ DECAP_INV_G11
XG11194 XI11_2/XI0/XI0_45/d__12_ XI11_2/XI0/XI0_45/d_12_ DECAP_INV_G11
XG11195 XI11_2/XI0/XI0_45/d__11_ XI11_2/XI0/XI0_45/d_11_ DECAP_INV_G11
XG11196 XI11_2/XI0/XI0_45/d__10_ XI11_2/XI0/XI0_45/d_10_ DECAP_INV_G11
XG11197 XI11_2/XI0/XI0_45/d__9_ XI11_2/XI0/XI0_45/d_9_ DECAP_INV_G11
XG11198 XI11_2/XI0/XI0_45/d__8_ XI11_2/XI0/XI0_45/d_8_ DECAP_INV_G11
XG11199 XI11_2/XI0/XI0_45/d__7_ XI11_2/XI0/XI0_45/d_7_ DECAP_INV_G11
XG11200 XI11_2/XI0/XI0_45/d__6_ XI11_2/XI0/XI0_45/d_6_ DECAP_INV_G11
XG11201 XI11_2/XI0/XI0_45/d__5_ XI11_2/XI0/XI0_45/d_5_ DECAP_INV_G11
XG11202 XI11_2/XI0/XI0_45/d__4_ XI11_2/XI0/XI0_45/d_4_ DECAP_INV_G11
XG11203 XI11_2/XI0/XI0_45/d__3_ XI11_2/XI0/XI0_45/d_3_ DECAP_INV_G11
XG11204 XI11_2/XI0/XI0_45/d__2_ XI11_2/XI0/XI0_45/d_2_ DECAP_INV_G11
XG11205 XI11_2/XI0/XI0_45/d__1_ XI11_2/XI0/XI0_45/d_1_ DECAP_INV_G11
XG11206 XI11_2/XI0/XI0_45/d__0_ XI11_2/XI0/XI0_45/d_0_ DECAP_INV_G11
XG11207 XI11_2/XI0/XI0_45/d_15_ XI11_2/XI0/XI0_45/d__15_ DECAP_INV_G11
XG11208 XI11_2/XI0/XI0_45/d_14_ XI11_2/XI0/XI0_45/d__14_ DECAP_INV_G11
XG11209 XI11_2/XI0/XI0_45/d_13_ XI11_2/XI0/XI0_45/d__13_ DECAP_INV_G11
XG11210 XI11_2/XI0/XI0_45/d_12_ XI11_2/XI0/XI0_45/d__12_ DECAP_INV_G11
XG11211 XI11_2/XI0/XI0_45/d_11_ XI11_2/XI0/XI0_45/d__11_ DECAP_INV_G11
XG11212 XI11_2/XI0/XI0_45/d_10_ XI11_2/XI0/XI0_45/d__10_ DECAP_INV_G11
XG11213 XI11_2/XI0/XI0_45/d_9_ XI11_2/XI0/XI0_45/d__9_ DECAP_INV_G11
XG11214 XI11_2/XI0/XI0_45/d_8_ XI11_2/XI0/XI0_45/d__8_ DECAP_INV_G11
XG11215 XI11_2/XI0/XI0_45/d_7_ XI11_2/XI0/XI0_45/d__7_ DECAP_INV_G11
XG11216 XI11_2/XI0/XI0_45/d_6_ XI11_2/XI0/XI0_45/d__6_ DECAP_INV_G11
XG11217 XI11_2/XI0/XI0_45/d_5_ XI11_2/XI0/XI0_45/d__5_ DECAP_INV_G11
XG11218 XI11_2/XI0/XI0_45/d_4_ XI11_2/XI0/XI0_45/d__4_ DECAP_INV_G11
XG11219 XI11_2/XI0/XI0_45/d_3_ XI11_2/XI0/XI0_45/d__3_ DECAP_INV_G11
XG11220 XI11_2/XI0/XI0_45/d_2_ XI11_2/XI0/XI0_45/d__2_ DECAP_INV_G11
XG11221 XI11_2/XI0/XI0_45/d_1_ XI11_2/XI0/XI0_45/d__1_ DECAP_INV_G11
XG11222 XI11_2/XI0/XI0_45/d_0_ XI11_2/XI0/XI0_45/d__0_ DECAP_INV_G11
XG11223 XI11_2/XI0/XI0_44/d__15_ XI11_2/XI0/XI0_44/d_15_ DECAP_INV_G11
XG11224 XI11_2/XI0/XI0_44/d__14_ XI11_2/XI0/XI0_44/d_14_ DECAP_INV_G11
XG11225 XI11_2/XI0/XI0_44/d__13_ XI11_2/XI0/XI0_44/d_13_ DECAP_INV_G11
XG11226 XI11_2/XI0/XI0_44/d__12_ XI11_2/XI0/XI0_44/d_12_ DECAP_INV_G11
XG11227 XI11_2/XI0/XI0_44/d__11_ XI11_2/XI0/XI0_44/d_11_ DECAP_INV_G11
XG11228 XI11_2/XI0/XI0_44/d__10_ XI11_2/XI0/XI0_44/d_10_ DECAP_INV_G11
XG11229 XI11_2/XI0/XI0_44/d__9_ XI11_2/XI0/XI0_44/d_9_ DECAP_INV_G11
XG11230 XI11_2/XI0/XI0_44/d__8_ XI11_2/XI0/XI0_44/d_8_ DECAP_INV_G11
XG11231 XI11_2/XI0/XI0_44/d__7_ XI11_2/XI0/XI0_44/d_7_ DECAP_INV_G11
XG11232 XI11_2/XI0/XI0_44/d__6_ XI11_2/XI0/XI0_44/d_6_ DECAP_INV_G11
XG11233 XI11_2/XI0/XI0_44/d__5_ XI11_2/XI0/XI0_44/d_5_ DECAP_INV_G11
XG11234 XI11_2/XI0/XI0_44/d__4_ XI11_2/XI0/XI0_44/d_4_ DECAP_INV_G11
XG11235 XI11_2/XI0/XI0_44/d__3_ XI11_2/XI0/XI0_44/d_3_ DECAP_INV_G11
XG11236 XI11_2/XI0/XI0_44/d__2_ XI11_2/XI0/XI0_44/d_2_ DECAP_INV_G11
XG11237 XI11_2/XI0/XI0_44/d__1_ XI11_2/XI0/XI0_44/d_1_ DECAP_INV_G11
XG11238 XI11_2/XI0/XI0_44/d__0_ XI11_2/XI0/XI0_44/d_0_ DECAP_INV_G11
XG11239 XI11_2/XI0/XI0_44/d_15_ XI11_2/XI0/XI0_44/d__15_ DECAP_INV_G11
XG11240 XI11_2/XI0/XI0_44/d_14_ XI11_2/XI0/XI0_44/d__14_ DECAP_INV_G11
XG11241 XI11_2/XI0/XI0_44/d_13_ XI11_2/XI0/XI0_44/d__13_ DECAP_INV_G11
XG11242 XI11_2/XI0/XI0_44/d_12_ XI11_2/XI0/XI0_44/d__12_ DECAP_INV_G11
XG11243 XI11_2/XI0/XI0_44/d_11_ XI11_2/XI0/XI0_44/d__11_ DECAP_INV_G11
XG11244 XI11_2/XI0/XI0_44/d_10_ XI11_2/XI0/XI0_44/d__10_ DECAP_INV_G11
XG11245 XI11_2/XI0/XI0_44/d_9_ XI11_2/XI0/XI0_44/d__9_ DECAP_INV_G11
XG11246 XI11_2/XI0/XI0_44/d_8_ XI11_2/XI0/XI0_44/d__8_ DECAP_INV_G11
XG11247 XI11_2/XI0/XI0_44/d_7_ XI11_2/XI0/XI0_44/d__7_ DECAP_INV_G11
XG11248 XI11_2/XI0/XI0_44/d_6_ XI11_2/XI0/XI0_44/d__6_ DECAP_INV_G11
XG11249 XI11_2/XI0/XI0_44/d_5_ XI11_2/XI0/XI0_44/d__5_ DECAP_INV_G11
XG11250 XI11_2/XI0/XI0_44/d_4_ XI11_2/XI0/XI0_44/d__4_ DECAP_INV_G11
XG11251 XI11_2/XI0/XI0_44/d_3_ XI11_2/XI0/XI0_44/d__3_ DECAP_INV_G11
XG11252 XI11_2/XI0/XI0_44/d_2_ XI11_2/XI0/XI0_44/d__2_ DECAP_INV_G11
XG11253 XI11_2/XI0/XI0_44/d_1_ XI11_2/XI0/XI0_44/d__1_ DECAP_INV_G11
XG11254 XI11_2/XI0/XI0_44/d_0_ XI11_2/XI0/XI0_44/d__0_ DECAP_INV_G11
XG11255 XI11_2/XI0/XI0_43/d__15_ XI11_2/XI0/XI0_43/d_15_ DECAP_INV_G11
XG11256 XI11_2/XI0/XI0_43/d__14_ XI11_2/XI0/XI0_43/d_14_ DECAP_INV_G11
XG11257 XI11_2/XI0/XI0_43/d__13_ XI11_2/XI0/XI0_43/d_13_ DECAP_INV_G11
XG11258 XI11_2/XI0/XI0_43/d__12_ XI11_2/XI0/XI0_43/d_12_ DECAP_INV_G11
XG11259 XI11_2/XI0/XI0_43/d__11_ XI11_2/XI0/XI0_43/d_11_ DECAP_INV_G11
XG11260 XI11_2/XI0/XI0_43/d__10_ XI11_2/XI0/XI0_43/d_10_ DECAP_INV_G11
XG11261 XI11_2/XI0/XI0_43/d__9_ XI11_2/XI0/XI0_43/d_9_ DECAP_INV_G11
XG11262 XI11_2/XI0/XI0_43/d__8_ XI11_2/XI0/XI0_43/d_8_ DECAP_INV_G11
XG11263 XI11_2/XI0/XI0_43/d__7_ XI11_2/XI0/XI0_43/d_7_ DECAP_INV_G11
XG11264 XI11_2/XI0/XI0_43/d__6_ XI11_2/XI0/XI0_43/d_6_ DECAP_INV_G11
XG11265 XI11_2/XI0/XI0_43/d__5_ XI11_2/XI0/XI0_43/d_5_ DECAP_INV_G11
XG11266 XI11_2/XI0/XI0_43/d__4_ XI11_2/XI0/XI0_43/d_4_ DECAP_INV_G11
XG11267 XI11_2/XI0/XI0_43/d__3_ XI11_2/XI0/XI0_43/d_3_ DECAP_INV_G11
XG11268 XI11_2/XI0/XI0_43/d__2_ XI11_2/XI0/XI0_43/d_2_ DECAP_INV_G11
XG11269 XI11_2/XI0/XI0_43/d__1_ XI11_2/XI0/XI0_43/d_1_ DECAP_INV_G11
XG11270 XI11_2/XI0/XI0_43/d__0_ XI11_2/XI0/XI0_43/d_0_ DECAP_INV_G11
XG11271 XI11_2/XI0/XI0_43/d_15_ XI11_2/XI0/XI0_43/d__15_ DECAP_INV_G11
XG11272 XI11_2/XI0/XI0_43/d_14_ XI11_2/XI0/XI0_43/d__14_ DECAP_INV_G11
XG11273 XI11_2/XI0/XI0_43/d_13_ XI11_2/XI0/XI0_43/d__13_ DECAP_INV_G11
XG11274 XI11_2/XI0/XI0_43/d_12_ XI11_2/XI0/XI0_43/d__12_ DECAP_INV_G11
XG11275 XI11_2/XI0/XI0_43/d_11_ XI11_2/XI0/XI0_43/d__11_ DECAP_INV_G11
XG11276 XI11_2/XI0/XI0_43/d_10_ XI11_2/XI0/XI0_43/d__10_ DECAP_INV_G11
XG11277 XI11_2/XI0/XI0_43/d_9_ XI11_2/XI0/XI0_43/d__9_ DECAP_INV_G11
XG11278 XI11_2/XI0/XI0_43/d_8_ XI11_2/XI0/XI0_43/d__8_ DECAP_INV_G11
XG11279 XI11_2/XI0/XI0_43/d_7_ XI11_2/XI0/XI0_43/d__7_ DECAP_INV_G11
XG11280 XI11_2/XI0/XI0_43/d_6_ XI11_2/XI0/XI0_43/d__6_ DECAP_INV_G11
XG11281 XI11_2/XI0/XI0_43/d_5_ XI11_2/XI0/XI0_43/d__5_ DECAP_INV_G11
XG11282 XI11_2/XI0/XI0_43/d_4_ XI11_2/XI0/XI0_43/d__4_ DECAP_INV_G11
XG11283 XI11_2/XI0/XI0_43/d_3_ XI11_2/XI0/XI0_43/d__3_ DECAP_INV_G11
XG11284 XI11_2/XI0/XI0_43/d_2_ XI11_2/XI0/XI0_43/d__2_ DECAP_INV_G11
XG11285 XI11_2/XI0/XI0_43/d_1_ XI11_2/XI0/XI0_43/d__1_ DECAP_INV_G11
XG11286 XI11_2/XI0/XI0_43/d_0_ XI11_2/XI0/XI0_43/d__0_ DECAP_INV_G11
XG11287 XI11_2/XI0/XI0_42/d__15_ XI11_2/XI0/XI0_42/d_15_ DECAP_INV_G11
XG11288 XI11_2/XI0/XI0_42/d__14_ XI11_2/XI0/XI0_42/d_14_ DECAP_INV_G11
XG11289 XI11_2/XI0/XI0_42/d__13_ XI11_2/XI0/XI0_42/d_13_ DECAP_INV_G11
XG11290 XI11_2/XI0/XI0_42/d__12_ XI11_2/XI0/XI0_42/d_12_ DECAP_INV_G11
XG11291 XI11_2/XI0/XI0_42/d__11_ XI11_2/XI0/XI0_42/d_11_ DECAP_INV_G11
XG11292 XI11_2/XI0/XI0_42/d__10_ XI11_2/XI0/XI0_42/d_10_ DECAP_INV_G11
XG11293 XI11_2/XI0/XI0_42/d__9_ XI11_2/XI0/XI0_42/d_9_ DECAP_INV_G11
XG11294 XI11_2/XI0/XI0_42/d__8_ XI11_2/XI0/XI0_42/d_8_ DECAP_INV_G11
XG11295 XI11_2/XI0/XI0_42/d__7_ XI11_2/XI0/XI0_42/d_7_ DECAP_INV_G11
XG11296 XI11_2/XI0/XI0_42/d__6_ XI11_2/XI0/XI0_42/d_6_ DECAP_INV_G11
XG11297 XI11_2/XI0/XI0_42/d__5_ XI11_2/XI0/XI0_42/d_5_ DECAP_INV_G11
XG11298 XI11_2/XI0/XI0_42/d__4_ XI11_2/XI0/XI0_42/d_4_ DECAP_INV_G11
XG11299 XI11_2/XI0/XI0_42/d__3_ XI11_2/XI0/XI0_42/d_3_ DECAP_INV_G11
XG11300 XI11_2/XI0/XI0_42/d__2_ XI11_2/XI0/XI0_42/d_2_ DECAP_INV_G11
XG11301 XI11_2/XI0/XI0_42/d__1_ XI11_2/XI0/XI0_42/d_1_ DECAP_INV_G11
XG11302 XI11_2/XI0/XI0_42/d__0_ XI11_2/XI0/XI0_42/d_0_ DECAP_INV_G11
XG11303 XI11_2/XI0/XI0_42/d_15_ XI11_2/XI0/XI0_42/d__15_ DECAP_INV_G11
XG11304 XI11_2/XI0/XI0_42/d_14_ XI11_2/XI0/XI0_42/d__14_ DECAP_INV_G11
XG11305 XI11_2/XI0/XI0_42/d_13_ XI11_2/XI0/XI0_42/d__13_ DECAP_INV_G11
XG11306 XI11_2/XI0/XI0_42/d_12_ XI11_2/XI0/XI0_42/d__12_ DECAP_INV_G11
XG11307 XI11_2/XI0/XI0_42/d_11_ XI11_2/XI0/XI0_42/d__11_ DECAP_INV_G11
XG11308 XI11_2/XI0/XI0_42/d_10_ XI11_2/XI0/XI0_42/d__10_ DECAP_INV_G11
XG11309 XI11_2/XI0/XI0_42/d_9_ XI11_2/XI0/XI0_42/d__9_ DECAP_INV_G11
XG11310 XI11_2/XI0/XI0_42/d_8_ XI11_2/XI0/XI0_42/d__8_ DECAP_INV_G11
XG11311 XI11_2/XI0/XI0_42/d_7_ XI11_2/XI0/XI0_42/d__7_ DECAP_INV_G11
XG11312 XI11_2/XI0/XI0_42/d_6_ XI11_2/XI0/XI0_42/d__6_ DECAP_INV_G11
XG11313 XI11_2/XI0/XI0_42/d_5_ XI11_2/XI0/XI0_42/d__5_ DECAP_INV_G11
XG11314 XI11_2/XI0/XI0_42/d_4_ XI11_2/XI0/XI0_42/d__4_ DECAP_INV_G11
XG11315 XI11_2/XI0/XI0_42/d_3_ XI11_2/XI0/XI0_42/d__3_ DECAP_INV_G11
XG11316 XI11_2/XI0/XI0_42/d_2_ XI11_2/XI0/XI0_42/d__2_ DECAP_INV_G11
XG11317 XI11_2/XI0/XI0_42/d_1_ XI11_2/XI0/XI0_42/d__1_ DECAP_INV_G11
XG11318 XI11_2/XI0/XI0_42/d_0_ XI11_2/XI0/XI0_42/d__0_ DECAP_INV_G11
XG11319 XI11_2/XI0/XI0_41/d__15_ XI11_2/XI0/XI0_41/d_15_ DECAP_INV_G11
XG11320 XI11_2/XI0/XI0_41/d__14_ XI11_2/XI0/XI0_41/d_14_ DECAP_INV_G11
XG11321 XI11_2/XI0/XI0_41/d__13_ XI11_2/XI0/XI0_41/d_13_ DECAP_INV_G11
XG11322 XI11_2/XI0/XI0_41/d__12_ XI11_2/XI0/XI0_41/d_12_ DECAP_INV_G11
XG11323 XI11_2/XI0/XI0_41/d__11_ XI11_2/XI0/XI0_41/d_11_ DECAP_INV_G11
XG11324 XI11_2/XI0/XI0_41/d__10_ XI11_2/XI0/XI0_41/d_10_ DECAP_INV_G11
XG11325 XI11_2/XI0/XI0_41/d__9_ XI11_2/XI0/XI0_41/d_9_ DECAP_INV_G11
XG11326 XI11_2/XI0/XI0_41/d__8_ XI11_2/XI0/XI0_41/d_8_ DECAP_INV_G11
XG11327 XI11_2/XI0/XI0_41/d__7_ XI11_2/XI0/XI0_41/d_7_ DECAP_INV_G11
XG11328 XI11_2/XI0/XI0_41/d__6_ XI11_2/XI0/XI0_41/d_6_ DECAP_INV_G11
XG11329 XI11_2/XI0/XI0_41/d__5_ XI11_2/XI0/XI0_41/d_5_ DECAP_INV_G11
XG11330 XI11_2/XI0/XI0_41/d__4_ XI11_2/XI0/XI0_41/d_4_ DECAP_INV_G11
XG11331 XI11_2/XI0/XI0_41/d__3_ XI11_2/XI0/XI0_41/d_3_ DECAP_INV_G11
XG11332 XI11_2/XI0/XI0_41/d__2_ XI11_2/XI0/XI0_41/d_2_ DECAP_INV_G11
XG11333 XI11_2/XI0/XI0_41/d__1_ XI11_2/XI0/XI0_41/d_1_ DECAP_INV_G11
XG11334 XI11_2/XI0/XI0_41/d__0_ XI11_2/XI0/XI0_41/d_0_ DECAP_INV_G11
XG11335 XI11_2/XI0/XI0_41/d_15_ XI11_2/XI0/XI0_41/d__15_ DECAP_INV_G11
XG11336 XI11_2/XI0/XI0_41/d_14_ XI11_2/XI0/XI0_41/d__14_ DECAP_INV_G11
XG11337 XI11_2/XI0/XI0_41/d_13_ XI11_2/XI0/XI0_41/d__13_ DECAP_INV_G11
XG11338 XI11_2/XI0/XI0_41/d_12_ XI11_2/XI0/XI0_41/d__12_ DECAP_INV_G11
XG11339 XI11_2/XI0/XI0_41/d_11_ XI11_2/XI0/XI0_41/d__11_ DECAP_INV_G11
XG11340 XI11_2/XI0/XI0_41/d_10_ XI11_2/XI0/XI0_41/d__10_ DECAP_INV_G11
XG11341 XI11_2/XI0/XI0_41/d_9_ XI11_2/XI0/XI0_41/d__9_ DECAP_INV_G11
XG11342 XI11_2/XI0/XI0_41/d_8_ XI11_2/XI0/XI0_41/d__8_ DECAP_INV_G11
XG11343 XI11_2/XI0/XI0_41/d_7_ XI11_2/XI0/XI0_41/d__7_ DECAP_INV_G11
XG11344 XI11_2/XI0/XI0_41/d_6_ XI11_2/XI0/XI0_41/d__6_ DECAP_INV_G11
XG11345 XI11_2/XI0/XI0_41/d_5_ XI11_2/XI0/XI0_41/d__5_ DECAP_INV_G11
XG11346 XI11_2/XI0/XI0_41/d_4_ XI11_2/XI0/XI0_41/d__4_ DECAP_INV_G11
XG11347 XI11_2/XI0/XI0_41/d_3_ XI11_2/XI0/XI0_41/d__3_ DECAP_INV_G11
XG11348 XI11_2/XI0/XI0_41/d_2_ XI11_2/XI0/XI0_41/d__2_ DECAP_INV_G11
XG11349 XI11_2/XI0/XI0_41/d_1_ XI11_2/XI0/XI0_41/d__1_ DECAP_INV_G11
XG11350 XI11_2/XI0/XI0_41/d_0_ XI11_2/XI0/XI0_41/d__0_ DECAP_INV_G11
XG11351 XI11_2/XI0/XI0_40/d__15_ XI11_2/XI0/XI0_40/d_15_ DECAP_INV_G11
XG11352 XI11_2/XI0/XI0_40/d__14_ XI11_2/XI0/XI0_40/d_14_ DECAP_INV_G11
XG11353 XI11_2/XI0/XI0_40/d__13_ XI11_2/XI0/XI0_40/d_13_ DECAP_INV_G11
XG11354 XI11_2/XI0/XI0_40/d__12_ XI11_2/XI0/XI0_40/d_12_ DECAP_INV_G11
XG11355 XI11_2/XI0/XI0_40/d__11_ XI11_2/XI0/XI0_40/d_11_ DECAP_INV_G11
XG11356 XI11_2/XI0/XI0_40/d__10_ XI11_2/XI0/XI0_40/d_10_ DECAP_INV_G11
XG11357 XI11_2/XI0/XI0_40/d__9_ XI11_2/XI0/XI0_40/d_9_ DECAP_INV_G11
XG11358 XI11_2/XI0/XI0_40/d__8_ XI11_2/XI0/XI0_40/d_8_ DECAP_INV_G11
XG11359 XI11_2/XI0/XI0_40/d__7_ XI11_2/XI0/XI0_40/d_7_ DECAP_INV_G11
XG11360 XI11_2/XI0/XI0_40/d__6_ XI11_2/XI0/XI0_40/d_6_ DECAP_INV_G11
XG11361 XI11_2/XI0/XI0_40/d__5_ XI11_2/XI0/XI0_40/d_5_ DECAP_INV_G11
XG11362 XI11_2/XI0/XI0_40/d__4_ XI11_2/XI0/XI0_40/d_4_ DECAP_INV_G11
XG11363 XI11_2/XI0/XI0_40/d__3_ XI11_2/XI0/XI0_40/d_3_ DECAP_INV_G11
XG11364 XI11_2/XI0/XI0_40/d__2_ XI11_2/XI0/XI0_40/d_2_ DECAP_INV_G11
XG11365 XI11_2/XI0/XI0_40/d__1_ XI11_2/XI0/XI0_40/d_1_ DECAP_INV_G11
XG11366 XI11_2/XI0/XI0_40/d__0_ XI11_2/XI0/XI0_40/d_0_ DECAP_INV_G11
XG11367 XI11_2/XI0/XI0_40/d_15_ XI11_2/XI0/XI0_40/d__15_ DECAP_INV_G11
XG11368 XI11_2/XI0/XI0_40/d_14_ XI11_2/XI0/XI0_40/d__14_ DECAP_INV_G11
XG11369 XI11_2/XI0/XI0_40/d_13_ XI11_2/XI0/XI0_40/d__13_ DECAP_INV_G11
XG11370 XI11_2/XI0/XI0_40/d_12_ XI11_2/XI0/XI0_40/d__12_ DECAP_INV_G11
XG11371 XI11_2/XI0/XI0_40/d_11_ XI11_2/XI0/XI0_40/d__11_ DECAP_INV_G11
XG11372 XI11_2/XI0/XI0_40/d_10_ XI11_2/XI0/XI0_40/d__10_ DECAP_INV_G11
XG11373 XI11_2/XI0/XI0_40/d_9_ XI11_2/XI0/XI0_40/d__9_ DECAP_INV_G11
XG11374 XI11_2/XI0/XI0_40/d_8_ XI11_2/XI0/XI0_40/d__8_ DECAP_INV_G11
XG11375 XI11_2/XI0/XI0_40/d_7_ XI11_2/XI0/XI0_40/d__7_ DECAP_INV_G11
XG11376 XI11_2/XI0/XI0_40/d_6_ XI11_2/XI0/XI0_40/d__6_ DECAP_INV_G11
XG11377 XI11_2/XI0/XI0_40/d_5_ XI11_2/XI0/XI0_40/d__5_ DECAP_INV_G11
XG11378 XI11_2/XI0/XI0_40/d_4_ XI11_2/XI0/XI0_40/d__4_ DECAP_INV_G11
XG11379 XI11_2/XI0/XI0_40/d_3_ XI11_2/XI0/XI0_40/d__3_ DECAP_INV_G11
XG11380 XI11_2/XI0/XI0_40/d_2_ XI11_2/XI0/XI0_40/d__2_ DECAP_INV_G11
XG11381 XI11_2/XI0/XI0_40/d_1_ XI11_2/XI0/XI0_40/d__1_ DECAP_INV_G11
XG11382 XI11_2/XI0/XI0_40/d_0_ XI11_2/XI0/XI0_40/d__0_ DECAP_INV_G11
XG11383 XI11_2/XI0/XI0_39/d__15_ XI11_2/XI0/XI0_39/d_15_ DECAP_INV_G11
XG11384 XI11_2/XI0/XI0_39/d__14_ XI11_2/XI0/XI0_39/d_14_ DECAP_INV_G11
XG11385 XI11_2/XI0/XI0_39/d__13_ XI11_2/XI0/XI0_39/d_13_ DECAP_INV_G11
XG11386 XI11_2/XI0/XI0_39/d__12_ XI11_2/XI0/XI0_39/d_12_ DECAP_INV_G11
XG11387 XI11_2/XI0/XI0_39/d__11_ XI11_2/XI0/XI0_39/d_11_ DECAP_INV_G11
XG11388 XI11_2/XI0/XI0_39/d__10_ XI11_2/XI0/XI0_39/d_10_ DECAP_INV_G11
XG11389 XI11_2/XI0/XI0_39/d__9_ XI11_2/XI0/XI0_39/d_9_ DECAP_INV_G11
XG11390 XI11_2/XI0/XI0_39/d__8_ XI11_2/XI0/XI0_39/d_8_ DECAP_INV_G11
XG11391 XI11_2/XI0/XI0_39/d__7_ XI11_2/XI0/XI0_39/d_7_ DECAP_INV_G11
XG11392 XI11_2/XI0/XI0_39/d__6_ XI11_2/XI0/XI0_39/d_6_ DECAP_INV_G11
XG11393 XI11_2/XI0/XI0_39/d__5_ XI11_2/XI0/XI0_39/d_5_ DECAP_INV_G11
XG11394 XI11_2/XI0/XI0_39/d__4_ XI11_2/XI0/XI0_39/d_4_ DECAP_INV_G11
XG11395 XI11_2/XI0/XI0_39/d__3_ XI11_2/XI0/XI0_39/d_3_ DECAP_INV_G11
XG11396 XI11_2/XI0/XI0_39/d__2_ XI11_2/XI0/XI0_39/d_2_ DECAP_INV_G11
XG11397 XI11_2/XI0/XI0_39/d__1_ XI11_2/XI0/XI0_39/d_1_ DECAP_INV_G11
XG11398 XI11_2/XI0/XI0_39/d__0_ XI11_2/XI0/XI0_39/d_0_ DECAP_INV_G11
XG11399 XI11_2/XI0/XI0_39/d_15_ XI11_2/XI0/XI0_39/d__15_ DECAP_INV_G11
XG11400 XI11_2/XI0/XI0_39/d_14_ XI11_2/XI0/XI0_39/d__14_ DECAP_INV_G11
XG11401 XI11_2/XI0/XI0_39/d_13_ XI11_2/XI0/XI0_39/d__13_ DECAP_INV_G11
XG11402 XI11_2/XI0/XI0_39/d_12_ XI11_2/XI0/XI0_39/d__12_ DECAP_INV_G11
XG11403 XI11_2/XI0/XI0_39/d_11_ XI11_2/XI0/XI0_39/d__11_ DECAP_INV_G11
XG11404 XI11_2/XI0/XI0_39/d_10_ XI11_2/XI0/XI0_39/d__10_ DECAP_INV_G11
XG11405 XI11_2/XI0/XI0_39/d_9_ XI11_2/XI0/XI0_39/d__9_ DECAP_INV_G11
XG11406 XI11_2/XI0/XI0_39/d_8_ XI11_2/XI0/XI0_39/d__8_ DECAP_INV_G11
XG11407 XI11_2/XI0/XI0_39/d_7_ XI11_2/XI0/XI0_39/d__7_ DECAP_INV_G11
XG11408 XI11_2/XI0/XI0_39/d_6_ XI11_2/XI0/XI0_39/d__6_ DECAP_INV_G11
XG11409 XI11_2/XI0/XI0_39/d_5_ XI11_2/XI0/XI0_39/d__5_ DECAP_INV_G11
XG11410 XI11_2/XI0/XI0_39/d_4_ XI11_2/XI0/XI0_39/d__4_ DECAP_INV_G11
XG11411 XI11_2/XI0/XI0_39/d_3_ XI11_2/XI0/XI0_39/d__3_ DECAP_INV_G11
XG11412 XI11_2/XI0/XI0_39/d_2_ XI11_2/XI0/XI0_39/d__2_ DECAP_INV_G11
XG11413 XI11_2/XI0/XI0_39/d_1_ XI11_2/XI0/XI0_39/d__1_ DECAP_INV_G11
XG11414 XI11_2/XI0/XI0_39/d_0_ XI11_2/XI0/XI0_39/d__0_ DECAP_INV_G11
XG11415 XI11_2/XI0/XI0_38/d__15_ XI11_2/XI0/XI0_38/d_15_ DECAP_INV_G11
XG11416 XI11_2/XI0/XI0_38/d__14_ XI11_2/XI0/XI0_38/d_14_ DECAP_INV_G11
XG11417 XI11_2/XI0/XI0_38/d__13_ XI11_2/XI0/XI0_38/d_13_ DECAP_INV_G11
XG11418 XI11_2/XI0/XI0_38/d__12_ XI11_2/XI0/XI0_38/d_12_ DECAP_INV_G11
XG11419 XI11_2/XI0/XI0_38/d__11_ XI11_2/XI0/XI0_38/d_11_ DECAP_INV_G11
XG11420 XI11_2/XI0/XI0_38/d__10_ XI11_2/XI0/XI0_38/d_10_ DECAP_INV_G11
XG11421 XI11_2/XI0/XI0_38/d__9_ XI11_2/XI0/XI0_38/d_9_ DECAP_INV_G11
XG11422 XI11_2/XI0/XI0_38/d__8_ XI11_2/XI0/XI0_38/d_8_ DECAP_INV_G11
XG11423 XI11_2/XI0/XI0_38/d__7_ XI11_2/XI0/XI0_38/d_7_ DECAP_INV_G11
XG11424 XI11_2/XI0/XI0_38/d__6_ XI11_2/XI0/XI0_38/d_6_ DECAP_INV_G11
XG11425 XI11_2/XI0/XI0_38/d__5_ XI11_2/XI0/XI0_38/d_5_ DECAP_INV_G11
XG11426 XI11_2/XI0/XI0_38/d__4_ XI11_2/XI0/XI0_38/d_4_ DECAP_INV_G11
XG11427 XI11_2/XI0/XI0_38/d__3_ XI11_2/XI0/XI0_38/d_3_ DECAP_INV_G11
XG11428 XI11_2/XI0/XI0_38/d__2_ XI11_2/XI0/XI0_38/d_2_ DECAP_INV_G11
XG11429 XI11_2/XI0/XI0_38/d__1_ XI11_2/XI0/XI0_38/d_1_ DECAP_INV_G11
XG11430 XI11_2/XI0/XI0_38/d__0_ XI11_2/XI0/XI0_38/d_0_ DECAP_INV_G11
XG11431 XI11_2/XI0/XI0_38/d_15_ XI11_2/XI0/XI0_38/d__15_ DECAP_INV_G11
XG11432 XI11_2/XI0/XI0_38/d_14_ XI11_2/XI0/XI0_38/d__14_ DECAP_INV_G11
XG11433 XI11_2/XI0/XI0_38/d_13_ XI11_2/XI0/XI0_38/d__13_ DECAP_INV_G11
XG11434 XI11_2/XI0/XI0_38/d_12_ XI11_2/XI0/XI0_38/d__12_ DECAP_INV_G11
XG11435 XI11_2/XI0/XI0_38/d_11_ XI11_2/XI0/XI0_38/d__11_ DECAP_INV_G11
XG11436 XI11_2/XI0/XI0_38/d_10_ XI11_2/XI0/XI0_38/d__10_ DECAP_INV_G11
XG11437 XI11_2/XI0/XI0_38/d_9_ XI11_2/XI0/XI0_38/d__9_ DECAP_INV_G11
XG11438 XI11_2/XI0/XI0_38/d_8_ XI11_2/XI0/XI0_38/d__8_ DECAP_INV_G11
XG11439 XI11_2/XI0/XI0_38/d_7_ XI11_2/XI0/XI0_38/d__7_ DECAP_INV_G11
XG11440 XI11_2/XI0/XI0_38/d_6_ XI11_2/XI0/XI0_38/d__6_ DECAP_INV_G11
XG11441 XI11_2/XI0/XI0_38/d_5_ XI11_2/XI0/XI0_38/d__5_ DECAP_INV_G11
XG11442 XI11_2/XI0/XI0_38/d_4_ XI11_2/XI0/XI0_38/d__4_ DECAP_INV_G11
XG11443 XI11_2/XI0/XI0_38/d_3_ XI11_2/XI0/XI0_38/d__3_ DECAP_INV_G11
XG11444 XI11_2/XI0/XI0_38/d_2_ XI11_2/XI0/XI0_38/d__2_ DECAP_INV_G11
XG11445 XI11_2/XI0/XI0_38/d_1_ XI11_2/XI0/XI0_38/d__1_ DECAP_INV_G11
XG11446 XI11_2/XI0/XI0_38/d_0_ XI11_2/XI0/XI0_38/d__0_ DECAP_INV_G11
XG11447 XI11_2/XI0/XI0_37/d__15_ XI11_2/XI0/XI0_37/d_15_ DECAP_INV_G11
XG11448 XI11_2/XI0/XI0_37/d__14_ XI11_2/XI0/XI0_37/d_14_ DECAP_INV_G11
XG11449 XI11_2/XI0/XI0_37/d__13_ XI11_2/XI0/XI0_37/d_13_ DECAP_INV_G11
XG11450 XI11_2/XI0/XI0_37/d__12_ XI11_2/XI0/XI0_37/d_12_ DECAP_INV_G11
XG11451 XI11_2/XI0/XI0_37/d__11_ XI11_2/XI0/XI0_37/d_11_ DECAP_INV_G11
XG11452 XI11_2/XI0/XI0_37/d__10_ XI11_2/XI0/XI0_37/d_10_ DECAP_INV_G11
XG11453 XI11_2/XI0/XI0_37/d__9_ XI11_2/XI0/XI0_37/d_9_ DECAP_INV_G11
XG11454 XI11_2/XI0/XI0_37/d__8_ XI11_2/XI0/XI0_37/d_8_ DECAP_INV_G11
XG11455 XI11_2/XI0/XI0_37/d__7_ XI11_2/XI0/XI0_37/d_7_ DECAP_INV_G11
XG11456 XI11_2/XI0/XI0_37/d__6_ XI11_2/XI0/XI0_37/d_6_ DECAP_INV_G11
XG11457 XI11_2/XI0/XI0_37/d__5_ XI11_2/XI0/XI0_37/d_5_ DECAP_INV_G11
XG11458 XI11_2/XI0/XI0_37/d__4_ XI11_2/XI0/XI0_37/d_4_ DECAP_INV_G11
XG11459 XI11_2/XI0/XI0_37/d__3_ XI11_2/XI0/XI0_37/d_3_ DECAP_INV_G11
XG11460 XI11_2/XI0/XI0_37/d__2_ XI11_2/XI0/XI0_37/d_2_ DECAP_INV_G11
XG11461 XI11_2/XI0/XI0_37/d__1_ XI11_2/XI0/XI0_37/d_1_ DECAP_INV_G11
XG11462 XI11_2/XI0/XI0_37/d__0_ XI11_2/XI0/XI0_37/d_0_ DECAP_INV_G11
XG11463 XI11_2/XI0/XI0_37/d_15_ XI11_2/XI0/XI0_37/d__15_ DECAP_INV_G11
XG11464 XI11_2/XI0/XI0_37/d_14_ XI11_2/XI0/XI0_37/d__14_ DECAP_INV_G11
XG11465 XI11_2/XI0/XI0_37/d_13_ XI11_2/XI0/XI0_37/d__13_ DECAP_INV_G11
XG11466 XI11_2/XI0/XI0_37/d_12_ XI11_2/XI0/XI0_37/d__12_ DECAP_INV_G11
XG11467 XI11_2/XI0/XI0_37/d_11_ XI11_2/XI0/XI0_37/d__11_ DECAP_INV_G11
XG11468 XI11_2/XI0/XI0_37/d_10_ XI11_2/XI0/XI0_37/d__10_ DECAP_INV_G11
XG11469 XI11_2/XI0/XI0_37/d_9_ XI11_2/XI0/XI0_37/d__9_ DECAP_INV_G11
XG11470 XI11_2/XI0/XI0_37/d_8_ XI11_2/XI0/XI0_37/d__8_ DECAP_INV_G11
XG11471 XI11_2/XI0/XI0_37/d_7_ XI11_2/XI0/XI0_37/d__7_ DECAP_INV_G11
XG11472 XI11_2/XI0/XI0_37/d_6_ XI11_2/XI0/XI0_37/d__6_ DECAP_INV_G11
XG11473 XI11_2/XI0/XI0_37/d_5_ XI11_2/XI0/XI0_37/d__5_ DECAP_INV_G11
XG11474 XI11_2/XI0/XI0_37/d_4_ XI11_2/XI0/XI0_37/d__4_ DECAP_INV_G11
XG11475 XI11_2/XI0/XI0_37/d_3_ XI11_2/XI0/XI0_37/d__3_ DECAP_INV_G11
XG11476 XI11_2/XI0/XI0_37/d_2_ XI11_2/XI0/XI0_37/d__2_ DECAP_INV_G11
XG11477 XI11_2/XI0/XI0_37/d_1_ XI11_2/XI0/XI0_37/d__1_ DECAP_INV_G11
XG11478 XI11_2/XI0/XI0_37/d_0_ XI11_2/XI0/XI0_37/d__0_ DECAP_INV_G11
XG11479 XI11_2/XI0/XI0_36/d__15_ XI11_2/XI0/XI0_36/d_15_ DECAP_INV_G11
XG11480 XI11_2/XI0/XI0_36/d__14_ XI11_2/XI0/XI0_36/d_14_ DECAP_INV_G11
XG11481 XI11_2/XI0/XI0_36/d__13_ XI11_2/XI0/XI0_36/d_13_ DECAP_INV_G11
XG11482 XI11_2/XI0/XI0_36/d__12_ XI11_2/XI0/XI0_36/d_12_ DECAP_INV_G11
XG11483 XI11_2/XI0/XI0_36/d__11_ XI11_2/XI0/XI0_36/d_11_ DECAP_INV_G11
XG11484 XI11_2/XI0/XI0_36/d__10_ XI11_2/XI0/XI0_36/d_10_ DECAP_INV_G11
XG11485 XI11_2/XI0/XI0_36/d__9_ XI11_2/XI0/XI0_36/d_9_ DECAP_INV_G11
XG11486 XI11_2/XI0/XI0_36/d__8_ XI11_2/XI0/XI0_36/d_8_ DECAP_INV_G11
XG11487 XI11_2/XI0/XI0_36/d__7_ XI11_2/XI0/XI0_36/d_7_ DECAP_INV_G11
XG11488 XI11_2/XI0/XI0_36/d__6_ XI11_2/XI0/XI0_36/d_6_ DECAP_INV_G11
XG11489 XI11_2/XI0/XI0_36/d__5_ XI11_2/XI0/XI0_36/d_5_ DECAP_INV_G11
XG11490 XI11_2/XI0/XI0_36/d__4_ XI11_2/XI0/XI0_36/d_4_ DECAP_INV_G11
XG11491 XI11_2/XI0/XI0_36/d__3_ XI11_2/XI0/XI0_36/d_3_ DECAP_INV_G11
XG11492 XI11_2/XI0/XI0_36/d__2_ XI11_2/XI0/XI0_36/d_2_ DECAP_INV_G11
XG11493 XI11_2/XI0/XI0_36/d__1_ XI11_2/XI0/XI0_36/d_1_ DECAP_INV_G11
XG11494 XI11_2/XI0/XI0_36/d__0_ XI11_2/XI0/XI0_36/d_0_ DECAP_INV_G11
XG11495 XI11_2/XI0/XI0_36/d_15_ XI11_2/XI0/XI0_36/d__15_ DECAP_INV_G11
XG11496 XI11_2/XI0/XI0_36/d_14_ XI11_2/XI0/XI0_36/d__14_ DECAP_INV_G11
XG11497 XI11_2/XI0/XI0_36/d_13_ XI11_2/XI0/XI0_36/d__13_ DECAP_INV_G11
XG11498 XI11_2/XI0/XI0_36/d_12_ XI11_2/XI0/XI0_36/d__12_ DECAP_INV_G11
XG11499 XI11_2/XI0/XI0_36/d_11_ XI11_2/XI0/XI0_36/d__11_ DECAP_INV_G11
XG11500 XI11_2/XI0/XI0_36/d_10_ XI11_2/XI0/XI0_36/d__10_ DECAP_INV_G11
XG11501 XI11_2/XI0/XI0_36/d_9_ XI11_2/XI0/XI0_36/d__9_ DECAP_INV_G11
XG11502 XI11_2/XI0/XI0_36/d_8_ XI11_2/XI0/XI0_36/d__8_ DECAP_INV_G11
XG11503 XI11_2/XI0/XI0_36/d_7_ XI11_2/XI0/XI0_36/d__7_ DECAP_INV_G11
XG11504 XI11_2/XI0/XI0_36/d_6_ XI11_2/XI0/XI0_36/d__6_ DECAP_INV_G11
XG11505 XI11_2/XI0/XI0_36/d_5_ XI11_2/XI0/XI0_36/d__5_ DECAP_INV_G11
XG11506 XI11_2/XI0/XI0_36/d_4_ XI11_2/XI0/XI0_36/d__4_ DECAP_INV_G11
XG11507 XI11_2/XI0/XI0_36/d_3_ XI11_2/XI0/XI0_36/d__3_ DECAP_INV_G11
XG11508 XI11_2/XI0/XI0_36/d_2_ XI11_2/XI0/XI0_36/d__2_ DECAP_INV_G11
XG11509 XI11_2/XI0/XI0_36/d_1_ XI11_2/XI0/XI0_36/d__1_ DECAP_INV_G11
XG11510 XI11_2/XI0/XI0_36/d_0_ XI11_2/XI0/XI0_36/d__0_ DECAP_INV_G11
XG11511 XI11_2/XI0/XI0_35/d__15_ XI11_2/XI0/XI0_35/d_15_ DECAP_INV_G11
XG11512 XI11_2/XI0/XI0_35/d__14_ XI11_2/XI0/XI0_35/d_14_ DECAP_INV_G11
XG11513 XI11_2/XI0/XI0_35/d__13_ XI11_2/XI0/XI0_35/d_13_ DECAP_INV_G11
XG11514 XI11_2/XI0/XI0_35/d__12_ XI11_2/XI0/XI0_35/d_12_ DECAP_INV_G11
XG11515 XI11_2/XI0/XI0_35/d__11_ XI11_2/XI0/XI0_35/d_11_ DECAP_INV_G11
XG11516 XI11_2/XI0/XI0_35/d__10_ XI11_2/XI0/XI0_35/d_10_ DECAP_INV_G11
XG11517 XI11_2/XI0/XI0_35/d__9_ XI11_2/XI0/XI0_35/d_9_ DECAP_INV_G11
XG11518 XI11_2/XI0/XI0_35/d__8_ XI11_2/XI0/XI0_35/d_8_ DECAP_INV_G11
XG11519 XI11_2/XI0/XI0_35/d__7_ XI11_2/XI0/XI0_35/d_7_ DECAP_INV_G11
XG11520 XI11_2/XI0/XI0_35/d__6_ XI11_2/XI0/XI0_35/d_6_ DECAP_INV_G11
XG11521 XI11_2/XI0/XI0_35/d__5_ XI11_2/XI0/XI0_35/d_5_ DECAP_INV_G11
XG11522 XI11_2/XI0/XI0_35/d__4_ XI11_2/XI0/XI0_35/d_4_ DECAP_INV_G11
XG11523 XI11_2/XI0/XI0_35/d__3_ XI11_2/XI0/XI0_35/d_3_ DECAP_INV_G11
XG11524 XI11_2/XI0/XI0_35/d__2_ XI11_2/XI0/XI0_35/d_2_ DECAP_INV_G11
XG11525 XI11_2/XI0/XI0_35/d__1_ XI11_2/XI0/XI0_35/d_1_ DECAP_INV_G11
XG11526 XI11_2/XI0/XI0_35/d__0_ XI11_2/XI0/XI0_35/d_0_ DECAP_INV_G11
XG11527 XI11_2/XI0/XI0_35/d_15_ XI11_2/XI0/XI0_35/d__15_ DECAP_INV_G11
XG11528 XI11_2/XI0/XI0_35/d_14_ XI11_2/XI0/XI0_35/d__14_ DECAP_INV_G11
XG11529 XI11_2/XI0/XI0_35/d_13_ XI11_2/XI0/XI0_35/d__13_ DECAP_INV_G11
XG11530 XI11_2/XI0/XI0_35/d_12_ XI11_2/XI0/XI0_35/d__12_ DECAP_INV_G11
XG11531 XI11_2/XI0/XI0_35/d_11_ XI11_2/XI0/XI0_35/d__11_ DECAP_INV_G11
XG11532 XI11_2/XI0/XI0_35/d_10_ XI11_2/XI0/XI0_35/d__10_ DECAP_INV_G11
XG11533 XI11_2/XI0/XI0_35/d_9_ XI11_2/XI0/XI0_35/d__9_ DECAP_INV_G11
XG11534 XI11_2/XI0/XI0_35/d_8_ XI11_2/XI0/XI0_35/d__8_ DECAP_INV_G11
XG11535 XI11_2/XI0/XI0_35/d_7_ XI11_2/XI0/XI0_35/d__7_ DECAP_INV_G11
XG11536 XI11_2/XI0/XI0_35/d_6_ XI11_2/XI0/XI0_35/d__6_ DECAP_INV_G11
XG11537 XI11_2/XI0/XI0_35/d_5_ XI11_2/XI0/XI0_35/d__5_ DECAP_INV_G11
XG11538 XI11_2/XI0/XI0_35/d_4_ XI11_2/XI0/XI0_35/d__4_ DECAP_INV_G11
XG11539 XI11_2/XI0/XI0_35/d_3_ XI11_2/XI0/XI0_35/d__3_ DECAP_INV_G11
XG11540 XI11_2/XI0/XI0_35/d_2_ XI11_2/XI0/XI0_35/d__2_ DECAP_INV_G11
XG11541 XI11_2/XI0/XI0_35/d_1_ XI11_2/XI0/XI0_35/d__1_ DECAP_INV_G11
XG11542 XI11_2/XI0/XI0_35/d_0_ XI11_2/XI0/XI0_35/d__0_ DECAP_INV_G11
XG11543 XI11_2/XI0/XI0_34/d__15_ XI11_2/XI0/XI0_34/d_15_ DECAP_INV_G11
XG11544 XI11_2/XI0/XI0_34/d__14_ XI11_2/XI0/XI0_34/d_14_ DECAP_INV_G11
XG11545 XI11_2/XI0/XI0_34/d__13_ XI11_2/XI0/XI0_34/d_13_ DECAP_INV_G11
XG11546 XI11_2/XI0/XI0_34/d__12_ XI11_2/XI0/XI0_34/d_12_ DECAP_INV_G11
XG11547 XI11_2/XI0/XI0_34/d__11_ XI11_2/XI0/XI0_34/d_11_ DECAP_INV_G11
XG11548 XI11_2/XI0/XI0_34/d__10_ XI11_2/XI0/XI0_34/d_10_ DECAP_INV_G11
XG11549 XI11_2/XI0/XI0_34/d__9_ XI11_2/XI0/XI0_34/d_9_ DECAP_INV_G11
XG11550 XI11_2/XI0/XI0_34/d__8_ XI11_2/XI0/XI0_34/d_8_ DECAP_INV_G11
XG11551 XI11_2/XI0/XI0_34/d__7_ XI11_2/XI0/XI0_34/d_7_ DECAP_INV_G11
XG11552 XI11_2/XI0/XI0_34/d__6_ XI11_2/XI0/XI0_34/d_6_ DECAP_INV_G11
XG11553 XI11_2/XI0/XI0_34/d__5_ XI11_2/XI0/XI0_34/d_5_ DECAP_INV_G11
XG11554 XI11_2/XI0/XI0_34/d__4_ XI11_2/XI0/XI0_34/d_4_ DECAP_INV_G11
XG11555 XI11_2/XI0/XI0_34/d__3_ XI11_2/XI0/XI0_34/d_3_ DECAP_INV_G11
XG11556 XI11_2/XI0/XI0_34/d__2_ XI11_2/XI0/XI0_34/d_2_ DECAP_INV_G11
XG11557 XI11_2/XI0/XI0_34/d__1_ XI11_2/XI0/XI0_34/d_1_ DECAP_INV_G11
XG11558 XI11_2/XI0/XI0_34/d__0_ XI11_2/XI0/XI0_34/d_0_ DECAP_INV_G11
XG11559 XI11_2/XI0/XI0_34/d_15_ XI11_2/XI0/XI0_34/d__15_ DECAP_INV_G11
XG11560 XI11_2/XI0/XI0_34/d_14_ XI11_2/XI0/XI0_34/d__14_ DECAP_INV_G11
XG11561 XI11_2/XI0/XI0_34/d_13_ XI11_2/XI0/XI0_34/d__13_ DECAP_INV_G11
XG11562 XI11_2/XI0/XI0_34/d_12_ XI11_2/XI0/XI0_34/d__12_ DECAP_INV_G11
XG11563 XI11_2/XI0/XI0_34/d_11_ XI11_2/XI0/XI0_34/d__11_ DECAP_INV_G11
XG11564 XI11_2/XI0/XI0_34/d_10_ XI11_2/XI0/XI0_34/d__10_ DECAP_INV_G11
XG11565 XI11_2/XI0/XI0_34/d_9_ XI11_2/XI0/XI0_34/d__9_ DECAP_INV_G11
XG11566 XI11_2/XI0/XI0_34/d_8_ XI11_2/XI0/XI0_34/d__8_ DECAP_INV_G11
XG11567 XI11_2/XI0/XI0_34/d_7_ XI11_2/XI0/XI0_34/d__7_ DECAP_INV_G11
XG11568 XI11_2/XI0/XI0_34/d_6_ XI11_2/XI0/XI0_34/d__6_ DECAP_INV_G11
XG11569 XI11_2/XI0/XI0_34/d_5_ XI11_2/XI0/XI0_34/d__5_ DECAP_INV_G11
XG11570 XI11_2/XI0/XI0_34/d_4_ XI11_2/XI0/XI0_34/d__4_ DECAP_INV_G11
XG11571 XI11_2/XI0/XI0_34/d_3_ XI11_2/XI0/XI0_34/d__3_ DECAP_INV_G11
XG11572 XI11_2/XI0/XI0_34/d_2_ XI11_2/XI0/XI0_34/d__2_ DECAP_INV_G11
XG11573 XI11_2/XI0/XI0_34/d_1_ XI11_2/XI0/XI0_34/d__1_ DECAP_INV_G11
XG11574 XI11_2/XI0/XI0_34/d_0_ XI11_2/XI0/XI0_34/d__0_ DECAP_INV_G11
XG11575 XI11_2/XI0/XI0_33/d__15_ XI11_2/XI0/XI0_33/d_15_ DECAP_INV_G11
XG11576 XI11_2/XI0/XI0_33/d__14_ XI11_2/XI0/XI0_33/d_14_ DECAP_INV_G11
XG11577 XI11_2/XI0/XI0_33/d__13_ XI11_2/XI0/XI0_33/d_13_ DECAP_INV_G11
XG11578 XI11_2/XI0/XI0_33/d__12_ XI11_2/XI0/XI0_33/d_12_ DECAP_INV_G11
XG11579 XI11_2/XI0/XI0_33/d__11_ XI11_2/XI0/XI0_33/d_11_ DECAP_INV_G11
XG11580 XI11_2/XI0/XI0_33/d__10_ XI11_2/XI0/XI0_33/d_10_ DECAP_INV_G11
XG11581 XI11_2/XI0/XI0_33/d__9_ XI11_2/XI0/XI0_33/d_9_ DECAP_INV_G11
XG11582 XI11_2/XI0/XI0_33/d__8_ XI11_2/XI0/XI0_33/d_8_ DECAP_INV_G11
XG11583 XI11_2/XI0/XI0_33/d__7_ XI11_2/XI0/XI0_33/d_7_ DECAP_INV_G11
XG11584 XI11_2/XI0/XI0_33/d__6_ XI11_2/XI0/XI0_33/d_6_ DECAP_INV_G11
XG11585 XI11_2/XI0/XI0_33/d__5_ XI11_2/XI0/XI0_33/d_5_ DECAP_INV_G11
XG11586 XI11_2/XI0/XI0_33/d__4_ XI11_2/XI0/XI0_33/d_4_ DECAP_INV_G11
XG11587 XI11_2/XI0/XI0_33/d__3_ XI11_2/XI0/XI0_33/d_3_ DECAP_INV_G11
XG11588 XI11_2/XI0/XI0_33/d__2_ XI11_2/XI0/XI0_33/d_2_ DECAP_INV_G11
XG11589 XI11_2/XI0/XI0_33/d__1_ XI11_2/XI0/XI0_33/d_1_ DECAP_INV_G11
XG11590 XI11_2/XI0/XI0_33/d__0_ XI11_2/XI0/XI0_33/d_0_ DECAP_INV_G11
XG11591 XI11_2/XI0/XI0_33/d_15_ XI11_2/XI0/XI0_33/d__15_ DECAP_INV_G11
XG11592 XI11_2/XI0/XI0_33/d_14_ XI11_2/XI0/XI0_33/d__14_ DECAP_INV_G11
XG11593 XI11_2/XI0/XI0_33/d_13_ XI11_2/XI0/XI0_33/d__13_ DECAP_INV_G11
XG11594 XI11_2/XI0/XI0_33/d_12_ XI11_2/XI0/XI0_33/d__12_ DECAP_INV_G11
XG11595 XI11_2/XI0/XI0_33/d_11_ XI11_2/XI0/XI0_33/d__11_ DECAP_INV_G11
XG11596 XI11_2/XI0/XI0_33/d_10_ XI11_2/XI0/XI0_33/d__10_ DECAP_INV_G11
XG11597 XI11_2/XI0/XI0_33/d_9_ XI11_2/XI0/XI0_33/d__9_ DECAP_INV_G11
XG11598 XI11_2/XI0/XI0_33/d_8_ XI11_2/XI0/XI0_33/d__8_ DECAP_INV_G11
XG11599 XI11_2/XI0/XI0_33/d_7_ XI11_2/XI0/XI0_33/d__7_ DECAP_INV_G11
XG11600 XI11_2/XI0/XI0_33/d_6_ XI11_2/XI0/XI0_33/d__6_ DECAP_INV_G11
XG11601 XI11_2/XI0/XI0_33/d_5_ XI11_2/XI0/XI0_33/d__5_ DECAP_INV_G11
XG11602 XI11_2/XI0/XI0_33/d_4_ XI11_2/XI0/XI0_33/d__4_ DECAP_INV_G11
XG11603 XI11_2/XI0/XI0_33/d_3_ XI11_2/XI0/XI0_33/d__3_ DECAP_INV_G11
XG11604 XI11_2/XI0/XI0_33/d_2_ XI11_2/XI0/XI0_33/d__2_ DECAP_INV_G11
XG11605 XI11_2/XI0/XI0_33/d_1_ XI11_2/XI0/XI0_33/d__1_ DECAP_INV_G11
XG11606 XI11_2/XI0/XI0_33/d_0_ XI11_2/XI0/XI0_33/d__0_ DECAP_INV_G11
XG11607 XI11_2/XI0/XI0_32/d__15_ XI11_2/XI0/XI0_32/d_15_ DECAP_INV_G11
XG11608 XI11_2/XI0/XI0_32/d__14_ XI11_2/XI0/XI0_32/d_14_ DECAP_INV_G11
XG11609 XI11_2/XI0/XI0_32/d__13_ XI11_2/XI0/XI0_32/d_13_ DECAP_INV_G11
XG11610 XI11_2/XI0/XI0_32/d__12_ XI11_2/XI0/XI0_32/d_12_ DECAP_INV_G11
XG11611 XI11_2/XI0/XI0_32/d__11_ XI11_2/XI0/XI0_32/d_11_ DECAP_INV_G11
XG11612 XI11_2/XI0/XI0_32/d__10_ XI11_2/XI0/XI0_32/d_10_ DECAP_INV_G11
XG11613 XI11_2/XI0/XI0_32/d__9_ XI11_2/XI0/XI0_32/d_9_ DECAP_INV_G11
XG11614 XI11_2/XI0/XI0_32/d__8_ XI11_2/XI0/XI0_32/d_8_ DECAP_INV_G11
XG11615 XI11_2/XI0/XI0_32/d__7_ XI11_2/XI0/XI0_32/d_7_ DECAP_INV_G11
XG11616 XI11_2/XI0/XI0_32/d__6_ XI11_2/XI0/XI0_32/d_6_ DECAP_INV_G11
XG11617 XI11_2/XI0/XI0_32/d__5_ XI11_2/XI0/XI0_32/d_5_ DECAP_INV_G11
XG11618 XI11_2/XI0/XI0_32/d__4_ XI11_2/XI0/XI0_32/d_4_ DECAP_INV_G11
XG11619 XI11_2/XI0/XI0_32/d__3_ XI11_2/XI0/XI0_32/d_3_ DECAP_INV_G11
XG11620 XI11_2/XI0/XI0_32/d__2_ XI11_2/XI0/XI0_32/d_2_ DECAP_INV_G11
XG11621 XI11_2/XI0/XI0_32/d__1_ XI11_2/XI0/XI0_32/d_1_ DECAP_INV_G11
XG11622 XI11_2/XI0/XI0_32/d__0_ XI11_2/XI0/XI0_32/d_0_ DECAP_INV_G11
XG11623 XI11_2/XI0/XI0_32/d_15_ XI11_2/XI0/XI0_32/d__15_ DECAP_INV_G11
XG11624 XI11_2/XI0/XI0_32/d_14_ XI11_2/XI0/XI0_32/d__14_ DECAP_INV_G11
XG11625 XI11_2/XI0/XI0_32/d_13_ XI11_2/XI0/XI0_32/d__13_ DECAP_INV_G11
XG11626 XI11_2/XI0/XI0_32/d_12_ XI11_2/XI0/XI0_32/d__12_ DECAP_INV_G11
XG11627 XI11_2/XI0/XI0_32/d_11_ XI11_2/XI0/XI0_32/d__11_ DECAP_INV_G11
XG11628 XI11_2/XI0/XI0_32/d_10_ XI11_2/XI0/XI0_32/d__10_ DECAP_INV_G11
XG11629 XI11_2/XI0/XI0_32/d_9_ XI11_2/XI0/XI0_32/d__9_ DECAP_INV_G11
XG11630 XI11_2/XI0/XI0_32/d_8_ XI11_2/XI0/XI0_32/d__8_ DECAP_INV_G11
XG11631 XI11_2/XI0/XI0_32/d_7_ XI11_2/XI0/XI0_32/d__7_ DECAP_INV_G11
XG11632 XI11_2/XI0/XI0_32/d_6_ XI11_2/XI0/XI0_32/d__6_ DECAP_INV_G11
XG11633 XI11_2/XI0/XI0_32/d_5_ XI11_2/XI0/XI0_32/d__5_ DECAP_INV_G11
XG11634 XI11_2/XI0/XI0_32/d_4_ XI11_2/XI0/XI0_32/d__4_ DECAP_INV_G11
XG11635 XI11_2/XI0/XI0_32/d_3_ XI11_2/XI0/XI0_32/d__3_ DECAP_INV_G11
XG11636 XI11_2/XI0/XI0_32/d_2_ XI11_2/XI0/XI0_32/d__2_ DECAP_INV_G11
XG11637 XI11_2/XI0/XI0_32/d_1_ XI11_2/XI0/XI0_32/d__1_ DECAP_INV_G11
XG11638 XI11_2/XI0/XI0_32/d_0_ XI11_2/XI0/XI0_32/d__0_ DECAP_INV_G11
XG11639 XI11_2/XI0/XI0_31/d__15_ XI11_2/XI0/XI0_31/d_15_ DECAP_INV_G11
XG11640 XI11_2/XI0/XI0_31/d__14_ XI11_2/XI0/XI0_31/d_14_ DECAP_INV_G11
XG11641 XI11_2/XI0/XI0_31/d__13_ XI11_2/XI0/XI0_31/d_13_ DECAP_INV_G11
XG11642 XI11_2/XI0/XI0_31/d__12_ XI11_2/XI0/XI0_31/d_12_ DECAP_INV_G11
XG11643 XI11_2/XI0/XI0_31/d__11_ XI11_2/XI0/XI0_31/d_11_ DECAP_INV_G11
XG11644 XI11_2/XI0/XI0_31/d__10_ XI11_2/XI0/XI0_31/d_10_ DECAP_INV_G11
XG11645 XI11_2/XI0/XI0_31/d__9_ XI11_2/XI0/XI0_31/d_9_ DECAP_INV_G11
XG11646 XI11_2/XI0/XI0_31/d__8_ XI11_2/XI0/XI0_31/d_8_ DECAP_INV_G11
XG11647 XI11_2/XI0/XI0_31/d__7_ XI11_2/XI0/XI0_31/d_7_ DECAP_INV_G11
XG11648 XI11_2/XI0/XI0_31/d__6_ XI11_2/XI0/XI0_31/d_6_ DECAP_INV_G11
XG11649 XI11_2/XI0/XI0_31/d__5_ XI11_2/XI0/XI0_31/d_5_ DECAP_INV_G11
XG11650 XI11_2/XI0/XI0_31/d__4_ XI11_2/XI0/XI0_31/d_4_ DECAP_INV_G11
XG11651 XI11_2/XI0/XI0_31/d__3_ XI11_2/XI0/XI0_31/d_3_ DECAP_INV_G11
XG11652 XI11_2/XI0/XI0_31/d__2_ XI11_2/XI0/XI0_31/d_2_ DECAP_INV_G11
XG11653 XI11_2/XI0/XI0_31/d__1_ XI11_2/XI0/XI0_31/d_1_ DECAP_INV_G11
XG11654 XI11_2/XI0/XI0_31/d__0_ XI11_2/XI0/XI0_31/d_0_ DECAP_INV_G11
XG11655 XI11_2/XI0/XI0_31/d_15_ XI11_2/XI0/XI0_31/d__15_ DECAP_INV_G11
XG11656 XI11_2/XI0/XI0_31/d_14_ XI11_2/XI0/XI0_31/d__14_ DECAP_INV_G11
XG11657 XI11_2/XI0/XI0_31/d_13_ XI11_2/XI0/XI0_31/d__13_ DECAP_INV_G11
XG11658 XI11_2/XI0/XI0_31/d_12_ XI11_2/XI0/XI0_31/d__12_ DECAP_INV_G11
XG11659 XI11_2/XI0/XI0_31/d_11_ XI11_2/XI0/XI0_31/d__11_ DECAP_INV_G11
XG11660 XI11_2/XI0/XI0_31/d_10_ XI11_2/XI0/XI0_31/d__10_ DECAP_INV_G11
XG11661 XI11_2/XI0/XI0_31/d_9_ XI11_2/XI0/XI0_31/d__9_ DECAP_INV_G11
XG11662 XI11_2/XI0/XI0_31/d_8_ XI11_2/XI0/XI0_31/d__8_ DECAP_INV_G11
XG11663 XI11_2/XI0/XI0_31/d_7_ XI11_2/XI0/XI0_31/d__7_ DECAP_INV_G11
XG11664 XI11_2/XI0/XI0_31/d_6_ XI11_2/XI0/XI0_31/d__6_ DECAP_INV_G11
XG11665 XI11_2/XI0/XI0_31/d_5_ XI11_2/XI0/XI0_31/d__5_ DECAP_INV_G11
XG11666 XI11_2/XI0/XI0_31/d_4_ XI11_2/XI0/XI0_31/d__4_ DECAP_INV_G11
XG11667 XI11_2/XI0/XI0_31/d_3_ XI11_2/XI0/XI0_31/d__3_ DECAP_INV_G11
XG11668 XI11_2/XI0/XI0_31/d_2_ XI11_2/XI0/XI0_31/d__2_ DECAP_INV_G11
XG11669 XI11_2/XI0/XI0_31/d_1_ XI11_2/XI0/XI0_31/d__1_ DECAP_INV_G11
XG11670 XI11_2/XI0/XI0_31/d_0_ XI11_2/XI0/XI0_31/d__0_ DECAP_INV_G11
XG11671 XI11_2/XI0/XI0_30/d__15_ XI11_2/XI0/XI0_30/d_15_ DECAP_INV_G11
XG11672 XI11_2/XI0/XI0_30/d__14_ XI11_2/XI0/XI0_30/d_14_ DECAP_INV_G11
XG11673 XI11_2/XI0/XI0_30/d__13_ XI11_2/XI0/XI0_30/d_13_ DECAP_INV_G11
XG11674 XI11_2/XI0/XI0_30/d__12_ XI11_2/XI0/XI0_30/d_12_ DECAP_INV_G11
XG11675 XI11_2/XI0/XI0_30/d__11_ XI11_2/XI0/XI0_30/d_11_ DECAP_INV_G11
XG11676 XI11_2/XI0/XI0_30/d__10_ XI11_2/XI0/XI0_30/d_10_ DECAP_INV_G11
XG11677 XI11_2/XI0/XI0_30/d__9_ XI11_2/XI0/XI0_30/d_9_ DECAP_INV_G11
XG11678 XI11_2/XI0/XI0_30/d__8_ XI11_2/XI0/XI0_30/d_8_ DECAP_INV_G11
XG11679 XI11_2/XI0/XI0_30/d__7_ XI11_2/XI0/XI0_30/d_7_ DECAP_INV_G11
XG11680 XI11_2/XI0/XI0_30/d__6_ XI11_2/XI0/XI0_30/d_6_ DECAP_INV_G11
XG11681 XI11_2/XI0/XI0_30/d__5_ XI11_2/XI0/XI0_30/d_5_ DECAP_INV_G11
XG11682 XI11_2/XI0/XI0_30/d__4_ XI11_2/XI0/XI0_30/d_4_ DECAP_INV_G11
XG11683 XI11_2/XI0/XI0_30/d__3_ XI11_2/XI0/XI0_30/d_3_ DECAP_INV_G11
XG11684 XI11_2/XI0/XI0_30/d__2_ XI11_2/XI0/XI0_30/d_2_ DECAP_INV_G11
XG11685 XI11_2/XI0/XI0_30/d__1_ XI11_2/XI0/XI0_30/d_1_ DECAP_INV_G11
XG11686 XI11_2/XI0/XI0_30/d__0_ XI11_2/XI0/XI0_30/d_0_ DECAP_INV_G11
XG11687 XI11_2/XI0/XI0_30/d_15_ XI11_2/XI0/XI0_30/d__15_ DECAP_INV_G11
XG11688 XI11_2/XI0/XI0_30/d_14_ XI11_2/XI0/XI0_30/d__14_ DECAP_INV_G11
XG11689 XI11_2/XI0/XI0_30/d_13_ XI11_2/XI0/XI0_30/d__13_ DECAP_INV_G11
XG11690 XI11_2/XI0/XI0_30/d_12_ XI11_2/XI0/XI0_30/d__12_ DECAP_INV_G11
XG11691 XI11_2/XI0/XI0_30/d_11_ XI11_2/XI0/XI0_30/d__11_ DECAP_INV_G11
XG11692 XI11_2/XI0/XI0_30/d_10_ XI11_2/XI0/XI0_30/d__10_ DECAP_INV_G11
XG11693 XI11_2/XI0/XI0_30/d_9_ XI11_2/XI0/XI0_30/d__9_ DECAP_INV_G11
XG11694 XI11_2/XI0/XI0_30/d_8_ XI11_2/XI0/XI0_30/d__8_ DECAP_INV_G11
XG11695 XI11_2/XI0/XI0_30/d_7_ XI11_2/XI0/XI0_30/d__7_ DECAP_INV_G11
XG11696 XI11_2/XI0/XI0_30/d_6_ XI11_2/XI0/XI0_30/d__6_ DECAP_INV_G11
XG11697 XI11_2/XI0/XI0_30/d_5_ XI11_2/XI0/XI0_30/d__5_ DECAP_INV_G11
XG11698 XI11_2/XI0/XI0_30/d_4_ XI11_2/XI0/XI0_30/d__4_ DECAP_INV_G11
XG11699 XI11_2/XI0/XI0_30/d_3_ XI11_2/XI0/XI0_30/d__3_ DECAP_INV_G11
XG11700 XI11_2/XI0/XI0_30/d_2_ XI11_2/XI0/XI0_30/d__2_ DECAP_INV_G11
XG11701 XI11_2/XI0/XI0_30/d_1_ XI11_2/XI0/XI0_30/d__1_ DECAP_INV_G11
XG11702 XI11_2/XI0/XI0_30/d_0_ XI11_2/XI0/XI0_30/d__0_ DECAP_INV_G11
XG11703 XI11_2/XI0/XI0_29/d__15_ XI11_2/XI0/XI0_29/d_15_ DECAP_INV_G11
XG11704 XI11_2/XI0/XI0_29/d__14_ XI11_2/XI0/XI0_29/d_14_ DECAP_INV_G11
XG11705 XI11_2/XI0/XI0_29/d__13_ XI11_2/XI0/XI0_29/d_13_ DECAP_INV_G11
XG11706 XI11_2/XI0/XI0_29/d__12_ XI11_2/XI0/XI0_29/d_12_ DECAP_INV_G11
XG11707 XI11_2/XI0/XI0_29/d__11_ XI11_2/XI0/XI0_29/d_11_ DECAP_INV_G11
XG11708 XI11_2/XI0/XI0_29/d__10_ XI11_2/XI0/XI0_29/d_10_ DECAP_INV_G11
XG11709 XI11_2/XI0/XI0_29/d__9_ XI11_2/XI0/XI0_29/d_9_ DECAP_INV_G11
XG11710 XI11_2/XI0/XI0_29/d__8_ XI11_2/XI0/XI0_29/d_8_ DECAP_INV_G11
XG11711 XI11_2/XI0/XI0_29/d__7_ XI11_2/XI0/XI0_29/d_7_ DECAP_INV_G11
XG11712 XI11_2/XI0/XI0_29/d__6_ XI11_2/XI0/XI0_29/d_6_ DECAP_INV_G11
XG11713 XI11_2/XI0/XI0_29/d__5_ XI11_2/XI0/XI0_29/d_5_ DECAP_INV_G11
XG11714 XI11_2/XI0/XI0_29/d__4_ XI11_2/XI0/XI0_29/d_4_ DECAP_INV_G11
XG11715 XI11_2/XI0/XI0_29/d__3_ XI11_2/XI0/XI0_29/d_3_ DECAP_INV_G11
XG11716 XI11_2/XI0/XI0_29/d__2_ XI11_2/XI0/XI0_29/d_2_ DECAP_INV_G11
XG11717 XI11_2/XI0/XI0_29/d__1_ XI11_2/XI0/XI0_29/d_1_ DECAP_INV_G11
XG11718 XI11_2/XI0/XI0_29/d__0_ XI11_2/XI0/XI0_29/d_0_ DECAP_INV_G11
XG11719 XI11_2/XI0/XI0_29/d_15_ XI11_2/XI0/XI0_29/d__15_ DECAP_INV_G11
XG11720 XI11_2/XI0/XI0_29/d_14_ XI11_2/XI0/XI0_29/d__14_ DECAP_INV_G11
XG11721 XI11_2/XI0/XI0_29/d_13_ XI11_2/XI0/XI0_29/d__13_ DECAP_INV_G11
XG11722 XI11_2/XI0/XI0_29/d_12_ XI11_2/XI0/XI0_29/d__12_ DECAP_INV_G11
XG11723 XI11_2/XI0/XI0_29/d_11_ XI11_2/XI0/XI0_29/d__11_ DECAP_INV_G11
XG11724 XI11_2/XI0/XI0_29/d_10_ XI11_2/XI0/XI0_29/d__10_ DECAP_INV_G11
XG11725 XI11_2/XI0/XI0_29/d_9_ XI11_2/XI0/XI0_29/d__9_ DECAP_INV_G11
XG11726 XI11_2/XI0/XI0_29/d_8_ XI11_2/XI0/XI0_29/d__8_ DECAP_INV_G11
XG11727 XI11_2/XI0/XI0_29/d_7_ XI11_2/XI0/XI0_29/d__7_ DECAP_INV_G11
XG11728 XI11_2/XI0/XI0_29/d_6_ XI11_2/XI0/XI0_29/d__6_ DECAP_INV_G11
XG11729 XI11_2/XI0/XI0_29/d_5_ XI11_2/XI0/XI0_29/d__5_ DECAP_INV_G11
XG11730 XI11_2/XI0/XI0_29/d_4_ XI11_2/XI0/XI0_29/d__4_ DECAP_INV_G11
XG11731 XI11_2/XI0/XI0_29/d_3_ XI11_2/XI0/XI0_29/d__3_ DECAP_INV_G11
XG11732 XI11_2/XI0/XI0_29/d_2_ XI11_2/XI0/XI0_29/d__2_ DECAP_INV_G11
XG11733 XI11_2/XI0/XI0_29/d_1_ XI11_2/XI0/XI0_29/d__1_ DECAP_INV_G11
XG11734 XI11_2/XI0/XI0_29/d_0_ XI11_2/XI0/XI0_29/d__0_ DECAP_INV_G11
XG11735 XI11_2/XI0/XI0_28/d__15_ XI11_2/XI0/XI0_28/d_15_ DECAP_INV_G11
XG11736 XI11_2/XI0/XI0_28/d__14_ XI11_2/XI0/XI0_28/d_14_ DECAP_INV_G11
XG11737 XI11_2/XI0/XI0_28/d__13_ XI11_2/XI0/XI0_28/d_13_ DECAP_INV_G11
XG11738 XI11_2/XI0/XI0_28/d__12_ XI11_2/XI0/XI0_28/d_12_ DECAP_INV_G11
XG11739 XI11_2/XI0/XI0_28/d__11_ XI11_2/XI0/XI0_28/d_11_ DECAP_INV_G11
XG11740 XI11_2/XI0/XI0_28/d__10_ XI11_2/XI0/XI0_28/d_10_ DECAP_INV_G11
XG11741 XI11_2/XI0/XI0_28/d__9_ XI11_2/XI0/XI0_28/d_9_ DECAP_INV_G11
XG11742 XI11_2/XI0/XI0_28/d__8_ XI11_2/XI0/XI0_28/d_8_ DECAP_INV_G11
XG11743 XI11_2/XI0/XI0_28/d__7_ XI11_2/XI0/XI0_28/d_7_ DECAP_INV_G11
XG11744 XI11_2/XI0/XI0_28/d__6_ XI11_2/XI0/XI0_28/d_6_ DECAP_INV_G11
XG11745 XI11_2/XI0/XI0_28/d__5_ XI11_2/XI0/XI0_28/d_5_ DECAP_INV_G11
XG11746 XI11_2/XI0/XI0_28/d__4_ XI11_2/XI0/XI0_28/d_4_ DECAP_INV_G11
XG11747 XI11_2/XI0/XI0_28/d__3_ XI11_2/XI0/XI0_28/d_3_ DECAP_INV_G11
XG11748 XI11_2/XI0/XI0_28/d__2_ XI11_2/XI0/XI0_28/d_2_ DECAP_INV_G11
XG11749 XI11_2/XI0/XI0_28/d__1_ XI11_2/XI0/XI0_28/d_1_ DECAP_INV_G11
XG11750 XI11_2/XI0/XI0_28/d__0_ XI11_2/XI0/XI0_28/d_0_ DECAP_INV_G11
XG11751 XI11_2/XI0/XI0_28/d_15_ XI11_2/XI0/XI0_28/d__15_ DECAP_INV_G11
XG11752 XI11_2/XI0/XI0_28/d_14_ XI11_2/XI0/XI0_28/d__14_ DECAP_INV_G11
XG11753 XI11_2/XI0/XI0_28/d_13_ XI11_2/XI0/XI0_28/d__13_ DECAP_INV_G11
XG11754 XI11_2/XI0/XI0_28/d_12_ XI11_2/XI0/XI0_28/d__12_ DECAP_INV_G11
XG11755 XI11_2/XI0/XI0_28/d_11_ XI11_2/XI0/XI0_28/d__11_ DECAP_INV_G11
XG11756 XI11_2/XI0/XI0_28/d_10_ XI11_2/XI0/XI0_28/d__10_ DECAP_INV_G11
XG11757 XI11_2/XI0/XI0_28/d_9_ XI11_2/XI0/XI0_28/d__9_ DECAP_INV_G11
XG11758 XI11_2/XI0/XI0_28/d_8_ XI11_2/XI0/XI0_28/d__8_ DECAP_INV_G11
XG11759 XI11_2/XI0/XI0_28/d_7_ XI11_2/XI0/XI0_28/d__7_ DECAP_INV_G11
XG11760 XI11_2/XI0/XI0_28/d_6_ XI11_2/XI0/XI0_28/d__6_ DECAP_INV_G11
XG11761 XI11_2/XI0/XI0_28/d_5_ XI11_2/XI0/XI0_28/d__5_ DECAP_INV_G11
XG11762 XI11_2/XI0/XI0_28/d_4_ XI11_2/XI0/XI0_28/d__4_ DECAP_INV_G11
XG11763 XI11_2/XI0/XI0_28/d_3_ XI11_2/XI0/XI0_28/d__3_ DECAP_INV_G11
XG11764 XI11_2/XI0/XI0_28/d_2_ XI11_2/XI0/XI0_28/d__2_ DECAP_INV_G11
XG11765 XI11_2/XI0/XI0_28/d_1_ XI11_2/XI0/XI0_28/d__1_ DECAP_INV_G11
XG11766 XI11_2/XI0/XI0_28/d_0_ XI11_2/XI0/XI0_28/d__0_ DECAP_INV_G11
XG11767 XI11_2/XI0/XI0_27/d__15_ XI11_2/XI0/XI0_27/d_15_ DECAP_INV_G11
XG11768 XI11_2/XI0/XI0_27/d__14_ XI11_2/XI0/XI0_27/d_14_ DECAP_INV_G11
XG11769 XI11_2/XI0/XI0_27/d__13_ XI11_2/XI0/XI0_27/d_13_ DECAP_INV_G11
XG11770 XI11_2/XI0/XI0_27/d__12_ XI11_2/XI0/XI0_27/d_12_ DECAP_INV_G11
XG11771 XI11_2/XI0/XI0_27/d__11_ XI11_2/XI0/XI0_27/d_11_ DECAP_INV_G11
XG11772 XI11_2/XI0/XI0_27/d__10_ XI11_2/XI0/XI0_27/d_10_ DECAP_INV_G11
XG11773 XI11_2/XI0/XI0_27/d__9_ XI11_2/XI0/XI0_27/d_9_ DECAP_INV_G11
XG11774 XI11_2/XI0/XI0_27/d__8_ XI11_2/XI0/XI0_27/d_8_ DECAP_INV_G11
XG11775 XI11_2/XI0/XI0_27/d__7_ XI11_2/XI0/XI0_27/d_7_ DECAP_INV_G11
XG11776 XI11_2/XI0/XI0_27/d__6_ XI11_2/XI0/XI0_27/d_6_ DECAP_INV_G11
XG11777 XI11_2/XI0/XI0_27/d__5_ XI11_2/XI0/XI0_27/d_5_ DECAP_INV_G11
XG11778 XI11_2/XI0/XI0_27/d__4_ XI11_2/XI0/XI0_27/d_4_ DECAP_INV_G11
XG11779 XI11_2/XI0/XI0_27/d__3_ XI11_2/XI0/XI0_27/d_3_ DECAP_INV_G11
XG11780 XI11_2/XI0/XI0_27/d__2_ XI11_2/XI0/XI0_27/d_2_ DECAP_INV_G11
XG11781 XI11_2/XI0/XI0_27/d__1_ XI11_2/XI0/XI0_27/d_1_ DECAP_INV_G11
XG11782 XI11_2/XI0/XI0_27/d__0_ XI11_2/XI0/XI0_27/d_0_ DECAP_INV_G11
XG11783 XI11_2/XI0/XI0_27/d_15_ XI11_2/XI0/XI0_27/d__15_ DECAP_INV_G11
XG11784 XI11_2/XI0/XI0_27/d_14_ XI11_2/XI0/XI0_27/d__14_ DECAP_INV_G11
XG11785 XI11_2/XI0/XI0_27/d_13_ XI11_2/XI0/XI0_27/d__13_ DECAP_INV_G11
XG11786 XI11_2/XI0/XI0_27/d_12_ XI11_2/XI0/XI0_27/d__12_ DECAP_INV_G11
XG11787 XI11_2/XI0/XI0_27/d_11_ XI11_2/XI0/XI0_27/d__11_ DECAP_INV_G11
XG11788 XI11_2/XI0/XI0_27/d_10_ XI11_2/XI0/XI0_27/d__10_ DECAP_INV_G11
XG11789 XI11_2/XI0/XI0_27/d_9_ XI11_2/XI0/XI0_27/d__9_ DECAP_INV_G11
XG11790 XI11_2/XI0/XI0_27/d_8_ XI11_2/XI0/XI0_27/d__8_ DECAP_INV_G11
XG11791 XI11_2/XI0/XI0_27/d_7_ XI11_2/XI0/XI0_27/d__7_ DECAP_INV_G11
XG11792 XI11_2/XI0/XI0_27/d_6_ XI11_2/XI0/XI0_27/d__6_ DECAP_INV_G11
XG11793 XI11_2/XI0/XI0_27/d_5_ XI11_2/XI0/XI0_27/d__5_ DECAP_INV_G11
XG11794 XI11_2/XI0/XI0_27/d_4_ XI11_2/XI0/XI0_27/d__4_ DECAP_INV_G11
XG11795 XI11_2/XI0/XI0_27/d_3_ XI11_2/XI0/XI0_27/d__3_ DECAP_INV_G11
XG11796 XI11_2/XI0/XI0_27/d_2_ XI11_2/XI0/XI0_27/d__2_ DECAP_INV_G11
XG11797 XI11_2/XI0/XI0_27/d_1_ XI11_2/XI0/XI0_27/d__1_ DECAP_INV_G11
XG11798 XI11_2/XI0/XI0_27/d_0_ XI11_2/XI0/XI0_27/d__0_ DECAP_INV_G11
XG11799 XI11_2/XI0/XI0_26/d__15_ XI11_2/XI0/XI0_26/d_15_ DECAP_INV_G11
XG11800 XI11_2/XI0/XI0_26/d__14_ XI11_2/XI0/XI0_26/d_14_ DECAP_INV_G11
XG11801 XI11_2/XI0/XI0_26/d__13_ XI11_2/XI0/XI0_26/d_13_ DECAP_INV_G11
XG11802 XI11_2/XI0/XI0_26/d__12_ XI11_2/XI0/XI0_26/d_12_ DECAP_INV_G11
XG11803 XI11_2/XI0/XI0_26/d__11_ XI11_2/XI0/XI0_26/d_11_ DECAP_INV_G11
XG11804 XI11_2/XI0/XI0_26/d__10_ XI11_2/XI0/XI0_26/d_10_ DECAP_INV_G11
XG11805 XI11_2/XI0/XI0_26/d__9_ XI11_2/XI0/XI0_26/d_9_ DECAP_INV_G11
XG11806 XI11_2/XI0/XI0_26/d__8_ XI11_2/XI0/XI0_26/d_8_ DECAP_INV_G11
XG11807 XI11_2/XI0/XI0_26/d__7_ XI11_2/XI0/XI0_26/d_7_ DECAP_INV_G11
XG11808 XI11_2/XI0/XI0_26/d__6_ XI11_2/XI0/XI0_26/d_6_ DECAP_INV_G11
XG11809 XI11_2/XI0/XI0_26/d__5_ XI11_2/XI0/XI0_26/d_5_ DECAP_INV_G11
XG11810 XI11_2/XI0/XI0_26/d__4_ XI11_2/XI0/XI0_26/d_4_ DECAP_INV_G11
XG11811 XI11_2/XI0/XI0_26/d__3_ XI11_2/XI0/XI0_26/d_3_ DECAP_INV_G11
XG11812 XI11_2/XI0/XI0_26/d__2_ XI11_2/XI0/XI0_26/d_2_ DECAP_INV_G11
XG11813 XI11_2/XI0/XI0_26/d__1_ XI11_2/XI0/XI0_26/d_1_ DECAP_INV_G11
XG11814 XI11_2/XI0/XI0_26/d__0_ XI11_2/XI0/XI0_26/d_0_ DECAP_INV_G11
XG11815 XI11_2/XI0/XI0_26/d_15_ XI11_2/XI0/XI0_26/d__15_ DECAP_INV_G11
XG11816 XI11_2/XI0/XI0_26/d_14_ XI11_2/XI0/XI0_26/d__14_ DECAP_INV_G11
XG11817 XI11_2/XI0/XI0_26/d_13_ XI11_2/XI0/XI0_26/d__13_ DECAP_INV_G11
XG11818 XI11_2/XI0/XI0_26/d_12_ XI11_2/XI0/XI0_26/d__12_ DECAP_INV_G11
XG11819 XI11_2/XI0/XI0_26/d_11_ XI11_2/XI0/XI0_26/d__11_ DECAP_INV_G11
XG11820 XI11_2/XI0/XI0_26/d_10_ XI11_2/XI0/XI0_26/d__10_ DECAP_INV_G11
XG11821 XI11_2/XI0/XI0_26/d_9_ XI11_2/XI0/XI0_26/d__9_ DECAP_INV_G11
XG11822 XI11_2/XI0/XI0_26/d_8_ XI11_2/XI0/XI0_26/d__8_ DECAP_INV_G11
XG11823 XI11_2/XI0/XI0_26/d_7_ XI11_2/XI0/XI0_26/d__7_ DECAP_INV_G11
XG11824 XI11_2/XI0/XI0_26/d_6_ XI11_2/XI0/XI0_26/d__6_ DECAP_INV_G11
XG11825 XI11_2/XI0/XI0_26/d_5_ XI11_2/XI0/XI0_26/d__5_ DECAP_INV_G11
XG11826 XI11_2/XI0/XI0_26/d_4_ XI11_2/XI0/XI0_26/d__4_ DECAP_INV_G11
XG11827 XI11_2/XI0/XI0_26/d_3_ XI11_2/XI0/XI0_26/d__3_ DECAP_INV_G11
XG11828 XI11_2/XI0/XI0_26/d_2_ XI11_2/XI0/XI0_26/d__2_ DECAP_INV_G11
XG11829 XI11_2/XI0/XI0_26/d_1_ XI11_2/XI0/XI0_26/d__1_ DECAP_INV_G11
XG11830 XI11_2/XI0/XI0_26/d_0_ XI11_2/XI0/XI0_26/d__0_ DECAP_INV_G11
XG11831 XI11_2/XI0/XI0_25/d__15_ XI11_2/XI0/XI0_25/d_15_ DECAP_INV_G11
XG11832 XI11_2/XI0/XI0_25/d__14_ XI11_2/XI0/XI0_25/d_14_ DECAP_INV_G11
XG11833 XI11_2/XI0/XI0_25/d__13_ XI11_2/XI0/XI0_25/d_13_ DECAP_INV_G11
XG11834 XI11_2/XI0/XI0_25/d__12_ XI11_2/XI0/XI0_25/d_12_ DECAP_INV_G11
XG11835 XI11_2/XI0/XI0_25/d__11_ XI11_2/XI0/XI0_25/d_11_ DECAP_INV_G11
XG11836 XI11_2/XI0/XI0_25/d__10_ XI11_2/XI0/XI0_25/d_10_ DECAP_INV_G11
XG11837 XI11_2/XI0/XI0_25/d__9_ XI11_2/XI0/XI0_25/d_9_ DECAP_INV_G11
XG11838 XI11_2/XI0/XI0_25/d__8_ XI11_2/XI0/XI0_25/d_8_ DECAP_INV_G11
XG11839 XI11_2/XI0/XI0_25/d__7_ XI11_2/XI0/XI0_25/d_7_ DECAP_INV_G11
XG11840 XI11_2/XI0/XI0_25/d__6_ XI11_2/XI0/XI0_25/d_6_ DECAP_INV_G11
XG11841 XI11_2/XI0/XI0_25/d__5_ XI11_2/XI0/XI0_25/d_5_ DECAP_INV_G11
XG11842 XI11_2/XI0/XI0_25/d__4_ XI11_2/XI0/XI0_25/d_4_ DECAP_INV_G11
XG11843 XI11_2/XI0/XI0_25/d__3_ XI11_2/XI0/XI0_25/d_3_ DECAP_INV_G11
XG11844 XI11_2/XI0/XI0_25/d__2_ XI11_2/XI0/XI0_25/d_2_ DECAP_INV_G11
XG11845 XI11_2/XI0/XI0_25/d__1_ XI11_2/XI0/XI0_25/d_1_ DECAP_INV_G11
XG11846 XI11_2/XI0/XI0_25/d__0_ XI11_2/XI0/XI0_25/d_0_ DECAP_INV_G11
XG11847 XI11_2/XI0/XI0_25/d_15_ XI11_2/XI0/XI0_25/d__15_ DECAP_INV_G11
XG11848 XI11_2/XI0/XI0_25/d_14_ XI11_2/XI0/XI0_25/d__14_ DECAP_INV_G11
XG11849 XI11_2/XI0/XI0_25/d_13_ XI11_2/XI0/XI0_25/d__13_ DECAP_INV_G11
XG11850 XI11_2/XI0/XI0_25/d_12_ XI11_2/XI0/XI0_25/d__12_ DECAP_INV_G11
XG11851 XI11_2/XI0/XI0_25/d_11_ XI11_2/XI0/XI0_25/d__11_ DECAP_INV_G11
XG11852 XI11_2/XI0/XI0_25/d_10_ XI11_2/XI0/XI0_25/d__10_ DECAP_INV_G11
XG11853 XI11_2/XI0/XI0_25/d_9_ XI11_2/XI0/XI0_25/d__9_ DECAP_INV_G11
XG11854 XI11_2/XI0/XI0_25/d_8_ XI11_2/XI0/XI0_25/d__8_ DECAP_INV_G11
XG11855 XI11_2/XI0/XI0_25/d_7_ XI11_2/XI0/XI0_25/d__7_ DECAP_INV_G11
XG11856 XI11_2/XI0/XI0_25/d_6_ XI11_2/XI0/XI0_25/d__6_ DECAP_INV_G11
XG11857 XI11_2/XI0/XI0_25/d_5_ XI11_2/XI0/XI0_25/d__5_ DECAP_INV_G11
XG11858 XI11_2/XI0/XI0_25/d_4_ XI11_2/XI0/XI0_25/d__4_ DECAP_INV_G11
XG11859 XI11_2/XI0/XI0_25/d_3_ XI11_2/XI0/XI0_25/d__3_ DECAP_INV_G11
XG11860 XI11_2/XI0/XI0_25/d_2_ XI11_2/XI0/XI0_25/d__2_ DECAP_INV_G11
XG11861 XI11_2/XI0/XI0_25/d_1_ XI11_2/XI0/XI0_25/d__1_ DECAP_INV_G11
XG11862 XI11_2/XI0/XI0_25/d_0_ XI11_2/XI0/XI0_25/d__0_ DECAP_INV_G11
XG11863 XI11_2/XI0/XI0_24/d__15_ XI11_2/XI0/XI0_24/d_15_ DECAP_INV_G11
XG11864 XI11_2/XI0/XI0_24/d__14_ XI11_2/XI0/XI0_24/d_14_ DECAP_INV_G11
XG11865 XI11_2/XI0/XI0_24/d__13_ XI11_2/XI0/XI0_24/d_13_ DECAP_INV_G11
XG11866 XI11_2/XI0/XI0_24/d__12_ XI11_2/XI0/XI0_24/d_12_ DECAP_INV_G11
XG11867 XI11_2/XI0/XI0_24/d__11_ XI11_2/XI0/XI0_24/d_11_ DECAP_INV_G11
XG11868 XI11_2/XI0/XI0_24/d__10_ XI11_2/XI0/XI0_24/d_10_ DECAP_INV_G11
XG11869 XI11_2/XI0/XI0_24/d__9_ XI11_2/XI0/XI0_24/d_9_ DECAP_INV_G11
XG11870 XI11_2/XI0/XI0_24/d__8_ XI11_2/XI0/XI0_24/d_8_ DECAP_INV_G11
XG11871 XI11_2/XI0/XI0_24/d__7_ XI11_2/XI0/XI0_24/d_7_ DECAP_INV_G11
XG11872 XI11_2/XI0/XI0_24/d__6_ XI11_2/XI0/XI0_24/d_6_ DECAP_INV_G11
XG11873 XI11_2/XI0/XI0_24/d__5_ XI11_2/XI0/XI0_24/d_5_ DECAP_INV_G11
XG11874 XI11_2/XI0/XI0_24/d__4_ XI11_2/XI0/XI0_24/d_4_ DECAP_INV_G11
XG11875 XI11_2/XI0/XI0_24/d__3_ XI11_2/XI0/XI0_24/d_3_ DECAP_INV_G11
XG11876 XI11_2/XI0/XI0_24/d__2_ XI11_2/XI0/XI0_24/d_2_ DECAP_INV_G11
XG11877 XI11_2/XI0/XI0_24/d__1_ XI11_2/XI0/XI0_24/d_1_ DECAP_INV_G11
XG11878 XI11_2/XI0/XI0_24/d__0_ XI11_2/XI0/XI0_24/d_0_ DECAP_INV_G11
XG11879 XI11_2/XI0/XI0_24/d_15_ XI11_2/XI0/XI0_24/d__15_ DECAP_INV_G11
XG11880 XI11_2/XI0/XI0_24/d_14_ XI11_2/XI0/XI0_24/d__14_ DECAP_INV_G11
XG11881 XI11_2/XI0/XI0_24/d_13_ XI11_2/XI0/XI0_24/d__13_ DECAP_INV_G11
XG11882 XI11_2/XI0/XI0_24/d_12_ XI11_2/XI0/XI0_24/d__12_ DECAP_INV_G11
XG11883 XI11_2/XI0/XI0_24/d_11_ XI11_2/XI0/XI0_24/d__11_ DECAP_INV_G11
XG11884 XI11_2/XI0/XI0_24/d_10_ XI11_2/XI0/XI0_24/d__10_ DECAP_INV_G11
XG11885 XI11_2/XI0/XI0_24/d_9_ XI11_2/XI0/XI0_24/d__9_ DECAP_INV_G11
XG11886 XI11_2/XI0/XI0_24/d_8_ XI11_2/XI0/XI0_24/d__8_ DECAP_INV_G11
XG11887 XI11_2/XI0/XI0_24/d_7_ XI11_2/XI0/XI0_24/d__7_ DECAP_INV_G11
XG11888 XI11_2/XI0/XI0_24/d_6_ XI11_2/XI0/XI0_24/d__6_ DECAP_INV_G11
XG11889 XI11_2/XI0/XI0_24/d_5_ XI11_2/XI0/XI0_24/d__5_ DECAP_INV_G11
XG11890 XI11_2/XI0/XI0_24/d_4_ XI11_2/XI0/XI0_24/d__4_ DECAP_INV_G11
XG11891 XI11_2/XI0/XI0_24/d_3_ XI11_2/XI0/XI0_24/d__3_ DECAP_INV_G11
XG11892 XI11_2/XI0/XI0_24/d_2_ XI11_2/XI0/XI0_24/d__2_ DECAP_INV_G11
XG11893 XI11_2/XI0/XI0_24/d_1_ XI11_2/XI0/XI0_24/d__1_ DECAP_INV_G11
XG11894 XI11_2/XI0/XI0_24/d_0_ XI11_2/XI0/XI0_24/d__0_ DECAP_INV_G11
XG11895 XI11_2/XI0/XI0_23/d__15_ XI11_2/XI0/XI0_23/d_15_ DECAP_INV_G11
XG11896 XI11_2/XI0/XI0_23/d__14_ XI11_2/XI0/XI0_23/d_14_ DECAP_INV_G11
XG11897 XI11_2/XI0/XI0_23/d__13_ XI11_2/XI0/XI0_23/d_13_ DECAP_INV_G11
XG11898 XI11_2/XI0/XI0_23/d__12_ XI11_2/XI0/XI0_23/d_12_ DECAP_INV_G11
XG11899 XI11_2/XI0/XI0_23/d__11_ XI11_2/XI0/XI0_23/d_11_ DECAP_INV_G11
XG11900 XI11_2/XI0/XI0_23/d__10_ XI11_2/XI0/XI0_23/d_10_ DECAP_INV_G11
XG11901 XI11_2/XI0/XI0_23/d__9_ XI11_2/XI0/XI0_23/d_9_ DECAP_INV_G11
XG11902 XI11_2/XI0/XI0_23/d__8_ XI11_2/XI0/XI0_23/d_8_ DECAP_INV_G11
XG11903 XI11_2/XI0/XI0_23/d__7_ XI11_2/XI0/XI0_23/d_7_ DECAP_INV_G11
XG11904 XI11_2/XI0/XI0_23/d__6_ XI11_2/XI0/XI0_23/d_6_ DECAP_INV_G11
XG11905 XI11_2/XI0/XI0_23/d__5_ XI11_2/XI0/XI0_23/d_5_ DECAP_INV_G11
XG11906 XI11_2/XI0/XI0_23/d__4_ XI11_2/XI0/XI0_23/d_4_ DECAP_INV_G11
XG11907 XI11_2/XI0/XI0_23/d__3_ XI11_2/XI0/XI0_23/d_3_ DECAP_INV_G11
XG11908 XI11_2/XI0/XI0_23/d__2_ XI11_2/XI0/XI0_23/d_2_ DECAP_INV_G11
XG11909 XI11_2/XI0/XI0_23/d__1_ XI11_2/XI0/XI0_23/d_1_ DECAP_INV_G11
XG11910 XI11_2/XI0/XI0_23/d__0_ XI11_2/XI0/XI0_23/d_0_ DECAP_INV_G11
XG11911 XI11_2/XI0/XI0_23/d_15_ XI11_2/XI0/XI0_23/d__15_ DECAP_INV_G11
XG11912 XI11_2/XI0/XI0_23/d_14_ XI11_2/XI0/XI0_23/d__14_ DECAP_INV_G11
XG11913 XI11_2/XI0/XI0_23/d_13_ XI11_2/XI0/XI0_23/d__13_ DECAP_INV_G11
XG11914 XI11_2/XI0/XI0_23/d_12_ XI11_2/XI0/XI0_23/d__12_ DECAP_INV_G11
XG11915 XI11_2/XI0/XI0_23/d_11_ XI11_2/XI0/XI0_23/d__11_ DECAP_INV_G11
XG11916 XI11_2/XI0/XI0_23/d_10_ XI11_2/XI0/XI0_23/d__10_ DECAP_INV_G11
XG11917 XI11_2/XI0/XI0_23/d_9_ XI11_2/XI0/XI0_23/d__9_ DECAP_INV_G11
XG11918 XI11_2/XI0/XI0_23/d_8_ XI11_2/XI0/XI0_23/d__8_ DECAP_INV_G11
XG11919 XI11_2/XI0/XI0_23/d_7_ XI11_2/XI0/XI0_23/d__7_ DECAP_INV_G11
XG11920 XI11_2/XI0/XI0_23/d_6_ XI11_2/XI0/XI0_23/d__6_ DECAP_INV_G11
XG11921 XI11_2/XI0/XI0_23/d_5_ XI11_2/XI0/XI0_23/d__5_ DECAP_INV_G11
XG11922 XI11_2/XI0/XI0_23/d_4_ XI11_2/XI0/XI0_23/d__4_ DECAP_INV_G11
XG11923 XI11_2/XI0/XI0_23/d_3_ XI11_2/XI0/XI0_23/d__3_ DECAP_INV_G11
XG11924 XI11_2/XI0/XI0_23/d_2_ XI11_2/XI0/XI0_23/d__2_ DECAP_INV_G11
XG11925 XI11_2/XI0/XI0_23/d_1_ XI11_2/XI0/XI0_23/d__1_ DECAP_INV_G11
XG11926 XI11_2/XI0/XI0_23/d_0_ XI11_2/XI0/XI0_23/d__0_ DECAP_INV_G11
XG11927 XI11_2/XI0/XI0_22/d__15_ XI11_2/XI0/XI0_22/d_15_ DECAP_INV_G11
XG11928 XI11_2/XI0/XI0_22/d__14_ XI11_2/XI0/XI0_22/d_14_ DECAP_INV_G11
XG11929 XI11_2/XI0/XI0_22/d__13_ XI11_2/XI0/XI0_22/d_13_ DECAP_INV_G11
XG11930 XI11_2/XI0/XI0_22/d__12_ XI11_2/XI0/XI0_22/d_12_ DECAP_INV_G11
XG11931 XI11_2/XI0/XI0_22/d__11_ XI11_2/XI0/XI0_22/d_11_ DECAP_INV_G11
XG11932 XI11_2/XI0/XI0_22/d__10_ XI11_2/XI0/XI0_22/d_10_ DECAP_INV_G11
XG11933 XI11_2/XI0/XI0_22/d__9_ XI11_2/XI0/XI0_22/d_9_ DECAP_INV_G11
XG11934 XI11_2/XI0/XI0_22/d__8_ XI11_2/XI0/XI0_22/d_8_ DECAP_INV_G11
XG11935 XI11_2/XI0/XI0_22/d__7_ XI11_2/XI0/XI0_22/d_7_ DECAP_INV_G11
XG11936 XI11_2/XI0/XI0_22/d__6_ XI11_2/XI0/XI0_22/d_6_ DECAP_INV_G11
XG11937 XI11_2/XI0/XI0_22/d__5_ XI11_2/XI0/XI0_22/d_5_ DECAP_INV_G11
XG11938 XI11_2/XI0/XI0_22/d__4_ XI11_2/XI0/XI0_22/d_4_ DECAP_INV_G11
XG11939 XI11_2/XI0/XI0_22/d__3_ XI11_2/XI0/XI0_22/d_3_ DECAP_INV_G11
XG11940 XI11_2/XI0/XI0_22/d__2_ XI11_2/XI0/XI0_22/d_2_ DECAP_INV_G11
XG11941 XI11_2/XI0/XI0_22/d__1_ XI11_2/XI0/XI0_22/d_1_ DECAP_INV_G11
XG11942 XI11_2/XI0/XI0_22/d__0_ XI11_2/XI0/XI0_22/d_0_ DECAP_INV_G11
XG11943 XI11_2/XI0/XI0_22/d_15_ XI11_2/XI0/XI0_22/d__15_ DECAP_INV_G11
XG11944 XI11_2/XI0/XI0_22/d_14_ XI11_2/XI0/XI0_22/d__14_ DECAP_INV_G11
XG11945 XI11_2/XI0/XI0_22/d_13_ XI11_2/XI0/XI0_22/d__13_ DECAP_INV_G11
XG11946 XI11_2/XI0/XI0_22/d_12_ XI11_2/XI0/XI0_22/d__12_ DECAP_INV_G11
XG11947 XI11_2/XI0/XI0_22/d_11_ XI11_2/XI0/XI0_22/d__11_ DECAP_INV_G11
XG11948 XI11_2/XI0/XI0_22/d_10_ XI11_2/XI0/XI0_22/d__10_ DECAP_INV_G11
XG11949 XI11_2/XI0/XI0_22/d_9_ XI11_2/XI0/XI0_22/d__9_ DECAP_INV_G11
XG11950 XI11_2/XI0/XI0_22/d_8_ XI11_2/XI0/XI0_22/d__8_ DECAP_INV_G11
XG11951 XI11_2/XI0/XI0_22/d_7_ XI11_2/XI0/XI0_22/d__7_ DECAP_INV_G11
XG11952 XI11_2/XI0/XI0_22/d_6_ XI11_2/XI0/XI0_22/d__6_ DECAP_INV_G11
XG11953 XI11_2/XI0/XI0_22/d_5_ XI11_2/XI0/XI0_22/d__5_ DECAP_INV_G11
XG11954 XI11_2/XI0/XI0_22/d_4_ XI11_2/XI0/XI0_22/d__4_ DECAP_INV_G11
XG11955 XI11_2/XI0/XI0_22/d_3_ XI11_2/XI0/XI0_22/d__3_ DECAP_INV_G11
XG11956 XI11_2/XI0/XI0_22/d_2_ XI11_2/XI0/XI0_22/d__2_ DECAP_INV_G11
XG11957 XI11_2/XI0/XI0_22/d_1_ XI11_2/XI0/XI0_22/d__1_ DECAP_INV_G11
XG11958 XI11_2/XI0/XI0_22/d_0_ XI11_2/XI0/XI0_22/d__0_ DECAP_INV_G11
XG11959 XI11_2/XI0/XI0_21/d__15_ XI11_2/XI0/XI0_21/d_15_ DECAP_INV_G11
XG11960 XI11_2/XI0/XI0_21/d__14_ XI11_2/XI0/XI0_21/d_14_ DECAP_INV_G11
XG11961 XI11_2/XI0/XI0_21/d__13_ XI11_2/XI0/XI0_21/d_13_ DECAP_INV_G11
XG11962 XI11_2/XI0/XI0_21/d__12_ XI11_2/XI0/XI0_21/d_12_ DECAP_INV_G11
XG11963 XI11_2/XI0/XI0_21/d__11_ XI11_2/XI0/XI0_21/d_11_ DECAP_INV_G11
XG11964 XI11_2/XI0/XI0_21/d__10_ XI11_2/XI0/XI0_21/d_10_ DECAP_INV_G11
XG11965 XI11_2/XI0/XI0_21/d__9_ XI11_2/XI0/XI0_21/d_9_ DECAP_INV_G11
XG11966 XI11_2/XI0/XI0_21/d__8_ XI11_2/XI0/XI0_21/d_8_ DECAP_INV_G11
XG11967 XI11_2/XI0/XI0_21/d__7_ XI11_2/XI0/XI0_21/d_7_ DECAP_INV_G11
XG11968 XI11_2/XI0/XI0_21/d__6_ XI11_2/XI0/XI0_21/d_6_ DECAP_INV_G11
XG11969 XI11_2/XI0/XI0_21/d__5_ XI11_2/XI0/XI0_21/d_5_ DECAP_INV_G11
XG11970 XI11_2/XI0/XI0_21/d__4_ XI11_2/XI0/XI0_21/d_4_ DECAP_INV_G11
XG11971 XI11_2/XI0/XI0_21/d__3_ XI11_2/XI0/XI0_21/d_3_ DECAP_INV_G11
XG11972 XI11_2/XI0/XI0_21/d__2_ XI11_2/XI0/XI0_21/d_2_ DECAP_INV_G11
XG11973 XI11_2/XI0/XI0_21/d__1_ XI11_2/XI0/XI0_21/d_1_ DECAP_INV_G11
XG11974 XI11_2/XI0/XI0_21/d__0_ XI11_2/XI0/XI0_21/d_0_ DECAP_INV_G11
XG11975 XI11_2/XI0/XI0_21/d_15_ XI11_2/XI0/XI0_21/d__15_ DECAP_INV_G11
XG11976 XI11_2/XI0/XI0_21/d_14_ XI11_2/XI0/XI0_21/d__14_ DECAP_INV_G11
XG11977 XI11_2/XI0/XI0_21/d_13_ XI11_2/XI0/XI0_21/d__13_ DECAP_INV_G11
XG11978 XI11_2/XI0/XI0_21/d_12_ XI11_2/XI0/XI0_21/d__12_ DECAP_INV_G11
XG11979 XI11_2/XI0/XI0_21/d_11_ XI11_2/XI0/XI0_21/d__11_ DECAP_INV_G11
XG11980 XI11_2/XI0/XI0_21/d_10_ XI11_2/XI0/XI0_21/d__10_ DECAP_INV_G11
XG11981 XI11_2/XI0/XI0_21/d_9_ XI11_2/XI0/XI0_21/d__9_ DECAP_INV_G11
XG11982 XI11_2/XI0/XI0_21/d_8_ XI11_2/XI0/XI0_21/d__8_ DECAP_INV_G11
XG11983 XI11_2/XI0/XI0_21/d_7_ XI11_2/XI0/XI0_21/d__7_ DECAP_INV_G11
XG11984 XI11_2/XI0/XI0_21/d_6_ XI11_2/XI0/XI0_21/d__6_ DECAP_INV_G11
XG11985 XI11_2/XI0/XI0_21/d_5_ XI11_2/XI0/XI0_21/d__5_ DECAP_INV_G11
XG11986 XI11_2/XI0/XI0_21/d_4_ XI11_2/XI0/XI0_21/d__4_ DECAP_INV_G11
XG11987 XI11_2/XI0/XI0_21/d_3_ XI11_2/XI0/XI0_21/d__3_ DECAP_INV_G11
XG11988 XI11_2/XI0/XI0_21/d_2_ XI11_2/XI0/XI0_21/d__2_ DECAP_INV_G11
XG11989 XI11_2/XI0/XI0_21/d_1_ XI11_2/XI0/XI0_21/d__1_ DECAP_INV_G11
XG11990 XI11_2/XI0/XI0_21/d_0_ XI11_2/XI0/XI0_21/d__0_ DECAP_INV_G11
XG11991 XI11_2/XI0/XI0_20/d__15_ XI11_2/XI0/XI0_20/d_15_ DECAP_INV_G11
XG11992 XI11_2/XI0/XI0_20/d__14_ XI11_2/XI0/XI0_20/d_14_ DECAP_INV_G11
XG11993 XI11_2/XI0/XI0_20/d__13_ XI11_2/XI0/XI0_20/d_13_ DECAP_INV_G11
XG11994 XI11_2/XI0/XI0_20/d__12_ XI11_2/XI0/XI0_20/d_12_ DECAP_INV_G11
XG11995 XI11_2/XI0/XI0_20/d__11_ XI11_2/XI0/XI0_20/d_11_ DECAP_INV_G11
XG11996 XI11_2/XI0/XI0_20/d__10_ XI11_2/XI0/XI0_20/d_10_ DECAP_INV_G11
XG11997 XI11_2/XI0/XI0_20/d__9_ XI11_2/XI0/XI0_20/d_9_ DECAP_INV_G11
XG11998 XI11_2/XI0/XI0_20/d__8_ XI11_2/XI0/XI0_20/d_8_ DECAP_INV_G11
XG11999 XI11_2/XI0/XI0_20/d__7_ XI11_2/XI0/XI0_20/d_7_ DECAP_INV_G11
XG12000 XI11_2/XI0/XI0_20/d__6_ XI11_2/XI0/XI0_20/d_6_ DECAP_INV_G11
XG12001 XI11_2/XI0/XI0_20/d__5_ XI11_2/XI0/XI0_20/d_5_ DECAP_INV_G11
XG12002 XI11_2/XI0/XI0_20/d__4_ XI11_2/XI0/XI0_20/d_4_ DECAP_INV_G11
XG12003 XI11_2/XI0/XI0_20/d__3_ XI11_2/XI0/XI0_20/d_3_ DECAP_INV_G11
XG12004 XI11_2/XI0/XI0_20/d__2_ XI11_2/XI0/XI0_20/d_2_ DECAP_INV_G11
XG12005 XI11_2/XI0/XI0_20/d__1_ XI11_2/XI0/XI0_20/d_1_ DECAP_INV_G11
XG12006 XI11_2/XI0/XI0_20/d__0_ XI11_2/XI0/XI0_20/d_0_ DECAP_INV_G11
XG12007 XI11_2/XI0/XI0_20/d_15_ XI11_2/XI0/XI0_20/d__15_ DECAP_INV_G11
XG12008 XI11_2/XI0/XI0_20/d_14_ XI11_2/XI0/XI0_20/d__14_ DECAP_INV_G11
XG12009 XI11_2/XI0/XI0_20/d_13_ XI11_2/XI0/XI0_20/d__13_ DECAP_INV_G11
XG12010 XI11_2/XI0/XI0_20/d_12_ XI11_2/XI0/XI0_20/d__12_ DECAP_INV_G11
XG12011 XI11_2/XI0/XI0_20/d_11_ XI11_2/XI0/XI0_20/d__11_ DECAP_INV_G11
XG12012 XI11_2/XI0/XI0_20/d_10_ XI11_2/XI0/XI0_20/d__10_ DECAP_INV_G11
XG12013 XI11_2/XI0/XI0_20/d_9_ XI11_2/XI0/XI0_20/d__9_ DECAP_INV_G11
XG12014 XI11_2/XI0/XI0_20/d_8_ XI11_2/XI0/XI0_20/d__8_ DECAP_INV_G11
XG12015 XI11_2/XI0/XI0_20/d_7_ XI11_2/XI0/XI0_20/d__7_ DECAP_INV_G11
XG12016 XI11_2/XI0/XI0_20/d_6_ XI11_2/XI0/XI0_20/d__6_ DECAP_INV_G11
XG12017 XI11_2/XI0/XI0_20/d_5_ XI11_2/XI0/XI0_20/d__5_ DECAP_INV_G11
XG12018 XI11_2/XI0/XI0_20/d_4_ XI11_2/XI0/XI0_20/d__4_ DECAP_INV_G11
XG12019 XI11_2/XI0/XI0_20/d_3_ XI11_2/XI0/XI0_20/d__3_ DECAP_INV_G11
XG12020 XI11_2/XI0/XI0_20/d_2_ XI11_2/XI0/XI0_20/d__2_ DECAP_INV_G11
XG12021 XI11_2/XI0/XI0_20/d_1_ XI11_2/XI0/XI0_20/d__1_ DECAP_INV_G11
XG12022 XI11_2/XI0/XI0_20/d_0_ XI11_2/XI0/XI0_20/d__0_ DECAP_INV_G11
XG12023 XI11_2/XI0/XI0_19/d__15_ XI11_2/XI0/XI0_19/d_15_ DECAP_INV_G11
XG12024 XI11_2/XI0/XI0_19/d__14_ XI11_2/XI0/XI0_19/d_14_ DECAP_INV_G11
XG12025 XI11_2/XI0/XI0_19/d__13_ XI11_2/XI0/XI0_19/d_13_ DECAP_INV_G11
XG12026 XI11_2/XI0/XI0_19/d__12_ XI11_2/XI0/XI0_19/d_12_ DECAP_INV_G11
XG12027 XI11_2/XI0/XI0_19/d__11_ XI11_2/XI0/XI0_19/d_11_ DECAP_INV_G11
XG12028 XI11_2/XI0/XI0_19/d__10_ XI11_2/XI0/XI0_19/d_10_ DECAP_INV_G11
XG12029 XI11_2/XI0/XI0_19/d__9_ XI11_2/XI0/XI0_19/d_9_ DECAP_INV_G11
XG12030 XI11_2/XI0/XI0_19/d__8_ XI11_2/XI0/XI0_19/d_8_ DECAP_INV_G11
XG12031 XI11_2/XI0/XI0_19/d__7_ XI11_2/XI0/XI0_19/d_7_ DECAP_INV_G11
XG12032 XI11_2/XI0/XI0_19/d__6_ XI11_2/XI0/XI0_19/d_6_ DECAP_INV_G11
XG12033 XI11_2/XI0/XI0_19/d__5_ XI11_2/XI0/XI0_19/d_5_ DECAP_INV_G11
XG12034 XI11_2/XI0/XI0_19/d__4_ XI11_2/XI0/XI0_19/d_4_ DECAP_INV_G11
XG12035 XI11_2/XI0/XI0_19/d__3_ XI11_2/XI0/XI0_19/d_3_ DECAP_INV_G11
XG12036 XI11_2/XI0/XI0_19/d__2_ XI11_2/XI0/XI0_19/d_2_ DECAP_INV_G11
XG12037 XI11_2/XI0/XI0_19/d__1_ XI11_2/XI0/XI0_19/d_1_ DECAP_INV_G11
XG12038 XI11_2/XI0/XI0_19/d__0_ XI11_2/XI0/XI0_19/d_0_ DECAP_INV_G11
XG12039 XI11_2/XI0/XI0_19/d_15_ XI11_2/XI0/XI0_19/d__15_ DECAP_INV_G11
XG12040 XI11_2/XI0/XI0_19/d_14_ XI11_2/XI0/XI0_19/d__14_ DECAP_INV_G11
XG12041 XI11_2/XI0/XI0_19/d_13_ XI11_2/XI0/XI0_19/d__13_ DECAP_INV_G11
XG12042 XI11_2/XI0/XI0_19/d_12_ XI11_2/XI0/XI0_19/d__12_ DECAP_INV_G11
XG12043 XI11_2/XI0/XI0_19/d_11_ XI11_2/XI0/XI0_19/d__11_ DECAP_INV_G11
XG12044 XI11_2/XI0/XI0_19/d_10_ XI11_2/XI0/XI0_19/d__10_ DECAP_INV_G11
XG12045 XI11_2/XI0/XI0_19/d_9_ XI11_2/XI0/XI0_19/d__9_ DECAP_INV_G11
XG12046 XI11_2/XI0/XI0_19/d_8_ XI11_2/XI0/XI0_19/d__8_ DECAP_INV_G11
XG12047 XI11_2/XI0/XI0_19/d_7_ XI11_2/XI0/XI0_19/d__7_ DECAP_INV_G11
XG12048 XI11_2/XI0/XI0_19/d_6_ XI11_2/XI0/XI0_19/d__6_ DECAP_INV_G11
XG12049 XI11_2/XI0/XI0_19/d_5_ XI11_2/XI0/XI0_19/d__5_ DECAP_INV_G11
XG12050 XI11_2/XI0/XI0_19/d_4_ XI11_2/XI0/XI0_19/d__4_ DECAP_INV_G11
XG12051 XI11_2/XI0/XI0_19/d_3_ XI11_2/XI0/XI0_19/d__3_ DECAP_INV_G11
XG12052 XI11_2/XI0/XI0_19/d_2_ XI11_2/XI0/XI0_19/d__2_ DECAP_INV_G11
XG12053 XI11_2/XI0/XI0_19/d_1_ XI11_2/XI0/XI0_19/d__1_ DECAP_INV_G11
XG12054 XI11_2/XI0/XI0_19/d_0_ XI11_2/XI0/XI0_19/d__0_ DECAP_INV_G11
XG12055 XI11_2/XI0/XI0_18/d__15_ XI11_2/XI0/XI0_18/d_15_ DECAP_INV_G11
XG12056 XI11_2/XI0/XI0_18/d__14_ XI11_2/XI0/XI0_18/d_14_ DECAP_INV_G11
XG12057 XI11_2/XI0/XI0_18/d__13_ XI11_2/XI0/XI0_18/d_13_ DECAP_INV_G11
XG12058 XI11_2/XI0/XI0_18/d__12_ XI11_2/XI0/XI0_18/d_12_ DECAP_INV_G11
XG12059 XI11_2/XI0/XI0_18/d__11_ XI11_2/XI0/XI0_18/d_11_ DECAP_INV_G11
XG12060 XI11_2/XI0/XI0_18/d__10_ XI11_2/XI0/XI0_18/d_10_ DECAP_INV_G11
XG12061 XI11_2/XI0/XI0_18/d__9_ XI11_2/XI0/XI0_18/d_9_ DECAP_INV_G11
XG12062 XI11_2/XI0/XI0_18/d__8_ XI11_2/XI0/XI0_18/d_8_ DECAP_INV_G11
XG12063 XI11_2/XI0/XI0_18/d__7_ XI11_2/XI0/XI0_18/d_7_ DECAP_INV_G11
XG12064 XI11_2/XI0/XI0_18/d__6_ XI11_2/XI0/XI0_18/d_6_ DECAP_INV_G11
XG12065 XI11_2/XI0/XI0_18/d__5_ XI11_2/XI0/XI0_18/d_5_ DECAP_INV_G11
XG12066 XI11_2/XI0/XI0_18/d__4_ XI11_2/XI0/XI0_18/d_4_ DECAP_INV_G11
XG12067 XI11_2/XI0/XI0_18/d__3_ XI11_2/XI0/XI0_18/d_3_ DECAP_INV_G11
XG12068 XI11_2/XI0/XI0_18/d__2_ XI11_2/XI0/XI0_18/d_2_ DECAP_INV_G11
XG12069 XI11_2/XI0/XI0_18/d__1_ XI11_2/XI0/XI0_18/d_1_ DECAP_INV_G11
XG12070 XI11_2/XI0/XI0_18/d__0_ XI11_2/XI0/XI0_18/d_0_ DECAP_INV_G11
XG12071 XI11_2/XI0/XI0_18/d_15_ XI11_2/XI0/XI0_18/d__15_ DECAP_INV_G11
XG12072 XI11_2/XI0/XI0_18/d_14_ XI11_2/XI0/XI0_18/d__14_ DECAP_INV_G11
XG12073 XI11_2/XI0/XI0_18/d_13_ XI11_2/XI0/XI0_18/d__13_ DECAP_INV_G11
XG12074 XI11_2/XI0/XI0_18/d_12_ XI11_2/XI0/XI0_18/d__12_ DECAP_INV_G11
XG12075 XI11_2/XI0/XI0_18/d_11_ XI11_2/XI0/XI0_18/d__11_ DECAP_INV_G11
XG12076 XI11_2/XI0/XI0_18/d_10_ XI11_2/XI0/XI0_18/d__10_ DECAP_INV_G11
XG12077 XI11_2/XI0/XI0_18/d_9_ XI11_2/XI0/XI0_18/d__9_ DECAP_INV_G11
XG12078 XI11_2/XI0/XI0_18/d_8_ XI11_2/XI0/XI0_18/d__8_ DECAP_INV_G11
XG12079 XI11_2/XI0/XI0_18/d_7_ XI11_2/XI0/XI0_18/d__7_ DECAP_INV_G11
XG12080 XI11_2/XI0/XI0_18/d_6_ XI11_2/XI0/XI0_18/d__6_ DECAP_INV_G11
XG12081 XI11_2/XI0/XI0_18/d_5_ XI11_2/XI0/XI0_18/d__5_ DECAP_INV_G11
XG12082 XI11_2/XI0/XI0_18/d_4_ XI11_2/XI0/XI0_18/d__4_ DECAP_INV_G11
XG12083 XI11_2/XI0/XI0_18/d_3_ XI11_2/XI0/XI0_18/d__3_ DECAP_INV_G11
XG12084 XI11_2/XI0/XI0_18/d_2_ XI11_2/XI0/XI0_18/d__2_ DECAP_INV_G11
XG12085 XI11_2/XI0/XI0_18/d_1_ XI11_2/XI0/XI0_18/d__1_ DECAP_INV_G11
XG12086 XI11_2/XI0/XI0_18/d_0_ XI11_2/XI0/XI0_18/d__0_ DECAP_INV_G11
XG12087 XI11_2/XI0/XI0_17/d__15_ XI11_2/XI0/XI0_17/d_15_ DECAP_INV_G11
XG12088 XI11_2/XI0/XI0_17/d__14_ XI11_2/XI0/XI0_17/d_14_ DECAP_INV_G11
XG12089 XI11_2/XI0/XI0_17/d__13_ XI11_2/XI0/XI0_17/d_13_ DECAP_INV_G11
XG12090 XI11_2/XI0/XI0_17/d__12_ XI11_2/XI0/XI0_17/d_12_ DECAP_INV_G11
XG12091 XI11_2/XI0/XI0_17/d__11_ XI11_2/XI0/XI0_17/d_11_ DECAP_INV_G11
XG12092 XI11_2/XI0/XI0_17/d__10_ XI11_2/XI0/XI0_17/d_10_ DECAP_INV_G11
XG12093 XI11_2/XI0/XI0_17/d__9_ XI11_2/XI0/XI0_17/d_9_ DECAP_INV_G11
XG12094 XI11_2/XI0/XI0_17/d__8_ XI11_2/XI0/XI0_17/d_8_ DECAP_INV_G11
XG12095 XI11_2/XI0/XI0_17/d__7_ XI11_2/XI0/XI0_17/d_7_ DECAP_INV_G11
XG12096 XI11_2/XI0/XI0_17/d__6_ XI11_2/XI0/XI0_17/d_6_ DECAP_INV_G11
XG12097 XI11_2/XI0/XI0_17/d__5_ XI11_2/XI0/XI0_17/d_5_ DECAP_INV_G11
XG12098 XI11_2/XI0/XI0_17/d__4_ XI11_2/XI0/XI0_17/d_4_ DECAP_INV_G11
XG12099 XI11_2/XI0/XI0_17/d__3_ XI11_2/XI0/XI0_17/d_3_ DECAP_INV_G11
XG12100 XI11_2/XI0/XI0_17/d__2_ XI11_2/XI0/XI0_17/d_2_ DECAP_INV_G11
XG12101 XI11_2/XI0/XI0_17/d__1_ XI11_2/XI0/XI0_17/d_1_ DECAP_INV_G11
XG12102 XI11_2/XI0/XI0_17/d__0_ XI11_2/XI0/XI0_17/d_0_ DECAP_INV_G11
XG12103 XI11_2/XI0/XI0_17/d_15_ XI11_2/XI0/XI0_17/d__15_ DECAP_INV_G11
XG12104 XI11_2/XI0/XI0_17/d_14_ XI11_2/XI0/XI0_17/d__14_ DECAP_INV_G11
XG12105 XI11_2/XI0/XI0_17/d_13_ XI11_2/XI0/XI0_17/d__13_ DECAP_INV_G11
XG12106 XI11_2/XI0/XI0_17/d_12_ XI11_2/XI0/XI0_17/d__12_ DECAP_INV_G11
XG12107 XI11_2/XI0/XI0_17/d_11_ XI11_2/XI0/XI0_17/d__11_ DECAP_INV_G11
XG12108 XI11_2/XI0/XI0_17/d_10_ XI11_2/XI0/XI0_17/d__10_ DECAP_INV_G11
XG12109 XI11_2/XI0/XI0_17/d_9_ XI11_2/XI0/XI0_17/d__9_ DECAP_INV_G11
XG12110 XI11_2/XI0/XI0_17/d_8_ XI11_2/XI0/XI0_17/d__8_ DECAP_INV_G11
XG12111 XI11_2/XI0/XI0_17/d_7_ XI11_2/XI0/XI0_17/d__7_ DECAP_INV_G11
XG12112 XI11_2/XI0/XI0_17/d_6_ XI11_2/XI0/XI0_17/d__6_ DECAP_INV_G11
XG12113 XI11_2/XI0/XI0_17/d_5_ XI11_2/XI0/XI0_17/d__5_ DECAP_INV_G11
XG12114 XI11_2/XI0/XI0_17/d_4_ XI11_2/XI0/XI0_17/d__4_ DECAP_INV_G11
XG12115 XI11_2/XI0/XI0_17/d_3_ XI11_2/XI0/XI0_17/d__3_ DECAP_INV_G11
XG12116 XI11_2/XI0/XI0_17/d_2_ XI11_2/XI0/XI0_17/d__2_ DECAP_INV_G11
XG12117 XI11_2/XI0/XI0_17/d_1_ XI11_2/XI0/XI0_17/d__1_ DECAP_INV_G11
XG12118 XI11_2/XI0/XI0_17/d_0_ XI11_2/XI0/XI0_17/d__0_ DECAP_INV_G11
XG12119 XI11_2/XI0/XI0_16/d__15_ XI11_2/XI0/XI0_16/d_15_ DECAP_INV_G11
XG12120 XI11_2/XI0/XI0_16/d__14_ XI11_2/XI0/XI0_16/d_14_ DECAP_INV_G11
XG12121 XI11_2/XI0/XI0_16/d__13_ XI11_2/XI0/XI0_16/d_13_ DECAP_INV_G11
XG12122 XI11_2/XI0/XI0_16/d__12_ XI11_2/XI0/XI0_16/d_12_ DECAP_INV_G11
XG12123 XI11_2/XI0/XI0_16/d__11_ XI11_2/XI0/XI0_16/d_11_ DECAP_INV_G11
XG12124 XI11_2/XI0/XI0_16/d__10_ XI11_2/XI0/XI0_16/d_10_ DECAP_INV_G11
XG12125 XI11_2/XI0/XI0_16/d__9_ XI11_2/XI0/XI0_16/d_9_ DECAP_INV_G11
XG12126 XI11_2/XI0/XI0_16/d__8_ XI11_2/XI0/XI0_16/d_8_ DECAP_INV_G11
XG12127 XI11_2/XI0/XI0_16/d__7_ XI11_2/XI0/XI0_16/d_7_ DECAP_INV_G11
XG12128 XI11_2/XI0/XI0_16/d__6_ XI11_2/XI0/XI0_16/d_6_ DECAP_INV_G11
XG12129 XI11_2/XI0/XI0_16/d__5_ XI11_2/XI0/XI0_16/d_5_ DECAP_INV_G11
XG12130 XI11_2/XI0/XI0_16/d__4_ XI11_2/XI0/XI0_16/d_4_ DECAP_INV_G11
XG12131 XI11_2/XI0/XI0_16/d__3_ XI11_2/XI0/XI0_16/d_3_ DECAP_INV_G11
XG12132 XI11_2/XI0/XI0_16/d__2_ XI11_2/XI0/XI0_16/d_2_ DECAP_INV_G11
XG12133 XI11_2/XI0/XI0_16/d__1_ XI11_2/XI0/XI0_16/d_1_ DECAP_INV_G11
XG12134 XI11_2/XI0/XI0_16/d__0_ XI11_2/XI0/XI0_16/d_0_ DECAP_INV_G11
XG12135 XI11_2/XI0/XI0_16/d_15_ XI11_2/XI0/XI0_16/d__15_ DECAP_INV_G11
XG12136 XI11_2/XI0/XI0_16/d_14_ XI11_2/XI0/XI0_16/d__14_ DECAP_INV_G11
XG12137 XI11_2/XI0/XI0_16/d_13_ XI11_2/XI0/XI0_16/d__13_ DECAP_INV_G11
XG12138 XI11_2/XI0/XI0_16/d_12_ XI11_2/XI0/XI0_16/d__12_ DECAP_INV_G11
XG12139 XI11_2/XI0/XI0_16/d_11_ XI11_2/XI0/XI0_16/d__11_ DECAP_INV_G11
XG12140 XI11_2/XI0/XI0_16/d_10_ XI11_2/XI0/XI0_16/d__10_ DECAP_INV_G11
XG12141 XI11_2/XI0/XI0_16/d_9_ XI11_2/XI0/XI0_16/d__9_ DECAP_INV_G11
XG12142 XI11_2/XI0/XI0_16/d_8_ XI11_2/XI0/XI0_16/d__8_ DECAP_INV_G11
XG12143 XI11_2/XI0/XI0_16/d_7_ XI11_2/XI0/XI0_16/d__7_ DECAP_INV_G11
XG12144 XI11_2/XI0/XI0_16/d_6_ XI11_2/XI0/XI0_16/d__6_ DECAP_INV_G11
XG12145 XI11_2/XI0/XI0_16/d_5_ XI11_2/XI0/XI0_16/d__5_ DECAP_INV_G11
XG12146 XI11_2/XI0/XI0_16/d_4_ XI11_2/XI0/XI0_16/d__4_ DECAP_INV_G11
XG12147 XI11_2/XI0/XI0_16/d_3_ XI11_2/XI0/XI0_16/d__3_ DECAP_INV_G11
XG12148 XI11_2/XI0/XI0_16/d_2_ XI11_2/XI0/XI0_16/d__2_ DECAP_INV_G11
XG12149 XI11_2/XI0/XI0_16/d_1_ XI11_2/XI0/XI0_16/d__1_ DECAP_INV_G11
XG12150 XI11_2/XI0/XI0_16/d_0_ XI11_2/XI0/XI0_16/d__0_ DECAP_INV_G11
XG12151 XI11_2/XI0/XI0_15/d__15_ XI11_2/XI0/XI0_15/d_15_ DECAP_INV_G11
XG12152 XI11_2/XI0/XI0_15/d__14_ XI11_2/XI0/XI0_15/d_14_ DECAP_INV_G11
XG12153 XI11_2/XI0/XI0_15/d__13_ XI11_2/XI0/XI0_15/d_13_ DECAP_INV_G11
XG12154 XI11_2/XI0/XI0_15/d__12_ XI11_2/XI0/XI0_15/d_12_ DECAP_INV_G11
XG12155 XI11_2/XI0/XI0_15/d__11_ XI11_2/XI0/XI0_15/d_11_ DECAP_INV_G11
XG12156 XI11_2/XI0/XI0_15/d__10_ XI11_2/XI0/XI0_15/d_10_ DECAP_INV_G11
XG12157 XI11_2/XI0/XI0_15/d__9_ XI11_2/XI0/XI0_15/d_9_ DECAP_INV_G11
XG12158 XI11_2/XI0/XI0_15/d__8_ XI11_2/XI0/XI0_15/d_8_ DECAP_INV_G11
XG12159 XI11_2/XI0/XI0_15/d__7_ XI11_2/XI0/XI0_15/d_7_ DECAP_INV_G11
XG12160 XI11_2/XI0/XI0_15/d__6_ XI11_2/XI0/XI0_15/d_6_ DECAP_INV_G11
XG12161 XI11_2/XI0/XI0_15/d__5_ XI11_2/XI0/XI0_15/d_5_ DECAP_INV_G11
XG12162 XI11_2/XI0/XI0_15/d__4_ XI11_2/XI0/XI0_15/d_4_ DECAP_INV_G11
XG12163 XI11_2/XI0/XI0_15/d__3_ XI11_2/XI0/XI0_15/d_3_ DECAP_INV_G11
XG12164 XI11_2/XI0/XI0_15/d__2_ XI11_2/XI0/XI0_15/d_2_ DECAP_INV_G11
XG12165 XI11_2/XI0/XI0_15/d__1_ XI11_2/XI0/XI0_15/d_1_ DECAP_INV_G11
XG12166 XI11_2/XI0/XI0_15/d__0_ XI11_2/XI0/XI0_15/d_0_ DECAP_INV_G11
XG12167 XI11_2/XI0/XI0_15/d_15_ XI11_2/XI0/XI0_15/d__15_ DECAP_INV_G11
XG12168 XI11_2/XI0/XI0_15/d_14_ XI11_2/XI0/XI0_15/d__14_ DECAP_INV_G11
XG12169 XI11_2/XI0/XI0_15/d_13_ XI11_2/XI0/XI0_15/d__13_ DECAP_INV_G11
XG12170 XI11_2/XI0/XI0_15/d_12_ XI11_2/XI0/XI0_15/d__12_ DECAP_INV_G11
XG12171 XI11_2/XI0/XI0_15/d_11_ XI11_2/XI0/XI0_15/d__11_ DECAP_INV_G11
XG12172 XI11_2/XI0/XI0_15/d_10_ XI11_2/XI0/XI0_15/d__10_ DECAP_INV_G11
XG12173 XI11_2/XI0/XI0_15/d_9_ XI11_2/XI0/XI0_15/d__9_ DECAP_INV_G11
XG12174 XI11_2/XI0/XI0_15/d_8_ XI11_2/XI0/XI0_15/d__8_ DECAP_INV_G11
XG12175 XI11_2/XI0/XI0_15/d_7_ XI11_2/XI0/XI0_15/d__7_ DECAP_INV_G11
XG12176 XI11_2/XI0/XI0_15/d_6_ XI11_2/XI0/XI0_15/d__6_ DECAP_INV_G11
XG12177 XI11_2/XI0/XI0_15/d_5_ XI11_2/XI0/XI0_15/d__5_ DECAP_INV_G11
XG12178 XI11_2/XI0/XI0_15/d_4_ XI11_2/XI0/XI0_15/d__4_ DECAP_INV_G11
XG12179 XI11_2/XI0/XI0_15/d_3_ XI11_2/XI0/XI0_15/d__3_ DECAP_INV_G11
XG12180 XI11_2/XI0/XI0_15/d_2_ XI11_2/XI0/XI0_15/d__2_ DECAP_INV_G11
XG12181 XI11_2/XI0/XI0_15/d_1_ XI11_2/XI0/XI0_15/d__1_ DECAP_INV_G11
XG12182 XI11_2/XI0/XI0_15/d_0_ XI11_2/XI0/XI0_15/d__0_ DECAP_INV_G11
XG12183 XI11_2/XI0/XI0_14/d__15_ XI11_2/XI0/XI0_14/d_15_ DECAP_INV_G11
XG12184 XI11_2/XI0/XI0_14/d__14_ XI11_2/XI0/XI0_14/d_14_ DECAP_INV_G11
XG12185 XI11_2/XI0/XI0_14/d__13_ XI11_2/XI0/XI0_14/d_13_ DECAP_INV_G11
XG12186 XI11_2/XI0/XI0_14/d__12_ XI11_2/XI0/XI0_14/d_12_ DECAP_INV_G11
XG12187 XI11_2/XI0/XI0_14/d__11_ XI11_2/XI0/XI0_14/d_11_ DECAP_INV_G11
XG12188 XI11_2/XI0/XI0_14/d__10_ XI11_2/XI0/XI0_14/d_10_ DECAP_INV_G11
XG12189 XI11_2/XI0/XI0_14/d__9_ XI11_2/XI0/XI0_14/d_9_ DECAP_INV_G11
XG12190 XI11_2/XI0/XI0_14/d__8_ XI11_2/XI0/XI0_14/d_8_ DECAP_INV_G11
XG12191 XI11_2/XI0/XI0_14/d__7_ XI11_2/XI0/XI0_14/d_7_ DECAP_INV_G11
XG12192 XI11_2/XI0/XI0_14/d__6_ XI11_2/XI0/XI0_14/d_6_ DECAP_INV_G11
XG12193 XI11_2/XI0/XI0_14/d__5_ XI11_2/XI0/XI0_14/d_5_ DECAP_INV_G11
XG12194 XI11_2/XI0/XI0_14/d__4_ XI11_2/XI0/XI0_14/d_4_ DECAP_INV_G11
XG12195 XI11_2/XI0/XI0_14/d__3_ XI11_2/XI0/XI0_14/d_3_ DECAP_INV_G11
XG12196 XI11_2/XI0/XI0_14/d__2_ XI11_2/XI0/XI0_14/d_2_ DECAP_INV_G11
XG12197 XI11_2/XI0/XI0_14/d__1_ XI11_2/XI0/XI0_14/d_1_ DECAP_INV_G11
XG12198 XI11_2/XI0/XI0_14/d__0_ XI11_2/XI0/XI0_14/d_0_ DECAP_INV_G11
XG12199 XI11_2/XI0/XI0_14/d_15_ XI11_2/XI0/XI0_14/d__15_ DECAP_INV_G11
XG12200 XI11_2/XI0/XI0_14/d_14_ XI11_2/XI0/XI0_14/d__14_ DECAP_INV_G11
XG12201 XI11_2/XI0/XI0_14/d_13_ XI11_2/XI0/XI0_14/d__13_ DECAP_INV_G11
XG12202 XI11_2/XI0/XI0_14/d_12_ XI11_2/XI0/XI0_14/d__12_ DECAP_INV_G11
XG12203 XI11_2/XI0/XI0_14/d_11_ XI11_2/XI0/XI0_14/d__11_ DECAP_INV_G11
XG12204 XI11_2/XI0/XI0_14/d_10_ XI11_2/XI0/XI0_14/d__10_ DECAP_INV_G11
XG12205 XI11_2/XI0/XI0_14/d_9_ XI11_2/XI0/XI0_14/d__9_ DECAP_INV_G11
XG12206 XI11_2/XI0/XI0_14/d_8_ XI11_2/XI0/XI0_14/d__8_ DECAP_INV_G11
XG12207 XI11_2/XI0/XI0_14/d_7_ XI11_2/XI0/XI0_14/d__7_ DECAP_INV_G11
XG12208 XI11_2/XI0/XI0_14/d_6_ XI11_2/XI0/XI0_14/d__6_ DECAP_INV_G11
XG12209 XI11_2/XI0/XI0_14/d_5_ XI11_2/XI0/XI0_14/d__5_ DECAP_INV_G11
XG12210 XI11_2/XI0/XI0_14/d_4_ XI11_2/XI0/XI0_14/d__4_ DECAP_INV_G11
XG12211 XI11_2/XI0/XI0_14/d_3_ XI11_2/XI0/XI0_14/d__3_ DECAP_INV_G11
XG12212 XI11_2/XI0/XI0_14/d_2_ XI11_2/XI0/XI0_14/d__2_ DECAP_INV_G11
XG12213 XI11_2/XI0/XI0_14/d_1_ XI11_2/XI0/XI0_14/d__1_ DECAP_INV_G11
XG12214 XI11_2/XI0/XI0_14/d_0_ XI11_2/XI0/XI0_14/d__0_ DECAP_INV_G11
XG12215 XI11_2/XI0/XI0_13/d__15_ XI11_2/XI0/XI0_13/d_15_ DECAP_INV_G11
XG12216 XI11_2/XI0/XI0_13/d__14_ XI11_2/XI0/XI0_13/d_14_ DECAP_INV_G11
XG12217 XI11_2/XI0/XI0_13/d__13_ XI11_2/XI0/XI0_13/d_13_ DECAP_INV_G11
XG12218 XI11_2/XI0/XI0_13/d__12_ XI11_2/XI0/XI0_13/d_12_ DECAP_INV_G11
XG12219 XI11_2/XI0/XI0_13/d__11_ XI11_2/XI0/XI0_13/d_11_ DECAP_INV_G11
XG12220 XI11_2/XI0/XI0_13/d__10_ XI11_2/XI0/XI0_13/d_10_ DECAP_INV_G11
XG12221 XI11_2/XI0/XI0_13/d__9_ XI11_2/XI0/XI0_13/d_9_ DECAP_INV_G11
XG12222 XI11_2/XI0/XI0_13/d__8_ XI11_2/XI0/XI0_13/d_8_ DECAP_INV_G11
XG12223 XI11_2/XI0/XI0_13/d__7_ XI11_2/XI0/XI0_13/d_7_ DECAP_INV_G11
XG12224 XI11_2/XI0/XI0_13/d__6_ XI11_2/XI0/XI0_13/d_6_ DECAP_INV_G11
XG12225 XI11_2/XI0/XI0_13/d__5_ XI11_2/XI0/XI0_13/d_5_ DECAP_INV_G11
XG12226 XI11_2/XI0/XI0_13/d__4_ XI11_2/XI0/XI0_13/d_4_ DECAP_INV_G11
XG12227 XI11_2/XI0/XI0_13/d__3_ XI11_2/XI0/XI0_13/d_3_ DECAP_INV_G11
XG12228 XI11_2/XI0/XI0_13/d__2_ XI11_2/XI0/XI0_13/d_2_ DECAP_INV_G11
XG12229 XI11_2/XI0/XI0_13/d__1_ XI11_2/XI0/XI0_13/d_1_ DECAP_INV_G11
XG12230 XI11_2/XI0/XI0_13/d__0_ XI11_2/XI0/XI0_13/d_0_ DECAP_INV_G11
XG12231 XI11_2/XI0/XI0_13/d_15_ XI11_2/XI0/XI0_13/d__15_ DECAP_INV_G11
XG12232 XI11_2/XI0/XI0_13/d_14_ XI11_2/XI0/XI0_13/d__14_ DECAP_INV_G11
XG12233 XI11_2/XI0/XI0_13/d_13_ XI11_2/XI0/XI0_13/d__13_ DECAP_INV_G11
XG12234 XI11_2/XI0/XI0_13/d_12_ XI11_2/XI0/XI0_13/d__12_ DECAP_INV_G11
XG12235 XI11_2/XI0/XI0_13/d_11_ XI11_2/XI0/XI0_13/d__11_ DECAP_INV_G11
XG12236 XI11_2/XI0/XI0_13/d_10_ XI11_2/XI0/XI0_13/d__10_ DECAP_INV_G11
XG12237 XI11_2/XI0/XI0_13/d_9_ XI11_2/XI0/XI0_13/d__9_ DECAP_INV_G11
XG12238 XI11_2/XI0/XI0_13/d_8_ XI11_2/XI0/XI0_13/d__8_ DECAP_INV_G11
XG12239 XI11_2/XI0/XI0_13/d_7_ XI11_2/XI0/XI0_13/d__7_ DECAP_INV_G11
XG12240 XI11_2/XI0/XI0_13/d_6_ XI11_2/XI0/XI0_13/d__6_ DECAP_INV_G11
XG12241 XI11_2/XI0/XI0_13/d_5_ XI11_2/XI0/XI0_13/d__5_ DECAP_INV_G11
XG12242 XI11_2/XI0/XI0_13/d_4_ XI11_2/XI0/XI0_13/d__4_ DECAP_INV_G11
XG12243 XI11_2/XI0/XI0_13/d_3_ XI11_2/XI0/XI0_13/d__3_ DECAP_INV_G11
XG12244 XI11_2/XI0/XI0_13/d_2_ XI11_2/XI0/XI0_13/d__2_ DECAP_INV_G11
XG12245 XI11_2/XI0/XI0_13/d_1_ XI11_2/XI0/XI0_13/d__1_ DECAP_INV_G11
XG12246 XI11_2/XI0/XI0_13/d_0_ XI11_2/XI0/XI0_13/d__0_ DECAP_INV_G11
XG12247 XI11_2/XI0/XI0_12/d__15_ XI11_2/XI0/XI0_12/d_15_ DECAP_INV_G11
XG12248 XI11_2/XI0/XI0_12/d__14_ XI11_2/XI0/XI0_12/d_14_ DECAP_INV_G11
XG12249 XI11_2/XI0/XI0_12/d__13_ XI11_2/XI0/XI0_12/d_13_ DECAP_INV_G11
XG12250 XI11_2/XI0/XI0_12/d__12_ XI11_2/XI0/XI0_12/d_12_ DECAP_INV_G11
XG12251 XI11_2/XI0/XI0_12/d__11_ XI11_2/XI0/XI0_12/d_11_ DECAP_INV_G11
XG12252 XI11_2/XI0/XI0_12/d__10_ XI11_2/XI0/XI0_12/d_10_ DECAP_INV_G11
XG12253 XI11_2/XI0/XI0_12/d__9_ XI11_2/XI0/XI0_12/d_9_ DECAP_INV_G11
XG12254 XI11_2/XI0/XI0_12/d__8_ XI11_2/XI0/XI0_12/d_8_ DECAP_INV_G11
XG12255 XI11_2/XI0/XI0_12/d__7_ XI11_2/XI0/XI0_12/d_7_ DECAP_INV_G11
XG12256 XI11_2/XI0/XI0_12/d__6_ XI11_2/XI0/XI0_12/d_6_ DECAP_INV_G11
XG12257 XI11_2/XI0/XI0_12/d__5_ XI11_2/XI0/XI0_12/d_5_ DECAP_INV_G11
XG12258 XI11_2/XI0/XI0_12/d__4_ XI11_2/XI0/XI0_12/d_4_ DECAP_INV_G11
XG12259 XI11_2/XI0/XI0_12/d__3_ XI11_2/XI0/XI0_12/d_3_ DECAP_INV_G11
XG12260 XI11_2/XI0/XI0_12/d__2_ XI11_2/XI0/XI0_12/d_2_ DECAP_INV_G11
XG12261 XI11_2/XI0/XI0_12/d__1_ XI11_2/XI0/XI0_12/d_1_ DECAP_INV_G11
XG12262 XI11_2/XI0/XI0_12/d__0_ XI11_2/XI0/XI0_12/d_0_ DECAP_INV_G11
XG12263 XI11_2/XI0/XI0_12/d_15_ XI11_2/XI0/XI0_12/d__15_ DECAP_INV_G11
XG12264 XI11_2/XI0/XI0_12/d_14_ XI11_2/XI0/XI0_12/d__14_ DECAP_INV_G11
XG12265 XI11_2/XI0/XI0_12/d_13_ XI11_2/XI0/XI0_12/d__13_ DECAP_INV_G11
XG12266 XI11_2/XI0/XI0_12/d_12_ XI11_2/XI0/XI0_12/d__12_ DECAP_INV_G11
XG12267 XI11_2/XI0/XI0_12/d_11_ XI11_2/XI0/XI0_12/d__11_ DECAP_INV_G11
XG12268 XI11_2/XI0/XI0_12/d_10_ XI11_2/XI0/XI0_12/d__10_ DECAP_INV_G11
XG12269 XI11_2/XI0/XI0_12/d_9_ XI11_2/XI0/XI0_12/d__9_ DECAP_INV_G11
XG12270 XI11_2/XI0/XI0_12/d_8_ XI11_2/XI0/XI0_12/d__8_ DECAP_INV_G11
XG12271 XI11_2/XI0/XI0_12/d_7_ XI11_2/XI0/XI0_12/d__7_ DECAP_INV_G11
XG12272 XI11_2/XI0/XI0_12/d_6_ XI11_2/XI0/XI0_12/d__6_ DECAP_INV_G11
XG12273 XI11_2/XI0/XI0_12/d_5_ XI11_2/XI0/XI0_12/d__5_ DECAP_INV_G11
XG12274 XI11_2/XI0/XI0_12/d_4_ XI11_2/XI0/XI0_12/d__4_ DECAP_INV_G11
XG12275 XI11_2/XI0/XI0_12/d_3_ XI11_2/XI0/XI0_12/d__3_ DECAP_INV_G11
XG12276 XI11_2/XI0/XI0_12/d_2_ XI11_2/XI0/XI0_12/d__2_ DECAP_INV_G11
XG12277 XI11_2/XI0/XI0_12/d_1_ XI11_2/XI0/XI0_12/d__1_ DECAP_INV_G11
XG12278 XI11_2/XI0/XI0_12/d_0_ XI11_2/XI0/XI0_12/d__0_ DECAP_INV_G11
XG12279 XI11_2/XI0/XI0_11/d__15_ XI11_2/XI0/XI0_11/d_15_ DECAP_INV_G11
XG12280 XI11_2/XI0/XI0_11/d__14_ XI11_2/XI0/XI0_11/d_14_ DECAP_INV_G11
XG12281 XI11_2/XI0/XI0_11/d__13_ XI11_2/XI0/XI0_11/d_13_ DECAP_INV_G11
XG12282 XI11_2/XI0/XI0_11/d__12_ XI11_2/XI0/XI0_11/d_12_ DECAP_INV_G11
XG12283 XI11_2/XI0/XI0_11/d__11_ XI11_2/XI0/XI0_11/d_11_ DECAP_INV_G11
XG12284 XI11_2/XI0/XI0_11/d__10_ XI11_2/XI0/XI0_11/d_10_ DECAP_INV_G11
XG12285 XI11_2/XI0/XI0_11/d__9_ XI11_2/XI0/XI0_11/d_9_ DECAP_INV_G11
XG12286 XI11_2/XI0/XI0_11/d__8_ XI11_2/XI0/XI0_11/d_8_ DECAP_INV_G11
XG12287 XI11_2/XI0/XI0_11/d__7_ XI11_2/XI0/XI0_11/d_7_ DECAP_INV_G11
XG12288 XI11_2/XI0/XI0_11/d__6_ XI11_2/XI0/XI0_11/d_6_ DECAP_INV_G11
XG12289 XI11_2/XI0/XI0_11/d__5_ XI11_2/XI0/XI0_11/d_5_ DECAP_INV_G11
XG12290 XI11_2/XI0/XI0_11/d__4_ XI11_2/XI0/XI0_11/d_4_ DECAP_INV_G11
XG12291 XI11_2/XI0/XI0_11/d__3_ XI11_2/XI0/XI0_11/d_3_ DECAP_INV_G11
XG12292 XI11_2/XI0/XI0_11/d__2_ XI11_2/XI0/XI0_11/d_2_ DECAP_INV_G11
XG12293 XI11_2/XI0/XI0_11/d__1_ XI11_2/XI0/XI0_11/d_1_ DECAP_INV_G11
XG12294 XI11_2/XI0/XI0_11/d__0_ XI11_2/XI0/XI0_11/d_0_ DECAP_INV_G11
XG12295 XI11_2/XI0/XI0_11/d_15_ XI11_2/XI0/XI0_11/d__15_ DECAP_INV_G11
XG12296 XI11_2/XI0/XI0_11/d_14_ XI11_2/XI0/XI0_11/d__14_ DECAP_INV_G11
XG12297 XI11_2/XI0/XI0_11/d_13_ XI11_2/XI0/XI0_11/d__13_ DECAP_INV_G11
XG12298 XI11_2/XI0/XI0_11/d_12_ XI11_2/XI0/XI0_11/d__12_ DECAP_INV_G11
XG12299 XI11_2/XI0/XI0_11/d_11_ XI11_2/XI0/XI0_11/d__11_ DECAP_INV_G11
XG12300 XI11_2/XI0/XI0_11/d_10_ XI11_2/XI0/XI0_11/d__10_ DECAP_INV_G11
XG12301 XI11_2/XI0/XI0_11/d_9_ XI11_2/XI0/XI0_11/d__9_ DECAP_INV_G11
XG12302 XI11_2/XI0/XI0_11/d_8_ XI11_2/XI0/XI0_11/d__8_ DECAP_INV_G11
XG12303 XI11_2/XI0/XI0_11/d_7_ XI11_2/XI0/XI0_11/d__7_ DECAP_INV_G11
XG12304 XI11_2/XI0/XI0_11/d_6_ XI11_2/XI0/XI0_11/d__6_ DECAP_INV_G11
XG12305 XI11_2/XI0/XI0_11/d_5_ XI11_2/XI0/XI0_11/d__5_ DECAP_INV_G11
XG12306 XI11_2/XI0/XI0_11/d_4_ XI11_2/XI0/XI0_11/d__4_ DECAP_INV_G11
XG12307 XI11_2/XI0/XI0_11/d_3_ XI11_2/XI0/XI0_11/d__3_ DECAP_INV_G11
XG12308 XI11_2/XI0/XI0_11/d_2_ XI11_2/XI0/XI0_11/d__2_ DECAP_INV_G11
XG12309 XI11_2/XI0/XI0_11/d_1_ XI11_2/XI0/XI0_11/d__1_ DECAP_INV_G11
XG12310 XI11_2/XI0/XI0_11/d_0_ XI11_2/XI0/XI0_11/d__0_ DECAP_INV_G11
XG12311 XI11_2/XI0/XI0_10/d__15_ XI11_2/XI0/XI0_10/d_15_ DECAP_INV_G11
XG12312 XI11_2/XI0/XI0_10/d__14_ XI11_2/XI0/XI0_10/d_14_ DECAP_INV_G11
XG12313 XI11_2/XI0/XI0_10/d__13_ XI11_2/XI0/XI0_10/d_13_ DECAP_INV_G11
XG12314 XI11_2/XI0/XI0_10/d__12_ XI11_2/XI0/XI0_10/d_12_ DECAP_INV_G11
XG12315 XI11_2/XI0/XI0_10/d__11_ XI11_2/XI0/XI0_10/d_11_ DECAP_INV_G11
XG12316 XI11_2/XI0/XI0_10/d__10_ XI11_2/XI0/XI0_10/d_10_ DECAP_INV_G11
XG12317 XI11_2/XI0/XI0_10/d__9_ XI11_2/XI0/XI0_10/d_9_ DECAP_INV_G11
XG12318 XI11_2/XI0/XI0_10/d__8_ XI11_2/XI0/XI0_10/d_8_ DECAP_INV_G11
XG12319 XI11_2/XI0/XI0_10/d__7_ XI11_2/XI0/XI0_10/d_7_ DECAP_INV_G11
XG12320 XI11_2/XI0/XI0_10/d__6_ XI11_2/XI0/XI0_10/d_6_ DECAP_INV_G11
XG12321 XI11_2/XI0/XI0_10/d__5_ XI11_2/XI0/XI0_10/d_5_ DECAP_INV_G11
XG12322 XI11_2/XI0/XI0_10/d__4_ XI11_2/XI0/XI0_10/d_4_ DECAP_INV_G11
XG12323 XI11_2/XI0/XI0_10/d__3_ XI11_2/XI0/XI0_10/d_3_ DECAP_INV_G11
XG12324 XI11_2/XI0/XI0_10/d__2_ XI11_2/XI0/XI0_10/d_2_ DECAP_INV_G11
XG12325 XI11_2/XI0/XI0_10/d__1_ XI11_2/XI0/XI0_10/d_1_ DECAP_INV_G11
XG12326 XI11_2/XI0/XI0_10/d__0_ XI11_2/XI0/XI0_10/d_0_ DECAP_INV_G11
XG12327 XI11_2/XI0/XI0_10/d_15_ XI11_2/XI0/XI0_10/d__15_ DECAP_INV_G11
XG12328 XI11_2/XI0/XI0_10/d_14_ XI11_2/XI0/XI0_10/d__14_ DECAP_INV_G11
XG12329 XI11_2/XI0/XI0_10/d_13_ XI11_2/XI0/XI0_10/d__13_ DECAP_INV_G11
XG12330 XI11_2/XI0/XI0_10/d_12_ XI11_2/XI0/XI0_10/d__12_ DECAP_INV_G11
XG12331 XI11_2/XI0/XI0_10/d_11_ XI11_2/XI0/XI0_10/d__11_ DECAP_INV_G11
XG12332 XI11_2/XI0/XI0_10/d_10_ XI11_2/XI0/XI0_10/d__10_ DECAP_INV_G11
XG12333 XI11_2/XI0/XI0_10/d_9_ XI11_2/XI0/XI0_10/d__9_ DECAP_INV_G11
XG12334 XI11_2/XI0/XI0_10/d_8_ XI11_2/XI0/XI0_10/d__8_ DECAP_INV_G11
XG12335 XI11_2/XI0/XI0_10/d_7_ XI11_2/XI0/XI0_10/d__7_ DECAP_INV_G11
XG12336 XI11_2/XI0/XI0_10/d_6_ XI11_2/XI0/XI0_10/d__6_ DECAP_INV_G11
XG12337 XI11_2/XI0/XI0_10/d_5_ XI11_2/XI0/XI0_10/d__5_ DECAP_INV_G11
XG12338 XI11_2/XI0/XI0_10/d_4_ XI11_2/XI0/XI0_10/d__4_ DECAP_INV_G11
XG12339 XI11_2/XI0/XI0_10/d_3_ XI11_2/XI0/XI0_10/d__3_ DECAP_INV_G11
XG12340 XI11_2/XI0/XI0_10/d_2_ XI11_2/XI0/XI0_10/d__2_ DECAP_INV_G11
XG12341 XI11_2/XI0/XI0_10/d_1_ XI11_2/XI0/XI0_10/d__1_ DECAP_INV_G11
XG12342 XI11_2/XI0/XI0_10/d_0_ XI11_2/XI0/XI0_10/d__0_ DECAP_INV_G11
XG12343 XI11_2/XI0/XI0_9/d__15_ XI11_2/XI0/XI0_9/d_15_ DECAP_INV_G11
XG12344 XI11_2/XI0/XI0_9/d__14_ XI11_2/XI0/XI0_9/d_14_ DECAP_INV_G11
XG12345 XI11_2/XI0/XI0_9/d__13_ XI11_2/XI0/XI0_9/d_13_ DECAP_INV_G11
XG12346 XI11_2/XI0/XI0_9/d__12_ XI11_2/XI0/XI0_9/d_12_ DECAP_INV_G11
XG12347 XI11_2/XI0/XI0_9/d__11_ XI11_2/XI0/XI0_9/d_11_ DECAP_INV_G11
XG12348 XI11_2/XI0/XI0_9/d__10_ XI11_2/XI0/XI0_9/d_10_ DECAP_INV_G11
XG12349 XI11_2/XI0/XI0_9/d__9_ XI11_2/XI0/XI0_9/d_9_ DECAP_INV_G11
XG12350 XI11_2/XI0/XI0_9/d__8_ XI11_2/XI0/XI0_9/d_8_ DECAP_INV_G11
XG12351 XI11_2/XI0/XI0_9/d__7_ XI11_2/XI0/XI0_9/d_7_ DECAP_INV_G11
XG12352 XI11_2/XI0/XI0_9/d__6_ XI11_2/XI0/XI0_9/d_6_ DECAP_INV_G11
XG12353 XI11_2/XI0/XI0_9/d__5_ XI11_2/XI0/XI0_9/d_5_ DECAP_INV_G11
XG12354 XI11_2/XI0/XI0_9/d__4_ XI11_2/XI0/XI0_9/d_4_ DECAP_INV_G11
XG12355 XI11_2/XI0/XI0_9/d__3_ XI11_2/XI0/XI0_9/d_3_ DECAP_INV_G11
XG12356 XI11_2/XI0/XI0_9/d__2_ XI11_2/XI0/XI0_9/d_2_ DECAP_INV_G11
XG12357 XI11_2/XI0/XI0_9/d__1_ XI11_2/XI0/XI0_9/d_1_ DECAP_INV_G11
XG12358 XI11_2/XI0/XI0_9/d__0_ XI11_2/XI0/XI0_9/d_0_ DECAP_INV_G11
XG12359 XI11_2/XI0/XI0_9/d_15_ XI11_2/XI0/XI0_9/d__15_ DECAP_INV_G11
XG12360 XI11_2/XI0/XI0_9/d_14_ XI11_2/XI0/XI0_9/d__14_ DECAP_INV_G11
XG12361 XI11_2/XI0/XI0_9/d_13_ XI11_2/XI0/XI0_9/d__13_ DECAP_INV_G11
XG12362 XI11_2/XI0/XI0_9/d_12_ XI11_2/XI0/XI0_9/d__12_ DECAP_INV_G11
XG12363 XI11_2/XI0/XI0_9/d_11_ XI11_2/XI0/XI0_9/d__11_ DECAP_INV_G11
XG12364 XI11_2/XI0/XI0_9/d_10_ XI11_2/XI0/XI0_9/d__10_ DECAP_INV_G11
XG12365 XI11_2/XI0/XI0_9/d_9_ XI11_2/XI0/XI0_9/d__9_ DECAP_INV_G11
XG12366 XI11_2/XI0/XI0_9/d_8_ XI11_2/XI0/XI0_9/d__8_ DECAP_INV_G11
XG12367 XI11_2/XI0/XI0_9/d_7_ XI11_2/XI0/XI0_9/d__7_ DECAP_INV_G11
XG12368 XI11_2/XI0/XI0_9/d_6_ XI11_2/XI0/XI0_9/d__6_ DECAP_INV_G11
XG12369 XI11_2/XI0/XI0_9/d_5_ XI11_2/XI0/XI0_9/d__5_ DECAP_INV_G11
XG12370 XI11_2/XI0/XI0_9/d_4_ XI11_2/XI0/XI0_9/d__4_ DECAP_INV_G11
XG12371 XI11_2/XI0/XI0_9/d_3_ XI11_2/XI0/XI0_9/d__3_ DECAP_INV_G11
XG12372 XI11_2/XI0/XI0_9/d_2_ XI11_2/XI0/XI0_9/d__2_ DECAP_INV_G11
XG12373 XI11_2/XI0/XI0_9/d_1_ XI11_2/XI0/XI0_9/d__1_ DECAP_INV_G11
XG12374 XI11_2/XI0/XI0_9/d_0_ XI11_2/XI0/XI0_9/d__0_ DECAP_INV_G11
XG12375 XI11_2/XI0/XI0_8/d__15_ XI11_2/XI0/XI0_8/d_15_ DECAP_INV_G11
XG12376 XI11_2/XI0/XI0_8/d__14_ XI11_2/XI0/XI0_8/d_14_ DECAP_INV_G11
XG12377 XI11_2/XI0/XI0_8/d__13_ XI11_2/XI0/XI0_8/d_13_ DECAP_INV_G11
XG12378 XI11_2/XI0/XI0_8/d__12_ XI11_2/XI0/XI0_8/d_12_ DECAP_INV_G11
XG12379 XI11_2/XI0/XI0_8/d__11_ XI11_2/XI0/XI0_8/d_11_ DECAP_INV_G11
XG12380 XI11_2/XI0/XI0_8/d__10_ XI11_2/XI0/XI0_8/d_10_ DECAP_INV_G11
XG12381 XI11_2/XI0/XI0_8/d__9_ XI11_2/XI0/XI0_8/d_9_ DECAP_INV_G11
XG12382 XI11_2/XI0/XI0_8/d__8_ XI11_2/XI0/XI0_8/d_8_ DECAP_INV_G11
XG12383 XI11_2/XI0/XI0_8/d__7_ XI11_2/XI0/XI0_8/d_7_ DECAP_INV_G11
XG12384 XI11_2/XI0/XI0_8/d__6_ XI11_2/XI0/XI0_8/d_6_ DECAP_INV_G11
XG12385 XI11_2/XI0/XI0_8/d__5_ XI11_2/XI0/XI0_8/d_5_ DECAP_INV_G11
XG12386 XI11_2/XI0/XI0_8/d__4_ XI11_2/XI0/XI0_8/d_4_ DECAP_INV_G11
XG12387 XI11_2/XI0/XI0_8/d__3_ XI11_2/XI0/XI0_8/d_3_ DECAP_INV_G11
XG12388 XI11_2/XI0/XI0_8/d__2_ XI11_2/XI0/XI0_8/d_2_ DECAP_INV_G11
XG12389 XI11_2/XI0/XI0_8/d__1_ XI11_2/XI0/XI0_8/d_1_ DECAP_INV_G11
XG12390 XI11_2/XI0/XI0_8/d__0_ XI11_2/XI0/XI0_8/d_0_ DECAP_INV_G11
XG12391 XI11_2/XI0/XI0_8/d_15_ XI11_2/XI0/XI0_8/d__15_ DECAP_INV_G11
XG12392 XI11_2/XI0/XI0_8/d_14_ XI11_2/XI0/XI0_8/d__14_ DECAP_INV_G11
XG12393 XI11_2/XI0/XI0_8/d_13_ XI11_2/XI0/XI0_8/d__13_ DECAP_INV_G11
XG12394 XI11_2/XI0/XI0_8/d_12_ XI11_2/XI0/XI0_8/d__12_ DECAP_INV_G11
XG12395 XI11_2/XI0/XI0_8/d_11_ XI11_2/XI0/XI0_8/d__11_ DECAP_INV_G11
XG12396 XI11_2/XI0/XI0_8/d_10_ XI11_2/XI0/XI0_8/d__10_ DECAP_INV_G11
XG12397 XI11_2/XI0/XI0_8/d_9_ XI11_2/XI0/XI0_8/d__9_ DECAP_INV_G11
XG12398 XI11_2/XI0/XI0_8/d_8_ XI11_2/XI0/XI0_8/d__8_ DECAP_INV_G11
XG12399 XI11_2/XI0/XI0_8/d_7_ XI11_2/XI0/XI0_8/d__7_ DECAP_INV_G11
XG12400 XI11_2/XI0/XI0_8/d_6_ XI11_2/XI0/XI0_8/d__6_ DECAP_INV_G11
XG12401 XI11_2/XI0/XI0_8/d_5_ XI11_2/XI0/XI0_8/d__5_ DECAP_INV_G11
XG12402 XI11_2/XI0/XI0_8/d_4_ XI11_2/XI0/XI0_8/d__4_ DECAP_INV_G11
XG12403 XI11_2/XI0/XI0_8/d_3_ XI11_2/XI0/XI0_8/d__3_ DECAP_INV_G11
XG12404 XI11_2/XI0/XI0_8/d_2_ XI11_2/XI0/XI0_8/d__2_ DECAP_INV_G11
XG12405 XI11_2/XI0/XI0_8/d_1_ XI11_2/XI0/XI0_8/d__1_ DECAP_INV_G11
XG12406 XI11_2/XI0/XI0_8/d_0_ XI11_2/XI0/XI0_8/d__0_ DECAP_INV_G11
XG12407 XI11_2/XI0/XI0_7/d__15_ XI11_2/XI0/XI0_7/d_15_ DECAP_INV_G11
XG12408 XI11_2/XI0/XI0_7/d__14_ XI11_2/XI0/XI0_7/d_14_ DECAP_INV_G11
XG12409 XI11_2/XI0/XI0_7/d__13_ XI11_2/XI0/XI0_7/d_13_ DECAP_INV_G11
XG12410 XI11_2/XI0/XI0_7/d__12_ XI11_2/XI0/XI0_7/d_12_ DECAP_INV_G11
XG12411 XI11_2/XI0/XI0_7/d__11_ XI11_2/XI0/XI0_7/d_11_ DECAP_INV_G11
XG12412 XI11_2/XI0/XI0_7/d__10_ XI11_2/XI0/XI0_7/d_10_ DECAP_INV_G11
XG12413 XI11_2/XI0/XI0_7/d__9_ XI11_2/XI0/XI0_7/d_9_ DECAP_INV_G11
XG12414 XI11_2/XI0/XI0_7/d__8_ XI11_2/XI0/XI0_7/d_8_ DECAP_INV_G11
XG12415 XI11_2/XI0/XI0_7/d__7_ XI11_2/XI0/XI0_7/d_7_ DECAP_INV_G11
XG12416 XI11_2/XI0/XI0_7/d__6_ XI11_2/XI0/XI0_7/d_6_ DECAP_INV_G11
XG12417 XI11_2/XI0/XI0_7/d__5_ XI11_2/XI0/XI0_7/d_5_ DECAP_INV_G11
XG12418 XI11_2/XI0/XI0_7/d__4_ XI11_2/XI0/XI0_7/d_4_ DECAP_INV_G11
XG12419 XI11_2/XI0/XI0_7/d__3_ XI11_2/XI0/XI0_7/d_3_ DECAP_INV_G11
XG12420 XI11_2/XI0/XI0_7/d__2_ XI11_2/XI0/XI0_7/d_2_ DECAP_INV_G11
XG12421 XI11_2/XI0/XI0_7/d__1_ XI11_2/XI0/XI0_7/d_1_ DECAP_INV_G11
XG12422 XI11_2/XI0/XI0_7/d__0_ XI11_2/XI0/XI0_7/d_0_ DECAP_INV_G11
XG12423 XI11_2/XI0/XI0_7/d_15_ XI11_2/XI0/XI0_7/d__15_ DECAP_INV_G11
XG12424 XI11_2/XI0/XI0_7/d_14_ XI11_2/XI0/XI0_7/d__14_ DECAP_INV_G11
XG12425 XI11_2/XI0/XI0_7/d_13_ XI11_2/XI0/XI0_7/d__13_ DECAP_INV_G11
XG12426 XI11_2/XI0/XI0_7/d_12_ XI11_2/XI0/XI0_7/d__12_ DECAP_INV_G11
XG12427 XI11_2/XI0/XI0_7/d_11_ XI11_2/XI0/XI0_7/d__11_ DECAP_INV_G11
XG12428 XI11_2/XI0/XI0_7/d_10_ XI11_2/XI0/XI0_7/d__10_ DECAP_INV_G11
XG12429 XI11_2/XI0/XI0_7/d_9_ XI11_2/XI0/XI0_7/d__9_ DECAP_INV_G11
XG12430 XI11_2/XI0/XI0_7/d_8_ XI11_2/XI0/XI0_7/d__8_ DECAP_INV_G11
XG12431 XI11_2/XI0/XI0_7/d_7_ XI11_2/XI0/XI0_7/d__7_ DECAP_INV_G11
XG12432 XI11_2/XI0/XI0_7/d_6_ XI11_2/XI0/XI0_7/d__6_ DECAP_INV_G11
XG12433 XI11_2/XI0/XI0_7/d_5_ XI11_2/XI0/XI0_7/d__5_ DECAP_INV_G11
XG12434 XI11_2/XI0/XI0_7/d_4_ XI11_2/XI0/XI0_7/d__4_ DECAP_INV_G11
XG12435 XI11_2/XI0/XI0_7/d_3_ XI11_2/XI0/XI0_7/d__3_ DECAP_INV_G11
XG12436 XI11_2/XI0/XI0_7/d_2_ XI11_2/XI0/XI0_7/d__2_ DECAP_INV_G11
XG12437 XI11_2/XI0/XI0_7/d_1_ XI11_2/XI0/XI0_7/d__1_ DECAP_INV_G11
XG12438 XI11_2/XI0/XI0_7/d_0_ XI11_2/XI0/XI0_7/d__0_ DECAP_INV_G11
XG12439 XI11_2/XI0/XI0_6/d__15_ XI11_2/XI0/XI0_6/d_15_ DECAP_INV_G11
XG12440 XI11_2/XI0/XI0_6/d__14_ XI11_2/XI0/XI0_6/d_14_ DECAP_INV_G11
XG12441 XI11_2/XI0/XI0_6/d__13_ XI11_2/XI0/XI0_6/d_13_ DECAP_INV_G11
XG12442 XI11_2/XI0/XI0_6/d__12_ XI11_2/XI0/XI0_6/d_12_ DECAP_INV_G11
XG12443 XI11_2/XI0/XI0_6/d__11_ XI11_2/XI0/XI0_6/d_11_ DECAP_INV_G11
XG12444 XI11_2/XI0/XI0_6/d__10_ XI11_2/XI0/XI0_6/d_10_ DECAP_INV_G11
XG12445 XI11_2/XI0/XI0_6/d__9_ XI11_2/XI0/XI0_6/d_9_ DECAP_INV_G11
XG12446 XI11_2/XI0/XI0_6/d__8_ XI11_2/XI0/XI0_6/d_8_ DECAP_INV_G11
XG12447 XI11_2/XI0/XI0_6/d__7_ XI11_2/XI0/XI0_6/d_7_ DECAP_INV_G11
XG12448 XI11_2/XI0/XI0_6/d__6_ XI11_2/XI0/XI0_6/d_6_ DECAP_INV_G11
XG12449 XI11_2/XI0/XI0_6/d__5_ XI11_2/XI0/XI0_6/d_5_ DECAP_INV_G11
XG12450 XI11_2/XI0/XI0_6/d__4_ XI11_2/XI0/XI0_6/d_4_ DECAP_INV_G11
XG12451 XI11_2/XI0/XI0_6/d__3_ XI11_2/XI0/XI0_6/d_3_ DECAP_INV_G11
XG12452 XI11_2/XI0/XI0_6/d__2_ XI11_2/XI0/XI0_6/d_2_ DECAP_INV_G11
XG12453 XI11_2/XI0/XI0_6/d__1_ XI11_2/XI0/XI0_6/d_1_ DECAP_INV_G11
XG12454 XI11_2/XI0/XI0_6/d__0_ XI11_2/XI0/XI0_6/d_0_ DECAP_INV_G11
XG12455 XI11_2/XI0/XI0_6/d_15_ XI11_2/XI0/XI0_6/d__15_ DECAP_INV_G11
XG12456 XI11_2/XI0/XI0_6/d_14_ XI11_2/XI0/XI0_6/d__14_ DECAP_INV_G11
XG12457 XI11_2/XI0/XI0_6/d_13_ XI11_2/XI0/XI0_6/d__13_ DECAP_INV_G11
XG12458 XI11_2/XI0/XI0_6/d_12_ XI11_2/XI0/XI0_6/d__12_ DECAP_INV_G11
XG12459 XI11_2/XI0/XI0_6/d_11_ XI11_2/XI0/XI0_6/d__11_ DECAP_INV_G11
XG12460 XI11_2/XI0/XI0_6/d_10_ XI11_2/XI0/XI0_6/d__10_ DECAP_INV_G11
XG12461 XI11_2/XI0/XI0_6/d_9_ XI11_2/XI0/XI0_6/d__9_ DECAP_INV_G11
XG12462 XI11_2/XI0/XI0_6/d_8_ XI11_2/XI0/XI0_6/d__8_ DECAP_INV_G11
XG12463 XI11_2/XI0/XI0_6/d_7_ XI11_2/XI0/XI0_6/d__7_ DECAP_INV_G11
XG12464 XI11_2/XI0/XI0_6/d_6_ XI11_2/XI0/XI0_6/d__6_ DECAP_INV_G11
XG12465 XI11_2/XI0/XI0_6/d_5_ XI11_2/XI0/XI0_6/d__5_ DECAP_INV_G11
XG12466 XI11_2/XI0/XI0_6/d_4_ XI11_2/XI0/XI0_6/d__4_ DECAP_INV_G11
XG12467 XI11_2/XI0/XI0_6/d_3_ XI11_2/XI0/XI0_6/d__3_ DECAP_INV_G11
XG12468 XI11_2/XI0/XI0_6/d_2_ XI11_2/XI0/XI0_6/d__2_ DECAP_INV_G11
XG12469 XI11_2/XI0/XI0_6/d_1_ XI11_2/XI0/XI0_6/d__1_ DECAP_INV_G11
XG12470 XI11_2/XI0/XI0_6/d_0_ XI11_2/XI0/XI0_6/d__0_ DECAP_INV_G11
XG12471 XI11_2/XI0/XI0_5/d__15_ XI11_2/XI0/XI0_5/d_15_ DECAP_INV_G11
XG12472 XI11_2/XI0/XI0_5/d__14_ XI11_2/XI0/XI0_5/d_14_ DECAP_INV_G11
XG12473 XI11_2/XI0/XI0_5/d__13_ XI11_2/XI0/XI0_5/d_13_ DECAP_INV_G11
XG12474 XI11_2/XI0/XI0_5/d__12_ XI11_2/XI0/XI0_5/d_12_ DECAP_INV_G11
XG12475 XI11_2/XI0/XI0_5/d__11_ XI11_2/XI0/XI0_5/d_11_ DECAP_INV_G11
XG12476 XI11_2/XI0/XI0_5/d__10_ XI11_2/XI0/XI0_5/d_10_ DECAP_INV_G11
XG12477 XI11_2/XI0/XI0_5/d__9_ XI11_2/XI0/XI0_5/d_9_ DECAP_INV_G11
XG12478 XI11_2/XI0/XI0_5/d__8_ XI11_2/XI0/XI0_5/d_8_ DECAP_INV_G11
XG12479 XI11_2/XI0/XI0_5/d__7_ XI11_2/XI0/XI0_5/d_7_ DECAP_INV_G11
XG12480 XI11_2/XI0/XI0_5/d__6_ XI11_2/XI0/XI0_5/d_6_ DECAP_INV_G11
XG12481 XI11_2/XI0/XI0_5/d__5_ XI11_2/XI0/XI0_5/d_5_ DECAP_INV_G11
XG12482 XI11_2/XI0/XI0_5/d__4_ XI11_2/XI0/XI0_5/d_4_ DECAP_INV_G11
XG12483 XI11_2/XI0/XI0_5/d__3_ XI11_2/XI0/XI0_5/d_3_ DECAP_INV_G11
XG12484 XI11_2/XI0/XI0_5/d__2_ XI11_2/XI0/XI0_5/d_2_ DECAP_INV_G11
XG12485 XI11_2/XI0/XI0_5/d__1_ XI11_2/XI0/XI0_5/d_1_ DECAP_INV_G11
XG12486 XI11_2/XI0/XI0_5/d__0_ XI11_2/XI0/XI0_5/d_0_ DECAP_INV_G11
XG12487 XI11_2/XI0/XI0_5/d_15_ XI11_2/XI0/XI0_5/d__15_ DECAP_INV_G11
XG12488 XI11_2/XI0/XI0_5/d_14_ XI11_2/XI0/XI0_5/d__14_ DECAP_INV_G11
XG12489 XI11_2/XI0/XI0_5/d_13_ XI11_2/XI0/XI0_5/d__13_ DECAP_INV_G11
XG12490 XI11_2/XI0/XI0_5/d_12_ XI11_2/XI0/XI0_5/d__12_ DECAP_INV_G11
XG12491 XI11_2/XI0/XI0_5/d_11_ XI11_2/XI0/XI0_5/d__11_ DECAP_INV_G11
XG12492 XI11_2/XI0/XI0_5/d_10_ XI11_2/XI0/XI0_5/d__10_ DECAP_INV_G11
XG12493 XI11_2/XI0/XI0_5/d_9_ XI11_2/XI0/XI0_5/d__9_ DECAP_INV_G11
XG12494 XI11_2/XI0/XI0_5/d_8_ XI11_2/XI0/XI0_5/d__8_ DECAP_INV_G11
XG12495 XI11_2/XI0/XI0_5/d_7_ XI11_2/XI0/XI0_5/d__7_ DECAP_INV_G11
XG12496 XI11_2/XI0/XI0_5/d_6_ XI11_2/XI0/XI0_5/d__6_ DECAP_INV_G11
XG12497 XI11_2/XI0/XI0_5/d_5_ XI11_2/XI0/XI0_5/d__5_ DECAP_INV_G11
XG12498 XI11_2/XI0/XI0_5/d_4_ XI11_2/XI0/XI0_5/d__4_ DECAP_INV_G11
XG12499 XI11_2/XI0/XI0_5/d_3_ XI11_2/XI0/XI0_5/d__3_ DECAP_INV_G11
XG12500 XI11_2/XI0/XI0_5/d_2_ XI11_2/XI0/XI0_5/d__2_ DECAP_INV_G11
XG12501 XI11_2/XI0/XI0_5/d_1_ XI11_2/XI0/XI0_5/d__1_ DECAP_INV_G11
XG12502 XI11_2/XI0/XI0_5/d_0_ XI11_2/XI0/XI0_5/d__0_ DECAP_INV_G11
XG12503 XI11_2/XI0/XI0_4/d__15_ XI11_2/XI0/XI0_4/d_15_ DECAP_INV_G11
XG12504 XI11_2/XI0/XI0_4/d__14_ XI11_2/XI0/XI0_4/d_14_ DECAP_INV_G11
XG12505 XI11_2/XI0/XI0_4/d__13_ XI11_2/XI0/XI0_4/d_13_ DECAP_INV_G11
XG12506 XI11_2/XI0/XI0_4/d__12_ XI11_2/XI0/XI0_4/d_12_ DECAP_INV_G11
XG12507 XI11_2/XI0/XI0_4/d__11_ XI11_2/XI0/XI0_4/d_11_ DECAP_INV_G11
XG12508 XI11_2/XI0/XI0_4/d__10_ XI11_2/XI0/XI0_4/d_10_ DECAP_INV_G11
XG12509 XI11_2/XI0/XI0_4/d__9_ XI11_2/XI0/XI0_4/d_9_ DECAP_INV_G11
XG12510 XI11_2/XI0/XI0_4/d__8_ XI11_2/XI0/XI0_4/d_8_ DECAP_INV_G11
XG12511 XI11_2/XI0/XI0_4/d__7_ XI11_2/XI0/XI0_4/d_7_ DECAP_INV_G11
XG12512 XI11_2/XI0/XI0_4/d__6_ XI11_2/XI0/XI0_4/d_6_ DECAP_INV_G11
XG12513 XI11_2/XI0/XI0_4/d__5_ XI11_2/XI0/XI0_4/d_5_ DECAP_INV_G11
XG12514 XI11_2/XI0/XI0_4/d__4_ XI11_2/XI0/XI0_4/d_4_ DECAP_INV_G11
XG12515 XI11_2/XI0/XI0_4/d__3_ XI11_2/XI0/XI0_4/d_3_ DECAP_INV_G11
XG12516 XI11_2/XI0/XI0_4/d__2_ XI11_2/XI0/XI0_4/d_2_ DECAP_INV_G11
XG12517 XI11_2/XI0/XI0_4/d__1_ XI11_2/XI0/XI0_4/d_1_ DECAP_INV_G11
XG12518 XI11_2/XI0/XI0_4/d__0_ XI11_2/XI0/XI0_4/d_0_ DECAP_INV_G11
XG12519 XI11_2/XI0/XI0_4/d_15_ XI11_2/XI0/XI0_4/d__15_ DECAP_INV_G11
XG12520 XI11_2/XI0/XI0_4/d_14_ XI11_2/XI0/XI0_4/d__14_ DECAP_INV_G11
XG12521 XI11_2/XI0/XI0_4/d_13_ XI11_2/XI0/XI0_4/d__13_ DECAP_INV_G11
XG12522 XI11_2/XI0/XI0_4/d_12_ XI11_2/XI0/XI0_4/d__12_ DECAP_INV_G11
XG12523 XI11_2/XI0/XI0_4/d_11_ XI11_2/XI0/XI0_4/d__11_ DECAP_INV_G11
XG12524 XI11_2/XI0/XI0_4/d_10_ XI11_2/XI0/XI0_4/d__10_ DECAP_INV_G11
XG12525 XI11_2/XI0/XI0_4/d_9_ XI11_2/XI0/XI0_4/d__9_ DECAP_INV_G11
XG12526 XI11_2/XI0/XI0_4/d_8_ XI11_2/XI0/XI0_4/d__8_ DECAP_INV_G11
XG12527 XI11_2/XI0/XI0_4/d_7_ XI11_2/XI0/XI0_4/d__7_ DECAP_INV_G11
XG12528 XI11_2/XI0/XI0_4/d_6_ XI11_2/XI0/XI0_4/d__6_ DECAP_INV_G11
XG12529 XI11_2/XI0/XI0_4/d_5_ XI11_2/XI0/XI0_4/d__5_ DECAP_INV_G11
XG12530 XI11_2/XI0/XI0_4/d_4_ XI11_2/XI0/XI0_4/d__4_ DECAP_INV_G11
XG12531 XI11_2/XI0/XI0_4/d_3_ XI11_2/XI0/XI0_4/d__3_ DECAP_INV_G11
XG12532 XI11_2/XI0/XI0_4/d_2_ XI11_2/XI0/XI0_4/d__2_ DECAP_INV_G11
XG12533 XI11_2/XI0/XI0_4/d_1_ XI11_2/XI0/XI0_4/d__1_ DECAP_INV_G11
XG12534 XI11_2/XI0/XI0_4/d_0_ XI11_2/XI0/XI0_4/d__0_ DECAP_INV_G11
XG12535 XI11_2/XI0/XI0_3/d__15_ XI11_2/XI0/XI0_3/d_15_ DECAP_INV_G11
XG12536 XI11_2/XI0/XI0_3/d__14_ XI11_2/XI0/XI0_3/d_14_ DECAP_INV_G11
XG12537 XI11_2/XI0/XI0_3/d__13_ XI11_2/XI0/XI0_3/d_13_ DECAP_INV_G11
XG12538 XI11_2/XI0/XI0_3/d__12_ XI11_2/XI0/XI0_3/d_12_ DECAP_INV_G11
XG12539 XI11_2/XI0/XI0_3/d__11_ XI11_2/XI0/XI0_3/d_11_ DECAP_INV_G11
XG12540 XI11_2/XI0/XI0_3/d__10_ XI11_2/XI0/XI0_3/d_10_ DECAP_INV_G11
XG12541 XI11_2/XI0/XI0_3/d__9_ XI11_2/XI0/XI0_3/d_9_ DECAP_INV_G11
XG12542 XI11_2/XI0/XI0_3/d__8_ XI11_2/XI0/XI0_3/d_8_ DECAP_INV_G11
XG12543 XI11_2/XI0/XI0_3/d__7_ XI11_2/XI0/XI0_3/d_7_ DECAP_INV_G11
XG12544 XI11_2/XI0/XI0_3/d__6_ XI11_2/XI0/XI0_3/d_6_ DECAP_INV_G11
XG12545 XI11_2/XI0/XI0_3/d__5_ XI11_2/XI0/XI0_3/d_5_ DECAP_INV_G11
XG12546 XI11_2/XI0/XI0_3/d__4_ XI11_2/XI0/XI0_3/d_4_ DECAP_INV_G11
XG12547 XI11_2/XI0/XI0_3/d__3_ XI11_2/XI0/XI0_3/d_3_ DECAP_INV_G11
XG12548 XI11_2/XI0/XI0_3/d__2_ XI11_2/XI0/XI0_3/d_2_ DECAP_INV_G11
XG12549 XI11_2/XI0/XI0_3/d__1_ XI11_2/XI0/XI0_3/d_1_ DECAP_INV_G11
XG12550 XI11_2/XI0/XI0_3/d__0_ XI11_2/XI0/XI0_3/d_0_ DECAP_INV_G11
XG12551 XI11_2/XI0/XI0_3/d_15_ XI11_2/XI0/XI0_3/d__15_ DECAP_INV_G11
XG12552 XI11_2/XI0/XI0_3/d_14_ XI11_2/XI0/XI0_3/d__14_ DECAP_INV_G11
XG12553 XI11_2/XI0/XI0_3/d_13_ XI11_2/XI0/XI0_3/d__13_ DECAP_INV_G11
XG12554 XI11_2/XI0/XI0_3/d_12_ XI11_2/XI0/XI0_3/d__12_ DECAP_INV_G11
XG12555 XI11_2/XI0/XI0_3/d_11_ XI11_2/XI0/XI0_3/d__11_ DECAP_INV_G11
XG12556 XI11_2/XI0/XI0_3/d_10_ XI11_2/XI0/XI0_3/d__10_ DECAP_INV_G11
XG12557 XI11_2/XI0/XI0_3/d_9_ XI11_2/XI0/XI0_3/d__9_ DECAP_INV_G11
XG12558 XI11_2/XI0/XI0_3/d_8_ XI11_2/XI0/XI0_3/d__8_ DECAP_INV_G11
XG12559 XI11_2/XI0/XI0_3/d_7_ XI11_2/XI0/XI0_3/d__7_ DECAP_INV_G11
XG12560 XI11_2/XI0/XI0_3/d_6_ XI11_2/XI0/XI0_3/d__6_ DECAP_INV_G11
XG12561 XI11_2/XI0/XI0_3/d_5_ XI11_2/XI0/XI0_3/d__5_ DECAP_INV_G11
XG12562 XI11_2/XI0/XI0_3/d_4_ XI11_2/XI0/XI0_3/d__4_ DECAP_INV_G11
XG12563 XI11_2/XI0/XI0_3/d_3_ XI11_2/XI0/XI0_3/d__3_ DECAP_INV_G11
XG12564 XI11_2/XI0/XI0_3/d_2_ XI11_2/XI0/XI0_3/d__2_ DECAP_INV_G11
XG12565 XI11_2/XI0/XI0_3/d_1_ XI11_2/XI0/XI0_3/d__1_ DECAP_INV_G11
XG12566 XI11_2/XI0/XI0_3/d_0_ XI11_2/XI0/XI0_3/d__0_ DECAP_INV_G11
XG12567 XI11_2/XI0/XI0_2/d__15_ XI11_2/XI0/XI0_2/d_15_ DECAP_INV_G11
XG12568 XI11_2/XI0/XI0_2/d__14_ XI11_2/XI0/XI0_2/d_14_ DECAP_INV_G11
XG12569 XI11_2/XI0/XI0_2/d__13_ XI11_2/XI0/XI0_2/d_13_ DECAP_INV_G11
XG12570 XI11_2/XI0/XI0_2/d__12_ XI11_2/XI0/XI0_2/d_12_ DECAP_INV_G11
XG12571 XI11_2/XI0/XI0_2/d__11_ XI11_2/XI0/XI0_2/d_11_ DECAP_INV_G11
XG12572 XI11_2/XI0/XI0_2/d__10_ XI11_2/XI0/XI0_2/d_10_ DECAP_INV_G11
XG12573 XI11_2/XI0/XI0_2/d__9_ XI11_2/XI0/XI0_2/d_9_ DECAP_INV_G11
XG12574 XI11_2/XI0/XI0_2/d__8_ XI11_2/XI0/XI0_2/d_8_ DECAP_INV_G11
XG12575 XI11_2/XI0/XI0_2/d__7_ XI11_2/XI0/XI0_2/d_7_ DECAP_INV_G11
XG12576 XI11_2/XI0/XI0_2/d__6_ XI11_2/XI0/XI0_2/d_6_ DECAP_INV_G11
XG12577 XI11_2/XI0/XI0_2/d__5_ XI11_2/XI0/XI0_2/d_5_ DECAP_INV_G11
XG12578 XI11_2/XI0/XI0_2/d__4_ XI11_2/XI0/XI0_2/d_4_ DECAP_INV_G11
XG12579 XI11_2/XI0/XI0_2/d__3_ XI11_2/XI0/XI0_2/d_3_ DECAP_INV_G11
XG12580 XI11_2/XI0/XI0_2/d__2_ XI11_2/XI0/XI0_2/d_2_ DECAP_INV_G11
XG12581 XI11_2/XI0/XI0_2/d__1_ XI11_2/XI0/XI0_2/d_1_ DECAP_INV_G11
XG12582 XI11_2/XI0/XI0_2/d__0_ XI11_2/XI0/XI0_2/d_0_ DECAP_INV_G11
XG12583 XI11_2/XI0/XI0_2/d_15_ XI11_2/XI0/XI0_2/d__15_ DECAP_INV_G11
XG12584 XI11_2/XI0/XI0_2/d_14_ XI11_2/XI0/XI0_2/d__14_ DECAP_INV_G11
XG12585 XI11_2/XI0/XI0_2/d_13_ XI11_2/XI0/XI0_2/d__13_ DECAP_INV_G11
XG12586 XI11_2/XI0/XI0_2/d_12_ XI11_2/XI0/XI0_2/d__12_ DECAP_INV_G11
XG12587 XI11_2/XI0/XI0_2/d_11_ XI11_2/XI0/XI0_2/d__11_ DECAP_INV_G11
XG12588 XI11_2/XI0/XI0_2/d_10_ XI11_2/XI0/XI0_2/d__10_ DECAP_INV_G11
XG12589 XI11_2/XI0/XI0_2/d_9_ XI11_2/XI0/XI0_2/d__9_ DECAP_INV_G11
XG12590 XI11_2/XI0/XI0_2/d_8_ XI11_2/XI0/XI0_2/d__8_ DECAP_INV_G11
XG12591 XI11_2/XI0/XI0_2/d_7_ XI11_2/XI0/XI0_2/d__7_ DECAP_INV_G11
XG12592 XI11_2/XI0/XI0_2/d_6_ XI11_2/XI0/XI0_2/d__6_ DECAP_INV_G11
XG12593 XI11_2/XI0/XI0_2/d_5_ XI11_2/XI0/XI0_2/d__5_ DECAP_INV_G11
XG12594 XI11_2/XI0/XI0_2/d_4_ XI11_2/XI0/XI0_2/d__4_ DECAP_INV_G11
XG12595 XI11_2/XI0/XI0_2/d_3_ XI11_2/XI0/XI0_2/d__3_ DECAP_INV_G11
XG12596 XI11_2/XI0/XI0_2/d_2_ XI11_2/XI0/XI0_2/d__2_ DECAP_INV_G11
XG12597 XI11_2/XI0/XI0_2/d_1_ XI11_2/XI0/XI0_2/d__1_ DECAP_INV_G11
XG12598 XI11_2/XI0/XI0_2/d_0_ XI11_2/XI0/XI0_2/d__0_ DECAP_INV_G11
XG12599 XI11_2/XI0/XI0_1/d__15_ XI11_2/XI0/XI0_1/d_15_ DECAP_INV_G11
XG12600 XI11_2/XI0/XI0_1/d__14_ XI11_2/XI0/XI0_1/d_14_ DECAP_INV_G11
XG12601 XI11_2/XI0/XI0_1/d__13_ XI11_2/XI0/XI0_1/d_13_ DECAP_INV_G11
XG12602 XI11_2/XI0/XI0_1/d__12_ XI11_2/XI0/XI0_1/d_12_ DECAP_INV_G11
XG12603 XI11_2/XI0/XI0_1/d__11_ XI11_2/XI0/XI0_1/d_11_ DECAP_INV_G11
XG12604 XI11_2/XI0/XI0_1/d__10_ XI11_2/XI0/XI0_1/d_10_ DECAP_INV_G11
XG12605 XI11_2/XI0/XI0_1/d__9_ XI11_2/XI0/XI0_1/d_9_ DECAP_INV_G11
XG12606 XI11_2/XI0/XI0_1/d__8_ XI11_2/XI0/XI0_1/d_8_ DECAP_INV_G11
XG12607 XI11_2/XI0/XI0_1/d__7_ XI11_2/XI0/XI0_1/d_7_ DECAP_INV_G11
XG12608 XI11_2/XI0/XI0_1/d__6_ XI11_2/XI0/XI0_1/d_6_ DECAP_INV_G11
XG12609 XI11_2/XI0/XI0_1/d__5_ XI11_2/XI0/XI0_1/d_5_ DECAP_INV_G11
XG12610 XI11_2/XI0/XI0_1/d__4_ XI11_2/XI0/XI0_1/d_4_ DECAP_INV_G11
XG12611 XI11_2/XI0/XI0_1/d__3_ XI11_2/XI0/XI0_1/d_3_ DECAP_INV_G11
XG12612 XI11_2/XI0/XI0_1/d__2_ XI11_2/XI0/XI0_1/d_2_ DECAP_INV_G11
XG12613 XI11_2/XI0/XI0_1/d__1_ XI11_2/XI0/XI0_1/d_1_ DECAP_INV_G11
XG12614 XI11_2/XI0/XI0_1/d__0_ XI11_2/XI0/XI0_1/d_0_ DECAP_INV_G11
XG12615 XI11_2/XI0/XI0_1/d_15_ XI11_2/XI0/XI0_1/d__15_ DECAP_INV_G11
XG12616 XI11_2/XI0/XI0_1/d_14_ XI11_2/XI0/XI0_1/d__14_ DECAP_INV_G11
XG12617 XI11_2/XI0/XI0_1/d_13_ XI11_2/XI0/XI0_1/d__13_ DECAP_INV_G11
XG12618 XI11_2/XI0/XI0_1/d_12_ XI11_2/XI0/XI0_1/d__12_ DECAP_INV_G11
XG12619 XI11_2/XI0/XI0_1/d_11_ XI11_2/XI0/XI0_1/d__11_ DECAP_INV_G11
XG12620 XI11_2/XI0/XI0_1/d_10_ XI11_2/XI0/XI0_1/d__10_ DECAP_INV_G11
XG12621 XI11_2/XI0/XI0_1/d_9_ XI11_2/XI0/XI0_1/d__9_ DECAP_INV_G11
XG12622 XI11_2/XI0/XI0_1/d_8_ XI11_2/XI0/XI0_1/d__8_ DECAP_INV_G11
XG12623 XI11_2/XI0/XI0_1/d_7_ XI11_2/XI0/XI0_1/d__7_ DECAP_INV_G11
XG12624 XI11_2/XI0/XI0_1/d_6_ XI11_2/XI0/XI0_1/d__6_ DECAP_INV_G11
XG12625 XI11_2/XI0/XI0_1/d_5_ XI11_2/XI0/XI0_1/d__5_ DECAP_INV_G11
XG12626 XI11_2/XI0/XI0_1/d_4_ XI11_2/XI0/XI0_1/d__4_ DECAP_INV_G11
XG12627 XI11_2/XI0/XI0_1/d_3_ XI11_2/XI0/XI0_1/d__3_ DECAP_INV_G11
XG12628 XI11_2/XI0/XI0_1/d_2_ XI11_2/XI0/XI0_1/d__2_ DECAP_INV_G11
XG12629 XI11_2/XI0/XI0_1/d_1_ XI11_2/XI0/XI0_1/d__1_ DECAP_INV_G11
XG12630 XI11_2/XI0/XI0_1/d_0_ XI11_2/XI0/XI0_1/d__0_ DECAP_INV_G11
XG12631 XI11_2/XI0/XI0_0/d__15_ XI11_2/XI0/XI0_0/d_15_ DECAP_INV_G11
XG12632 XI11_2/XI0/XI0_0/d__14_ XI11_2/XI0/XI0_0/d_14_ DECAP_INV_G11
XG12633 XI11_2/XI0/XI0_0/d__13_ XI11_2/XI0/XI0_0/d_13_ DECAP_INV_G11
XG12634 XI11_2/XI0/XI0_0/d__12_ XI11_2/XI0/XI0_0/d_12_ DECAP_INV_G11
XG12635 XI11_2/XI0/XI0_0/d__11_ XI11_2/XI0/XI0_0/d_11_ DECAP_INV_G11
XG12636 XI11_2/XI0/XI0_0/d__10_ XI11_2/XI0/XI0_0/d_10_ DECAP_INV_G11
XG12637 XI11_2/XI0/XI0_0/d__9_ XI11_2/XI0/XI0_0/d_9_ DECAP_INV_G11
XG12638 XI11_2/XI0/XI0_0/d__8_ XI11_2/XI0/XI0_0/d_8_ DECAP_INV_G11
XG12639 XI11_2/XI0/XI0_0/d__7_ XI11_2/XI0/XI0_0/d_7_ DECAP_INV_G11
XG12640 XI11_2/XI0/XI0_0/d__6_ XI11_2/XI0/XI0_0/d_6_ DECAP_INV_G11
XG12641 XI11_2/XI0/XI0_0/d__5_ XI11_2/XI0/XI0_0/d_5_ DECAP_INV_G11
XG12642 XI11_2/XI0/XI0_0/d__4_ XI11_2/XI0/XI0_0/d_4_ DECAP_INV_G11
XG12643 XI11_2/XI0/XI0_0/d__3_ XI11_2/XI0/XI0_0/d_3_ DECAP_INV_G11
XG12644 XI11_2/XI0/XI0_0/d__2_ XI11_2/XI0/XI0_0/d_2_ DECAP_INV_G11
XG12645 XI11_2/XI0/XI0_0/d__1_ XI11_2/XI0/XI0_0/d_1_ DECAP_INV_G11
XG12646 XI11_2/XI0/XI0_0/d__0_ XI11_2/XI0/XI0_0/d_0_ DECAP_INV_G11
XG12647 XI11_2/XI0/XI0_0/d_15_ XI11_2/XI0/XI0_0/d__15_ DECAP_INV_G11
XG12648 XI11_2/XI0/XI0_0/d_14_ XI11_2/XI0/XI0_0/d__14_ DECAP_INV_G11
XG12649 XI11_2/XI0/XI0_0/d_13_ XI11_2/XI0/XI0_0/d__13_ DECAP_INV_G11
XG12650 XI11_2/XI0/XI0_0/d_12_ XI11_2/XI0/XI0_0/d__12_ DECAP_INV_G11
XG12651 XI11_2/XI0/XI0_0/d_11_ XI11_2/XI0/XI0_0/d__11_ DECAP_INV_G11
XG12652 XI11_2/XI0/XI0_0/d_10_ XI11_2/XI0/XI0_0/d__10_ DECAP_INV_G11
XG12653 XI11_2/XI0/XI0_0/d_9_ XI11_2/XI0/XI0_0/d__9_ DECAP_INV_G11
XG12654 XI11_2/XI0/XI0_0/d_8_ XI11_2/XI0/XI0_0/d__8_ DECAP_INV_G11
XG12655 XI11_2/XI0/XI0_0/d_7_ XI11_2/XI0/XI0_0/d__7_ DECAP_INV_G11
XG12656 XI11_2/XI0/XI0_0/d_6_ XI11_2/XI0/XI0_0/d__6_ DECAP_INV_G11
XG12657 XI11_2/XI0/XI0_0/d_5_ XI11_2/XI0/XI0_0/d__5_ DECAP_INV_G11
XG12658 XI11_2/XI0/XI0_0/d_4_ XI11_2/XI0/XI0_0/d__4_ DECAP_INV_G11
XG12659 XI11_2/XI0/XI0_0/d_3_ XI11_2/XI0/XI0_0/d__3_ DECAP_INV_G11
XG12660 XI11_2/XI0/XI0_0/d_2_ XI11_2/XI0/XI0_0/d__2_ DECAP_INV_G11
XG12661 XI11_2/XI0/XI0_0/d_1_ XI11_2/XI0/XI0_0/d__1_ DECAP_INV_G11
XG12662 XI11_2/XI0/XI0_0/d_0_ XI11_2/XI0/XI0_0/d__0_ DECAP_INV_G11
XG12663 XI11_1/XI3/net17 XI11_1/XI3/net5 DECAP_INV_G7
XG12664 XI11_1/XI3/net5 XI11_1/preck DECAP_INV_G8
XG12665 sck_bar XI11_1/XI3/net018 DECAP_INV_G9
XG12666 XI11_1/XI3/net018 XI11_1/XI3/net012 DECAP_INV_G9
XG12667 XI11_1/XI3/net014 XI11_1/XI3/net7 DECAP_INV_G9
XG12668 XI11_1/XI3/net012 XI11_1/XI3/net014 DECAP_INV_G9
XG12669 XI11_1/XI4/net063 XI11_1/XI4/net0112 DECAP_INV_G10
XG12670 XI11_1/XI4/net26 XI11_1/XI4/net089 DECAP_INV_G10
XG12671 XI11_1/XI4/data_out XI11_1/XI4/data_out_ DECAP_INV_G10
XG12672 XI11_1/XI4/net20 XI11_1/XI4/net0103 DECAP_INV_G10
XG12673 XI11_1/net12 XI11_1/XI4/net32 DECAP_INV_G7
XG12674 XI11_1/net9 XI11_1/XI4/net52 DECAP_INV_G7
XG12675 XI11_1/XI4/data_out_ XI11_1/XI4/data_out DECAP_INV_G10
XG12676 XI11_1/XI0/XI0_63/d__15_ XI11_1/XI0/XI0_63/d_15_ DECAP_INV_G11
XG12677 XI11_1/XI0/XI0_63/d__14_ XI11_1/XI0/XI0_63/d_14_ DECAP_INV_G11
XG12678 XI11_1/XI0/XI0_63/d__13_ XI11_1/XI0/XI0_63/d_13_ DECAP_INV_G11
XG12679 XI11_1/XI0/XI0_63/d__12_ XI11_1/XI0/XI0_63/d_12_ DECAP_INV_G11
XG12680 XI11_1/XI0/XI0_63/d__11_ XI11_1/XI0/XI0_63/d_11_ DECAP_INV_G11
XG12681 XI11_1/XI0/XI0_63/d__10_ XI11_1/XI0/XI0_63/d_10_ DECAP_INV_G11
XG12682 XI11_1/XI0/XI0_63/d__9_ XI11_1/XI0/XI0_63/d_9_ DECAP_INV_G11
XG12683 XI11_1/XI0/XI0_63/d__8_ XI11_1/XI0/XI0_63/d_8_ DECAP_INV_G11
XG12684 XI11_1/XI0/XI0_63/d__7_ XI11_1/XI0/XI0_63/d_7_ DECAP_INV_G11
XG12685 XI11_1/XI0/XI0_63/d__6_ XI11_1/XI0/XI0_63/d_6_ DECAP_INV_G11
XG12686 XI11_1/XI0/XI0_63/d__5_ XI11_1/XI0/XI0_63/d_5_ DECAP_INV_G11
XG12687 XI11_1/XI0/XI0_63/d__4_ XI11_1/XI0/XI0_63/d_4_ DECAP_INV_G11
XG12688 XI11_1/XI0/XI0_63/d__3_ XI11_1/XI0/XI0_63/d_3_ DECAP_INV_G11
XG12689 XI11_1/XI0/XI0_63/d__2_ XI11_1/XI0/XI0_63/d_2_ DECAP_INV_G11
XG12690 XI11_1/XI0/XI0_63/d__1_ XI11_1/XI0/XI0_63/d_1_ DECAP_INV_G11
XG12691 XI11_1/XI0/XI0_63/d__0_ XI11_1/XI0/XI0_63/d_0_ DECAP_INV_G11
XG12692 XI11_1/XI0/XI0_63/d_15_ XI11_1/XI0/XI0_63/d__15_ DECAP_INV_G11
XG12693 XI11_1/XI0/XI0_63/d_14_ XI11_1/XI0/XI0_63/d__14_ DECAP_INV_G11
XG12694 XI11_1/XI0/XI0_63/d_13_ XI11_1/XI0/XI0_63/d__13_ DECAP_INV_G11
XG12695 XI11_1/XI0/XI0_63/d_12_ XI11_1/XI0/XI0_63/d__12_ DECAP_INV_G11
XG12696 XI11_1/XI0/XI0_63/d_11_ XI11_1/XI0/XI0_63/d__11_ DECAP_INV_G11
XG12697 XI11_1/XI0/XI0_63/d_10_ XI11_1/XI0/XI0_63/d__10_ DECAP_INV_G11
XG12698 XI11_1/XI0/XI0_63/d_9_ XI11_1/XI0/XI0_63/d__9_ DECAP_INV_G11
XG12699 XI11_1/XI0/XI0_63/d_8_ XI11_1/XI0/XI0_63/d__8_ DECAP_INV_G11
XG12700 XI11_1/XI0/XI0_63/d_7_ XI11_1/XI0/XI0_63/d__7_ DECAP_INV_G11
XG12701 XI11_1/XI0/XI0_63/d_6_ XI11_1/XI0/XI0_63/d__6_ DECAP_INV_G11
XG12702 XI11_1/XI0/XI0_63/d_5_ XI11_1/XI0/XI0_63/d__5_ DECAP_INV_G11
XG12703 XI11_1/XI0/XI0_63/d_4_ XI11_1/XI0/XI0_63/d__4_ DECAP_INV_G11
XG12704 XI11_1/XI0/XI0_63/d_3_ XI11_1/XI0/XI0_63/d__3_ DECAP_INV_G11
XG12705 XI11_1/XI0/XI0_63/d_2_ XI11_1/XI0/XI0_63/d__2_ DECAP_INV_G11
XG12706 XI11_1/XI0/XI0_63/d_1_ XI11_1/XI0/XI0_63/d__1_ DECAP_INV_G11
XG12707 XI11_1/XI0/XI0_63/d_0_ XI11_1/XI0/XI0_63/d__0_ DECAP_INV_G11
XG12708 XI11_1/XI0/XI0_62/d__15_ XI11_1/XI0/XI0_62/d_15_ DECAP_INV_G11
XG12709 XI11_1/XI0/XI0_62/d__14_ XI11_1/XI0/XI0_62/d_14_ DECAP_INV_G11
XG12710 XI11_1/XI0/XI0_62/d__13_ XI11_1/XI0/XI0_62/d_13_ DECAP_INV_G11
XG12711 XI11_1/XI0/XI0_62/d__12_ XI11_1/XI0/XI0_62/d_12_ DECAP_INV_G11
XG12712 XI11_1/XI0/XI0_62/d__11_ XI11_1/XI0/XI0_62/d_11_ DECAP_INV_G11
XG12713 XI11_1/XI0/XI0_62/d__10_ XI11_1/XI0/XI0_62/d_10_ DECAP_INV_G11
XG12714 XI11_1/XI0/XI0_62/d__9_ XI11_1/XI0/XI0_62/d_9_ DECAP_INV_G11
XG12715 XI11_1/XI0/XI0_62/d__8_ XI11_1/XI0/XI0_62/d_8_ DECAP_INV_G11
XG12716 XI11_1/XI0/XI0_62/d__7_ XI11_1/XI0/XI0_62/d_7_ DECAP_INV_G11
XG12717 XI11_1/XI0/XI0_62/d__6_ XI11_1/XI0/XI0_62/d_6_ DECAP_INV_G11
XG12718 XI11_1/XI0/XI0_62/d__5_ XI11_1/XI0/XI0_62/d_5_ DECAP_INV_G11
XG12719 XI11_1/XI0/XI0_62/d__4_ XI11_1/XI0/XI0_62/d_4_ DECAP_INV_G11
XG12720 XI11_1/XI0/XI0_62/d__3_ XI11_1/XI0/XI0_62/d_3_ DECAP_INV_G11
XG12721 XI11_1/XI0/XI0_62/d__2_ XI11_1/XI0/XI0_62/d_2_ DECAP_INV_G11
XG12722 XI11_1/XI0/XI0_62/d__1_ XI11_1/XI0/XI0_62/d_1_ DECAP_INV_G11
XG12723 XI11_1/XI0/XI0_62/d__0_ XI11_1/XI0/XI0_62/d_0_ DECAP_INV_G11
XG12724 XI11_1/XI0/XI0_62/d_15_ XI11_1/XI0/XI0_62/d__15_ DECAP_INV_G11
XG12725 XI11_1/XI0/XI0_62/d_14_ XI11_1/XI0/XI0_62/d__14_ DECAP_INV_G11
XG12726 XI11_1/XI0/XI0_62/d_13_ XI11_1/XI0/XI0_62/d__13_ DECAP_INV_G11
XG12727 XI11_1/XI0/XI0_62/d_12_ XI11_1/XI0/XI0_62/d__12_ DECAP_INV_G11
XG12728 XI11_1/XI0/XI0_62/d_11_ XI11_1/XI0/XI0_62/d__11_ DECAP_INV_G11
XG12729 XI11_1/XI0/XI0_62/d_10_ XI11_1/XI0/XI0_62/d__10_ DECAP_INV_G11
XG12730 XI11_1/XI0/XI0_62/d_9_ XI11_1/XI0/XI0_62/d__9_ DECAP_INV_G11
XG12731 XI11_1/XI0/XI0_62/d_8_ XI11_1/XI0/XI0_62/d__8_ DECAP_INV_G11
XG12732 XI11_1/XI0/XI0_62/d_7_ XI11_1/XI0/XI0_62/d__7_ DECAP_INV_G11
XG12733 XI11_1/XI0/XI0_62/d_6_ XI11_1/XI0/XI0_62/d__6_ DECAP_INV_G11
XG12734 XI11_1/XI0/XI0_62/d_5_ XI11_1/XI0/XI0_62/d__5_ DECAP_INV_G11
XG12735 XI11_1/XI0/XI0_62/d_4_ XI11_1/XI0/XI0_62/d__4_ DECAP_INV_G11
XG12736 XI11_1/XI0/XI0_62/d_3_ XI11_1/XI0/XI0_62/d__3_ DECAP_INV_G11
XG12737 XI11_1/XI0/XI0_62/d_2_ XI11_1/XI0/XI0_62/d__2_ DECAP_INV_G11
XG12738 XI11_1/XI0/XI0_62/d_1_ XI11_1/XI0/XI0_62/d__1_ DECAP_INV_G11
XG12739 XI11_1/XI0/XI0_62/d_0_ XI11_1/XI0/XI0_62/d__0_ DECAP_INV_G11
XG12740 XI11_1/XI0/XI0_61/d__15_ XI11_1/XI0/XI0_61/d_15_ DECAP_INV_G11
XG12741 XI11_1/XI0/XI0_61/d__14_ XI11_1/XI0/XI0_61/d_14_ DECAP_INV_G11
XG12742 XI11_1/XI0/XI0_61/d__13_ XI11_1/XI0/XI0_61/d_13_ DECAP_INV_G11
XG12743 XI11_1/XI0/XI0_61/d__12_ XI11_1/XI0/XI0_61/d_12_ DECAP_INV_G11
XG12744 XI11_1/XI0/XI0_61/d__11_ XI11_1/XI0/XI0_61/d_11_ DECAP_INV_G11
XG12745 XI11_1/XI0/XI0_61/d__10_ XI11_1/XI0/XI0_61/d_10_ DECAP_INV_G11
XG12746 XI11_1/XI0/XI0_61/d__9_ XI11_1/XI0/XI0_61/d_9_ DECAP_INV_G11
XG12747 XI11_1/XI0/XI0_61/d__8_ XI11_1/XI0/XI0_61/d_8_ DECAP_INV_G11
XG12748 XI11_1/XI0/XI0_61/d__7_ XI11_1/XI0/XI0_61/d_7_ DECAP_INV_G11
XG12749 XI11_1/XI0/XI0_61/d__6_ XI11_1/XI0/XI0_61/d_6_ DECAP_INV_G11
XG12750 XI11_1/XI0/XI0_61/d__5_ XI11_1/XI0/XI0_61/d_5_ DECAP_INV_G11
XG12751 XI11_1/XI0/XI0_61/d__4_ XI11_1/XI0/XI0_61/d_4_ DECAP_INV_G11
XG12752 XI11_1/XI0/XI0_61/d__3_ XI11_1/XI0/XI0_61/d_3_ DECAP_INV_G11
XG12753 XI11_1/XI0/XI0_61/d__2_ XI11_1/XI0/XI0_61/d_2_ DECAP_INV_G11
XG12754 XI11_1/XI0/XI0_61/d__1_ XI11_1/XI0/XI0_61/d_1_ DECAP_INV_G11
XG12755 XI11_1/XI0/XI0_61/d__0_ XI11_1/XI0/XI0_61/d_0_ DECAP_INV_G11
XG12756 XI11_1/XI0/XI0_61/d_15_ XI11_1/XI0/XI0_61/d__15_ DECAP_INV_G11
XG12757 XI11_1/XI0/XI0_61/d_14_ XI11_1/XI0/XI0_61/d__14_ DECAP_INV_G11
XG12758 XI11_1/XI0/XI0_61/d_13_ XI11_1/XI0/XI0_61/d__13_ DECAP_INV_G11
XG12759 XI11_1/XI0/XI0_61/d_12_ XI11_1/XI0/XI0_61/d__12_ DECAP_INV_G11
XG12760 XI11_1/XI0/XI0_61/d_11_ XI11_1/XI0/XI0_61/d__11_ DECAP_INV_G11
XG12761 XI11_1/XI0/XI0_61/d_10_ XI11_1/XI0/XI0_61/d__10_ DECAP_INV_G11
XG12762 XI11_1/XI0/XI0_61/d_9_ XI11_1/XI0/XI0_61/d__9_ DECAP_INV_G11
XG12763 XI11_1/XI0/XI0_61/d_8_ XI11_1/XI0/XI0_61/d__8_ DECAP_INV_G11
XG12764 XI11_1/XI0/XI0_61/d_7_ XI11_1/XI0/XI0_61/d__7_ DECAP_INV_G11
XG12765 XI11_1/XI0/XI0_61/d_6_ XI11_1/XI0/XI0_61/d__6_ DECAP_INV_G11
XG12766 XI11_1/XI0/XI0_61/d_5_ XI11_1/XI0/XI0_61/d__5_ DECAP_INV_G11
XG12767 XI11_1/XI0/XI0_61/d_4_ XI11_1/XI0/XI0_61/d__4_ DECAP_INV_G11
XG12768 XI11_1/XI0/XI0_61/d_3_ XI11_1/XI0/XI0_61/d__3_ DECAP_INV_G11
XG12769 XI11_1/XI0/XI0_61/d_2_ XI11_1/XI0/XI0_61/d__2_ DECAP_INV_G11
XG12770 XI11_1/XI0/XI0_61/d_1_ XI11_1/XI0/XI0_61/d__1_ DECAP_INV_G11
XG12771 XI11_1/XI0/XI0_61/d_0_ XI11_1/XI0/XI0_61/d__0_ DECAP_INV_G11
XG12772 XI11_1/XI0/XI0_60/d__15_ XI11_1/XI0/XI0_60/d_15_ DECAP_INV_G11
XG12773 XI11_1/XI0/XI0_60/d__14_ XI11_1/XI0/XI0_60/d_14_ DECAP_INV_G11
XG12774 XI11_1/XI0/XI0_60/d__13_ XI11_1/XI0/XI0_60/d_13_ DECAP_INV_G11
XG12775 XI11_1/XI0/XI0_60/d__12_ XI11_1/XI0/XI0_60/d_12_ DECAP_INV_G11
XG12776 XI11_1/XI0/XI0_60/d__11_ XI11_1/XI0/XI0_60/d_11_ DECAP_INV_G11
XG12777 XI11_1/XI0/XI0_60/d__10_ XI11_1/XI0/XI0_60/d_10_ DECAP_INV_G11
XG12778 XI11_1/XI0/XI0_60/d__9_ XI11_1/XI0/XI0_60/d_9_ DECAP_INV_G11
XG12779 XI11_1/XI0/XI0_60/d__8_ XI11_1/XI0/XI0_60/d_8_ DECAP_INV_G11
XG12780 XI11_1/XI0/XI0_60/d__7_ XI11_1/XI0/XI0_60/d_7_ DECAP_INV_G11
XG12781 XI11_1/XI0/XI0_60/d__6_ XI11_1/XI0/XI0_60/d_6_ DECAP_INV_G11
XG12782 XI11_1/XI0/XI0_60/d__5_ XI11_1/XI0/XI0_60/d_5_ DECAP_INV_G11
XG12783 XI11_1/XI0/XI0_60/d__4_ XI11_1/XI0/XI0_60/d_4_ DECAP_INV_G11
XG12784 XI11_1/XI0/XI0_60/d__3_ XI11_1/XI0/XI0_60/d_3_ DECAP_INV_G11
XG12785 XI11_1/XI0/XI0_60/d__2_ XI11_1/XI0/XI0_60/d_2_ DECAP_INV_G11
XG12786 XI11_1/XI0/XI0_60/d__1_ XI11_1/XI0/XI0_60/d_1_ DECAP_INV_G11
XG12787 XI11_1/XI0/XI0_60/d__0_ XI11_1/XI0/XI0_60/d_0_ DECAP_INV_G11
XG12788 XI11_1/XI0/XI0_60/d_15_ XI11_1/XI0/XI0_60/d__15_ DECAP_INV_G11
XG12789 XI11_1/XI0/XI0_60/d_14_ XI11_1/XI0/XI0_60/d__14_ DECAP_INV_G11
XG12790 XI11_1/XI0/XI0_60/d_13_ XI11_1/XI0/XI0_60/d__13_ DECAP_INV_G11
XG12791 XI11_1/XI0/XI0_60/d_12_ XI11_1/XI0/XI0_60/d__12_ DECAP_INV_G11
XG12792 XI11_1/XI0/XI0_60/d_11_ XI11_1/XI0/XI0_60/d__11_ DECAP_INV_G11
XG12793 XI11_1/XI0/XI0_60/d_10_ XI11_1/XI0/XI0_60/d__10_ DECAP_INV_G11
XG12794 XI11_1/XI0/XI0_60/d_9_ XI11_1/XI0/XI0_60/d__9_ DECAP_INV_G11
XG12795 XI11_1/XI0/XI0_60/d_8_ XI11_1/XI0/XI0_60/d__8_ DECAP_INV_G11
XG12796 XI11_1/XI0/XI0_60/d_7_ XI11_1/XI0/XI0_60/d__7_ DECAP_INV_G11
XG12797 XI11_1/XI0/XI0_60/d_6_ XI11_1/XI0/XI0_60/d__6_ DECAP_INV_G11
XG12798 XI11_1/XI0/XI0_60/d_5_ XI11_1/XI0/XI0_60/d__5_ DECAP_INV_G11
XG12799 XI11_1/XI0/XI0_60/d_4_ XI11_1/XI0/XI0_60/d__4_ DECAP_INV_G11
XG12800 XI11_1/XI0/XI0_60/d_3_ XI11_1/XI0/XI0_60/d__3_ DECAP_INV_G11
XG12801 XI11_1/XI0/XI0_60/d_2_ XI11_1/XI0/XI0_60/d__2_ DECAP_INV_G11
XG12802 XI11_1/XI0/XI0_60/d_1_ XI11_1/XI0/XI0_60/d__1_ DECAP_INV_G11
XG12803 XI11_1/XI0/XI0_60/d_0_ XI11_1/XI0/XI0_60/d__0_ DECAP_INV_G11
XG12804 XI11_1/XI0/XI0_59/d__15_ XI11_1/XI0/XI0_59/d_15_ DECAP_INV_G11
XG12805 XI11_1/XI0/XI0_59/d__14_ XI11_1/XI0/XI0_59/d_14_ DECAP_INV_G11
XG12806 XI11_1/XI0/XI0_59/d__13_ XI11_1/XI0/XI0_59/d_13_ DECAP_INV_G11
XG12807 XI11_1/XI0/XI0_59/d__12_ XI11_1/XI0/XI0_59/d_12_ DECAP_INV_G11
XG12808 XI11_1/XI0/XI0_59/d__11_ XI11_1/XI0/XI0_59/d_11_ DECAP_INV_G11
XG12809 XI11_1/XI0/XI0_59/d__10_ XI11_1/XI0/XI0_59/d_10_ DECAP_INV_G11
XG12810 XI11_1/XI0/XI0_59/d__9_ XI11_1/XI0/XI0_59/d_9_ DECAP_INV_G11
XG12811 XI11_1/XI0/XI0_59/d__8_ XI11_1/XI0/XI0_59/d_8_ DECAP_INV_G11
XG12812 XI11_1/XI0/XI0_59/d__7_ XI11_1/XI0/XI0_59/d_7_ DECAP_INV_G11
XG12813 XI11_1/XI0/XI0_59/d__6_ XI11_1/XI0/XI0_59/d_6_ DECAP_INV_G11
XG12814 XI11_1/XI0/XI0_59/d__5_ XI11_1/XI0/XI0_59/d_5_ DECAP_INV_G11
XG12815 XI11_1/XI0/XI0_59/d__4_ XI11_1/XI0/XI0_59/d_4_ DECAP_INV_G11
XG12816 XI11_1/XI0/XI0_59/d__3_ XI11_1/XI0/XI0_59/d_3_ DECAP_INV_G11
XG12817 XI11_1/XI0/XI0_59/d__2_ XI11_1/XI0/XI0_59/d_2_ DECAP_INV_G11
XG12818 XI11_1/XI0/XI0_59/d__1_ XI11_1/XI0/XI0_59/d_1_ DECAP_INV_G11
XG12819 XI11_1/XI0/XI0_59/d__0_ XI11_1/XI0/XI0_59/d_0_ DECAP_INV_G11
XG12820 XI11_1/XI0/XI0_59/d_15_ XI11_1/XI0/XI0_59/d__15_ DECAP_INV_G11
XG12821 XI11_1/XI0/XI0_59/d_14_ XI11_1/XI0/XI0_59/d__14_ DECAP_INV_G11
XG12822 XI11_1/XI0/XI0_59/d_13_ XI11_1/XI0/XI0_59/d__13_ DECAP_INV_G11
XG12823 XI11_1/XI0/XI0_59/d_12_ XI11_1/XI0/XI0_59/d__12_ DECAP_INV_G11
XG12824 XI11_1/XI0/XI0_59/d_11_ XI11_1/XI0/XI0_59/d__11_ DECAP_INV_G11
XG12825 XI11_1/XI0/XI0_59/d_10_ XI11_1/XI0/XI0_59/d__10_ DECAP_INV_G11
XG12826 XI11_1/XI0/XI0_59/d_9_ XI11_1/XI0/XI0_59/d__9_ DECAP_INV_G11
XG12827 XI11_1/XI0/XI0_59/d_8_ XI11_1/XI0/XI0_59/d__8_ DECAP_INV_G11
XG12828 XI11_1/XI0/XI0_59/d_7_ XI11_1/XI0/XI0_59/d__7_ DECAP_INV_G11
XG12829 XI11_1/XI0/XI0_59/d_6_ XI11_1/XI0/XI0_59/d__6_ DECAP_INV_G11
XG12830 XI11_1/XI0/XI0_59/d_5_ XI11_1/XI0/XI0_59/d__5_ DECAP_INV_G11
XG12831 XI11_1/XI0/XI0_59/d_4_ XI11_1/XI0/XI0_59/d__4_ DECAP_INV_G11
XG12832 XI11_1/XI0/XI0_59/d_3_ XI11_1/XI0/XI0_59/d__3_ DECAP_INV_G11
XG12833 XI11_1/XI0/XI0_59/d_2_ XI11_1/XI0/XI0_59/d__2_ DECAP_INV_G11
XG12834 XI11_1/XI0/XI0_59/d_1_ XI11_1/XI0/XI0_59/d__1_ DECAP_INV_G11
XG12835 XI11_1/XI0/XI0_59/d_0_ XI11_1/XI0/XI0_59/d__0_ DECAP_INV_G11
XG12836 XI11_1/XI0/XI0_58/d__15_ XI11_1/XI0/XI0_58/d_15_ DECAP_INV_G11
XG12837 XI11_1/XI0/XI0_58/d__14_ XI11_1/XI0/XI0_58/d_14_ DECAP_INV_G11
XG12838 XI11_1/XI0/XI0_58/d__13_ XI11_1/XI0/XI0_58/d_13_ DECAP_INV_G11
XG12839 XI11_1/XI0/XI0_58/d__12_ XI11_1/XI0/XI0_58/d_12_ DECAP_INV_G11
XG12840 XI11_1/XI0/XI0_58/d__11_ XI11_1/XI0/XI0_58/d_11_ DECAP_INV_G11
XG12841 XI11_1/XI0/XI0_58/d__10_ XI11_1/XI0/XI0_58/d_10_ DECAP_INV_G11
XG12842 XI11_1/XI0/XI0_58/d__9_ XI11_1/XI0/XI0_58/d_9_ DECAP_INV_G11
XG12843 XI11_1/XI0/XI0_58/d__8_ XI11_1/XI0/XI0_58/d_8_ DECAP_INV_G11
XG12844 XI11_1/XI0/XI0_58/d__7_ XI11_1/XI0/XI0_58/d_7_ DECAP_INV_G11
XG12845 XI11_1/XI0/XI0_58/d__6_ XI11_1/XI0/XI0_58/d_6_ DECAP_INV_G11
XG12846 XI11_1/XI0/XI0_58/d__5_ XI11_1/XI0/XI0_58/d_5_ DECAP_INV_G11
XG12847 XI11_1/XI0/XI0_58/d__4_ XI11_1/XI0/XI0_58/d_4_ DECAP_INV_G11
XG12848 XI11_1/XI0/XI0_58/d__3_ XI11_1/XI0/XI0_58/d_3_ DECAP_INV_G11
XG12849 XI11_1/XI0/XI0_58/d__2_ XI11_1/XI0/XI0_58/d_2_ DECAP_INV_G11
XG12850 XI11_1/XI0/XI0_58/d__1_ XI11_1/XI0/XI0_58/d_1_ DECAP_INV_G11
XG12851 XI11_1/XI0/XI0_58/d__0_ XI11_1/XI0/XI0_58/d_0_ DECAP_INV_G11
XG12852 XI11_1/XI0/XI0_58/d_15_ XI11_1/XI0/XI0_58/d__15_ DECAP_INV_G11
XG12853 XI11_1/XI0/XI0_58/d_14_ XI11_1/XI0/XI0_58/d__14_ DECAP_INV_G11
XG12854 XI11_1/XI0/XI0_58/d_13_ XI11_1/XI0/XI0_58/d__13_ DECAP_INV_G11
XG12855 XI11_1/XI0/XI0_58/d_12_ XI11_1/XI0/XI0_58/d__12_ DECAP_INV_G11
XG12856 XI11_1/XI0/XI0_58/d_11_ XI11_1/XI0/XI0_58/d__11_ DECAP_INV_G11
XG12857 XI11_1/XI0/XI0_58/d_10_ XI11_1/XI0/XI0_58/d__10_ DECAP_INV_G11
XG12858 XI11_1/XI0/XI0_58/d_9_ XI11_1/XI0/XI0_58/d__9_ DECAP_INV_G11
XG12859 XI11_1/XI0/XI0_58/d_8_ XI11_1/XI0/XI0_58/d__8_ DECAP_INV_G11
XG12860 XI11_1/XI0/XI0_58/d_7_ XI11_1/XI0/XI0_58/d__7_ DECAP_INV_G11
XG12861 XI11_1/XI0/XI0_58/d_6_ XI11_1/XI0/XI0_58/d__6_ DECAP_INV_G11
XG12862 XI11_1/XI0/XI0_58/d_5_ XI11_1/XI0/XI0_58/d__5_ DECAP_INV_G11
XG12863 XI11_1/XI0/XI0_58/d_4_ XI11_1/XI0/XI0_58/d__4_ DECAP_INV_G11
XG12864 XI11_1/XI0/XI0_58/d_3_ XI11_1/XI0/XI0_58/d__3_ DECAP_INV_G11
XG12865 XI11_1/XI0/XI0_58/d_2_ XI11_1/XI0/XI0_58/d__2_ DECAP_INV_G11
XG12866 XI11_1/XI0/XI0_58/d_1_ XI11_1/XI0/XI0_58/d__1_ DECAP_INV_G11
XG12867 XI11_1/XI0/XI0_58/d_0_ XI11_1/XI0/XI0_58/d__0_ DECAP_INV_G11
XG12868 XI11_1/XI0/XI0_57/d__15_ XI11_1/XI0/XI0_57/d_15_ DECAP_INV_G11
XG12869 XI11_1/XI0/XI0_57/d__14_ XI11_1/XI0/XI0_57/d_14_ DECAP_INV_G11
XG12870 XI11_1/XI0/XI0_57/d__13_ XI11_1/XI0/XI0_57/d_13_ DECAP_INV_G11
XG12871 XI11_1/XI0/XI0_57/d__12_ XI11_1/XI0/XI0_57/d_12_ DECAP_INV_G11
XG12872 XI11_1/XI0/XI0_57/d__11_ XI11_1/XI0/XI0_57/d_11_ DECAP_INV_G11
XG12873 XI11_1/XI0/XI0_57/d__10_ XI11_1/XI0/XI0_57/d_10_ DECAP_INV_G11
XG12874 XI11_1/XI0/XI0_57/d__9_ XI11_1/XI0/XI0_57/d_9_ DECAP_INV_G11
XG12875 XI11_1/XI0/XI0_57/d__8_ XI11_1/XI0/XI0_57/d_8_ DECAP_INV_G11
XG12876 XI11_1/XI0/XI0_57/d__7_ XI11_1/XI0/XI0_57/d_7_ DECAP_INV_G11
XG12877 XI11_1/XI0/XI0_57/d__6_ XI11_1/XI0/XI0_57/d_6_ DECAP_INV_G11
XG12878 XI11_1/XI0/XI0_57/d__5_ XI11_1/XI0/XI0_57/d_5_ DECAP_INV_G11
XG12879 XI11_1/XI0/XI0_57/d__4_ XI11_1/XI0/XI0_57/d_4_ DECAP_INV_G11
XG12880 XI11_1/XI0/XI0_57/d__3_ XI11_1/XI0/XI0_57/d_3_ DECAP_INV_G11
XG12881 XI11_1/XI0/XI0_57/d__2_ XI11_1/XI0/XI0_57/d_2_ DECAP_INV_G11
XG12882 XI11_1/XI0/XI0_57/d__1_ XI11_1/XI0/XI0_57/d_1_ DECAP_INV_G11
XG12883 XI11_1/XI0/XI0_57/d__0_ XI11_1/XI0/XI0_57/d_0_ DECAP_INV_G11
XG12884 XI11_1/XI0/XI0_57/d_15_ XI11_1/XI0/XI0_57/d__15_ DECAP_INV_G11
XG12885 XI11_1/XI0/XI0_57/d_14_ XI11_1/XI0/XI0_57/d__14_ DECAP_INV_G11
XG12886 XI11_1/XI0/XI0_57/d_13_ XI11_1/XI0/XI0_57/d__13_ DECAP_INV_G11
XG12887 XI11_1/XI0/XI0_57/d_12_ XI11_1/XI0/XI0_57/d__12_ DECAP_INV_G11
XG12888 XI11_1/XI0/XI0_57/d_11_ XI11_1/XI0/XI0_57/d__11_ DECAP_INV_G11
XG12889 XI11_1/XI0/XI0_57/d_10_ XI11_1/XI0/XI0_57/d__10_ DECAP_INV_G11
XG12890 XI11_1/XI0/XI0_57/d_9_ XI11_1/XI0/XI0_57/d__9_ DECAP_INV_G11
XG12891 XI11_1/XI0/XI0_57/d_8_ XI11_1/XI0/XI0_57/d__8_ DECAP_INV_G11
XG12892 XI11_1/XI0/XI0_57/d_7_ XI11_1/XI0/XI0_57/d__7_ DECAP_INV_G11
XG12893 XI11_1/XI0/XI0_57/d_6_ XI11_1/XI0/XI0_57/d__6_ DECAP_INV_G11
XG12894 XI11_1/XI0/XI0_57/d_5_ XI11_1/XI0/XI0_57/d__5_ DECAP_INV_G11
XG12895 XI11_1/XI0/XI0_57/d_4_ XI11_1/XI0/XI0_57/d__4_ DECAP_INV_G11
XG12896 XI11_1/XI0/XI0_57/d_3_ XI11_1/XI0/XI0_57/d__3_ DECAP_INV_G11
XG12897 XI11_1/XI0/XI0_57/d_2_ XI11_1/XI0/XI0_57/d__2_ DECAP_INV_G11
XG12898 XI11_1/XI0/XI0_57/d_1_ XI11_1/XI0/XI0_57/d__1_ DECAP_INV_G11
XG12899 XI11_1/XI0/XI0_57/d_0_ XI11_1/XI0/XI0_57/d__0_ DECAP_INV_G11
XG12900 XI11_1/XI0/XI0_56/d__15_ XI11_1/XI0/XI0_56/d_15_ DECAP_INV_G11
XG12901 XI11_1/XI0/XI0_56/d__14_ XI11_1/XI0/XI0_56/d_14_ DECAP_INV_G11
XG12902 XI11_1/XI0/XI0_56/d__13_ XI11_1/XI0/XI0_56/d_13_ DECAP_INV_G11
XG12903 XI11_1/XI0/XI0_56/d__12_ XI11_1/XI0/XI0_56/d_12_ DECAP_INV_G11
XG12904 XI11_1/XI0/XI0_56/d__11_ XI11_1/XI0/XI0_56/d_11_ DECAP_INV_G11
XG12905 XI11_1/XI0/XI0_56/d__10_ XI11_1/XI0/XI0_56/d_10_ DECAP_INV_G11
XG12906 XI11_1/XI0/XI0_56/d__9_ XI11_1/XI0/XI0_56/d_9_ DECAP_INV_G11
XG12907 XI11_1/XI0/XI0_56/d__8_ XI11_1/XI0/XI0_56/d_8_ DECAP_INV_G11
XG12908 XI11_1/XI0/XI0_56/d__7_ XI11_1/XI0/XI0_56/d_7_ DECAP_INV_G11
XG12909 XI11_1/XI0/XI0_56/d__6_ XI11_1/XI0/XI0_56/d_6_ DECAP_INV_G11
XG12910 XI11_1/XI0/XI0_56/d__5_ XI11_1/XI0/XI0_56/d_5_ DECAP_INV_G11
XG12911 XI11_1/XI0/XI0_56/d__4_ XI11_1/XI0/XI0_56/d_4_ DECAP_INV_G11
XG12912 XI11_1/XI0/XI0_56/d__3_ XI11_1/XI0/XI0_56/d_3_ DECAP_INV_G11
XG12913 XI11_1/XI0/XI0_56/d__2_ XI11_1/XI0/XI0_56/d_2_ DECAP_INV_G11
XG12914 XI11_1/XI0/XI0_56/d__1_ XI11_1/XI0/XI0_56/d_1_ DECAP_INV_G11
XG12915 XI11_1/XI0/XI0_56/d__0_ XI11_1/XI0/XI0_56/d_0_ DECAP_INV_G11
XG12916 XI11_1/XI0/XI0_56/d_15_ XI11_1/XI0/XI0_56/d__15_ DECAP_INV_G11
XG12917 XI11_1/XI0/XI0_56/d_14_ XI11_1/XI0/XI0_56/d__14_ DECAP_INV_G11
XG12918 XI11_1/XI0/XI0_56/d_13_ XI11_1/XI0/XI0_56/d__13_ DECAP_INV_G11
XG12919 XI11_1/XI0/XI0_56/d_12_ XI11_1/XI0/XI0_56/d__12_ DECAP_INV_G11
XG12920 XI11_1/XI0/XI0_56/d_11_ XI11_1/XI0/XI0_56/d__11_ DECAP_INV_G11
XG12921 XI11_1/XI0/XI0_56/d_10_ XI11_1/XI0/XI0_56/d__10_ DECAP_INV_G11
XG12922 XI11_1/XI0/XI0_56/d_9_ XI11_1/XI0/XI0_56/d__9_ DECAP_INV_G11
XG12923 XI11_1/XI0/XI0_56/d_8_ XI11_1/XI0/XI0_56/d__8_ DECAP_INV_G11
XG12924 XI11_1/XI0/XI0_56/d_7_ XI11_1/XI0/XI0_56/d__7_ DECAP_INV_G11
XG12925 XI11_1/XI0/XI0_56/d_6_ XI11_1/XI0/XI0_56/d__6_ DECAP_INV_G11
XG12926 XI11_1/XI0/XI0_56/d_5_ XI11_1/XI0/XI0_56/d__5_ DECAP_INV_G11
XG12927 XI11_1/XI0/XI0_56/d_4_ XI11_1/XI0/XI0_56/d__4_ DECAP_INV_G11
XG12928 XI11_1/XI0/XI0_56/d_3_ XI11_1/XI0/XI0_56/d__3_ DECAP_INV_G11
XG12929 XI11_1/XI0/XI0_56/d_2_ XI11_1/XI0/XI0_56/d__2_ DECAP_INV_G11
XG12930 XI11_1/XI0/XI0_56/d_1_ XI11_1/XI0/XI0_56/d__1_ DECAP_INV_G11
XG12931 XI11_1/XI0/XI0_56/d_0_ XI11_1/XI0/XI0_56/d__0_ DECAP_INV_G11
XG12932 XI11_1/XI0/XI0_55/d__15_ XI11_1/XI0/XI0_55/d_15_ DECAP_INV_G11
XG12933 XI11_1/XI0/XI0_55/d__14_ XI11_1/XI0/XI0_55/d_14_ DECAP_INV_G11
XG12934 XI11_1/XI0/XI0_55/d__13_ XI11_1/XI0/XI0_55/d_13_ DECAP_INV_G11
XG12935 XI11_1/XI0/XI0_55/d__12_ XI11_1/XI0/XI0_55/d_12_ DECAP_INV_G11
XG12936 XI11_1/XI0/XI0_55/d__11_ XI11_1/XI0/XI0_55/d_11_ DECAP_INV_G11
XG12937 XI11_1/XI0/XI0_55/d__10_ XI11_1/XI0/XI0_55/d_10_ DECAP_INV_G11
XG12938 XI11_1/XI0/XI0_55/d__9_ XI11_1/XI0/XI0_55/d_9_ DECAP_INV_G11
XG12939 XI11_1/XI0/XI0_55/d__8_ XI11_1/XI0/XI0_55/d_8_ DECAP_INV_G11
XG12940 XI11_1/XI0/XI0_55/d__7_ XI11_1/XI0/XI0_55/d_7_ DECAP_INV_G11
XG12941 XI11_1/XI0/XI0_55/d__6_ XI11_1/XI0/XI0_55/d_6_ DECAP_INV_G11
XG12942 XI11_1/XI0/XI0_55/d__5_ XI11_1/XI0/XI0_55/d_5_ DECAP_INV_G11
XG12943 XI11_1/XI0/XI0_55/d__4_ XI11_1/XI0/XI0_55/d_4_ DECAP_INV_G11
XG12944 XI11_1/XI0/XI0_55/d__3_ XI11_1/XI0/XI0_55/d_3_ DECAP_INV_G11
XG12945 XI11_1/XI0/XI0_55/d__2_ XI11_1/XI0/XI0_55/d_2_ DECAP_INV_G11
XG12946 XI11_1/XI0/XI0_55/d__1_ XI11_1/XI0/XI0_55/d_1_ DECAP_INV_G11
XG12947 XI11_1/XI0/XI0_55/d__0_ XI11_1/XI0/XI0_55/d_0_ DECAP_INV_G11
XG12948 XI11_1/XI0/XI0_55/d_15_ XI11_1/XI0/XI0_55/d__15_ DECAP_INV_G11
XG12949 XI11_1/XI0/XI0_55/d_14_ XI11_1/XI0/XI0_55/d__14_ DECAP_INV_G11
XG12950 XI11_1/XI0/XI0_55/d_13_ XI11_1/XI0/XI0_55/d__13_ DECAP_INV_G11
XG12951 XI11_1/XI0/XI0_55/d_12_ XI11_1/XI0/XI0_55/d__12_ DECAP_INV_G11
XG12952 XI11_1/XI0/XI0_55/d_11_ XI11_1/XI0/XI0_55/d__11_ DECAP_INV_G11
XG12953 XI11_1/XI0/XI0_55/d_10_ XI11_1/XI0/XI0_55/d__10_ DECAP_INV_G11
XG12954 XI11_1/XI0/XI0_55/d_9_ XI11_1/XI0/XI0_55/d__9_ DECAP_INV_G11
XG12955 XI11_1/XI0/XI0_55/d_8_ XI11_1/XI0/XI0_55/d__8_ DECAP_INV_G11
XG12956 XI11_1/XI0/XI0_55/d_7_ XI11_1/XI0/XI0_55/d__7_ DECAP_INV_G11
XG12957 XI11_1/XI0/XI0_55/d_6_ XI11_1/XI0/XI0_55/d__6_ DECAP_INV_G11
XG12958 XI11_1/XI0/XI0_55/d_5_ XI11_1/XI0/XI0_55/d__5_ DECAP_INV_G11
XG12959 XI11_1/XI0/XI0_55/d_4_ XI11_1/XI0/XI0_55/d__4_ DECAP_INV_G11
XG12960 XI11_1/XI0/XI0_55/d_3_ XI11_1/XI0/XI0_55/d__3_ DECAP_INV_G11
XG12961 XI11_1/XI0/XI0_55/d_2_ XI11_1/XI0/XI0_55/d__2_ DECAP_INV_G11
XG12962 XI11_1/XI0/XI0_55/d_1_ XI11_1/XI0/XI0_55/d__1_ DECAP_INV_G11
XG12963 XI11_1/XI0/XI0_55/d_0_ XI11_1/XI0/XI0_55/d__0_ DECAP_INV_G11
XG12964 XI11_1/XI0/XI0_54/d__15_ XI11_1/XI0/XI0_54/d_15_ DECAP_INV_G11
XG12965 XI11_1/XI0/XI0_54/d__14_ XI11_1/XI0/XI0_54/d_14_ DECAP_INV_G11
XG12966 XI11_1/XI0/XI0_54/d__13_ XI11_1/XI0/XI0_54/d_13_ DECAP_INV_G11
XG12967 XI11_1/XI0/XI0_54/d__12_ XI11_1/XI0/XI0_54/d_12_ DECAP_INV_G11
XG12968 XI11_1/XI0/XI0_54/d__11_ XI11_1/XI0/XI0_54/d_11_ DECAP_INV_G11
XG12969 XI11_1/XI0/XI0_54/d__10_ XI11_1/XI0/XI0_54/d_10_ DECAP_INV_G11
XG12970 XI11_1/XI0/XI0_54/d__9_ XI11_1/XI0/XI0_54/d_9_ DECAP_INV_G11
XG12971 XI11_1/XI0/XI0_54/d__8_ XI11_1/XI0/XI0_54/d_8_ DECAP_INV_G11
XG12972 XI11_1/XI0/XI0_54/d__7_ XI11_1/XI0/XI0_54/d_7_ DECAP_INV_G11
XG12973 XI11_1/XI0/XI0_54/d__6_ XI11_1/XI0/XI0_54/d_6_ DECAP_INV_G11
XG12974 XI11_1/XI0/XI0_54/d__5_ XI11_1/XI0/XI0_54/d_5_ DECAP_INV_G11
XG12975 XI11_1/XI0/XI0_54/d__4_ XI11_1/XI0/XI0_54/d_4_ DECAP_INV_G11
XG12976 XI11_1/XI0/XI0_54/d__3_ XI11_1/XI0/XI0_54/d_3_ DECAP_INV_G11
XG12977 XI11_1/XI0/XI0_54/d__2_ XI11_1/XI0/XI0_54/d_2_ DECAP_INV_G11
XG12978 XI11_1/XI0/XI0_54/d__1_ XI11_1/XI0/XI0_54/d_1_ DECAP_INV_G11
XG12979 XI11_1/XI0/XI0_54/d__0_ XI11_1/XI0/XI0_54/d_0_ DECAP_INV_G11
XG12980 XI11_1/XI0/XI0_54/d_15_ XI11_1/XI0/XI0_54/d__15_ DECAP_INV_G11
XG12981 XI11_1/XI0/XI0_54/d_14_ XI11_1/XI0/XI0_54/d__14_ DECAP_INV_G11
XG12982 XI11_1/XI0/XI0_54/d_13_ XI11_1/XI0/XI0_54/d__13_ DECAP_INV_G11
XG12983 XI11_1/XI0/XI0_54/d_12_ XI11_1/XI0/XI0_54/d__12_ DECAP_INV_G11
XG12984 XI11_1/XI0/XI0_54/d_11_ XI11_1/XI0/XI0_54/d__11_ DECAP_INV_G11
XG12985 XI11_1/XI0/XI0_54/d_10_ XI11_1/XI0/XI0_54/d__10_ DECAP_INV_G11
XG12986 XI11_1/XI0/XI0_54/d_9_ XI11_1/XI0/XI0_54/d__9_ DECAP_INV_G11
XG12987 XI11_1/XI0/XI0_54/d_8_ XI11_1/XI0/XI0_54/d__8_ DECAP_INV_G11
XG12988 XI11_1/XI0/XI0_54/d_7_ XI11_1/XI0/XI0_54/d__7_ DECAP_INV_G11
XG12989 XI11_1/XI0/XI0_54/d_6_ XI11_1/XI0/XI0_54/d__6_ DECAP_INV_G11
XG12990 XI11_1/XI0/XI0_54/d_5_ XI11_1/XI0/XI0_54/d__5_ DECAP_INV_G11
XG12991 XI11_1/XI0/XI0_54/d_4_ XI11_1/XI0/XI0_54/d__4_ DECAP_INV_G11
XG12992 XI11_1/XI0/XI0_54/d_3_ XI11_1/XI0/XI0_54/d__3_ DECAP_INV_G11
XG12993 XI11_1/XI0/XI0_54/d_2_ XI11_1/XI0/XI0_54/d__2_ DECAP_INV_G11
XG12994 XI11_1/XI0/XI0_54/d_1_ XI11_1/XI0/XI0_54/d__1_ DECAP_INV_G11
XG12995 XI11_1/XI0/XI0_54/d_0_ XI11_1/XI0/XI0_54/d__0_ DECAP_INV_G11
XG12996 XI11_1/XI0/XI0_53/d__15_ XI11_1/XI0/XI0_53/d_15_ DECAP_INV_G11
XG12997 XI11_1/XI0/XI0_53/d__14_ XI11_1/XI0/XI0_53/d_14_ DECAP_INV_G11
XG12998 XI11_1/XI0/XI0_53/d__13_ XI11_1/XI0/XI0_53/d_13_ DECAP_INV_G11
XG12999 XI11_1/XI0/XI0_53/d__12_ XI11_1/XI0/XI0_53/d_12_ DECAP_INV_G11
XG13000 XI11_1/XI0/XI0_53/d__11_ XI11_1/XI0/XI0_53/d_11_ DECAP_INV_G11
XG13001 XI11_1/XI0/XI0_53/d__10_ XI11_1/XI0/XI0_53/d_10_ DECAP_INV_G11
XG13002 XI11_1/XI0/XI0_53/d__9_ XI11_1/XI0/XI0_53/d_9_ DECAP_INV_G11
XG13003 XI11_1/XI0/XI0_53/d__8_ XI11_1/XI0/XI0_53/d_8_ DECAP_INV_G11
XG13004 XI11_1/XI0/XI0_53/d__7_ XI11_1/XI0/XI0_53/d_7_ DECAP_INV_G11
XG13005 XI11_1/XI0/XI0_53/d__6_ XI11_1/XI0/XI0_53/d_6_ DECAP_INV_G11
XG13006 XI11_1/XI0/XI0_53/d__5_ XI11_1/XI0/XI0_53/d_5_ DECAP_INV_G11
XG13007 XI11_1/XI0/XI0_53/d__4_ XI11_1/XI0/XI0_53/d_4_ DECAP_INV_G11
XG13008 XI11_1/XI0/XI0_53/d__3_ XI11_1/XI0/XI0_53/d_3_ DECAP_INV_G11
XG13009 XI11_1/XI0/XI0_53/d__2_ XI11_1/XI0/XI0_53/d_2_ DECAP_INV_G11
XG13010 XI11_1/XI0/XI0_53/d__1_ XI11_1/XI0/XI0_53/d_1_ DECAP_INV_G11
XG13011 XI11_1/XI0/XI0_53/d__0_ XI11_1/XI0/XI0_53/d_0_ DECAP_INV_G11
XG13012 XI11_1/XI0/XI0_53/d_15_ XI11_1/XI0/XI0_53/d__15_ DECAP_INV_G11
XG13013 XI11_1/XI0/XI0_53/d_14_ XI11_1/XI0/XI0_53/d__14_ DECAP_INV_G11
XG13014 XI11_1/XI0/XI0_53/d_13_ XI11_1/XI0/XI0_53/d__13_ DECAP_INV_G11
XG13015 XI11_1/XI0/XI0_53/d_12_ XI11_1/XI0/XI0_53/d__12_ DECAP_INV_G11
XG13016 XI11_1/XI0/XI0_53/d_11_ XI11_1/XI0/XI0_53/d__11_ DECAP_INV_G11
XG13017 XI11_1/XI0/XI0_53/d_10_ XI11_1/XI0/XI0_53/d__10_ DECAP_INV_G11
XG13018 XI11_1/XI0/XI0_53/d_9_ XI11_1/XI0/XI0_53/d__9_ DECAP_INV_G11
XG13019 XI11_1/XI0/XI0_53/d_8_ XI11_1/XI0/XI0_53/d__8_ DECAP_INV_G11
XG13020 XI11_1/XI0/XI0_53/d_7_ XI11_1/XI0/XI0_53/d__7_ DECAP_INV_G11
XG13021 XI11_1/XI0/XI0_53/d_6_ XI11_1/XI0/XI0_53/d__6_ DECAP_INV_G11
XG13022 XI11_1/XI0/XI0_53/d_5_ XI11_1/XI0/XI0_53/d__5_ DECAP_INV_G11
XG13023 XI11_1/XI0/XI0_53/d_4_ XI11_1/XI0/XI0_53/d__4_ DECAP_INV_G11
XG13024 XI11_1/XI0/XI0_53/d_3_ XI11_1/XI0/XI0_53/d__3_ DECAP_INV_G11
XG13025 XI11_1/XI0/XI0_53/d_2_ XI11_1/XI0/XI0_53/d__2_ DECAP_INV_G11
XG13026 XI11_1/XI0/XI0_53/d_1_ XI11_1/XI0/XI0_53/d__1_ DECAP_INV_G11
XG13027 XI11_1/XI0/XI0_53/d_0_ XI11_1/XI0/XI0_53/d__0_ DECAP_INV_G11
XG13028 XI11_1/XI0/XI0_52/d__15_ XI11_1/XI0/XI0_52/d_15_ DECAP_INV_G11
XG13029 XI11_1/XI0/XI0_52/d__14_ XI11_1/XI0/XI0_52/d_14_ DECAP_INV_G11
XG13030 XI11_1/XI0/XI0_52/d__13_ XI11_1/XI0/XI0_52/d_13_ DECAP_INV_G11
XG13031 XI11_1/XI0/XI0_52/d__12_ XI11_1/XI0/XI0_52/d_12_ DECAP_INV_G11
XG13032 XI11_1/XI0/XI0_52/d__11_ XI11_1/XI0/XI0_52/d_11_ DECAP_INV_G11
XG13033 XI11_1/XI0/XI0_52/d__10_ XI11_1/XI0/XI0_52/d_10_ DECAP_INV_G11
XG13034 XI11_1/XI0/XI0_52/d__9_ XI11_1/XI0/XI0_52/d_9_ DECAP_INV_G11
XG13035 XI11_1/XI0/XI0_52/d__8_ XI11_1/XI0/XI0_52/d_8_ DECAP_INV_G11
XG13036 XI11_1/XI0/XI0_52/d__7_ XI11_1/XI0/XI0_52/d_7_ DECAP_INV_G11
XG13037 XI11_1/XI0/XI0_52/d__6_ XI11_1/XI0/XI0_52/d_6_ DECAP_INV_G11
XG13038 XI11_1/XI0/XI0_52/d__5_ XI11_1/XI0/XI0_52/d_5_ DECAP_INV_G11
XG13039 XI11_1/XI0/XI0_52/d__4_ XI11_1/XI0/XI0_52/d_4_ DECAP_INV_G11
XG13040 XI11_1/XI0/XI0_52/d__3_ XI11_1/XI0/XI0_52/d_3_ DECAP_INV_G11
XG13041 XI11_1/XI0/XI0_52/d__2_ XI11_1/XI0/XI0_52/d_2_ DECAP_INV_G11
XG13042 XI11_1/XI0/XI0_52/d__1_ XI11_1/XI0/XI0_52/d_1_ DECAP_INV_G11
XG13043 XI11_1/XI0/XI0_52/d__0_ XI11_1/XI0/XI0_52/d_0_ DECAP_INV_G11
XG13044 XI11_1/XI0/XI0_52/d_15_ XI11_1/XI0/XI0_52/d__15_ DECAP_INV_G11
XG13045 XI11_1/XI0/XI0_52/d_14_ XI11_1/XI0/XI0_52/d__14_ DECAP_INV_G11
XG13046 XI11_1/XI0/XI0_52/d_13_ XI11_1/XI0/XI0_52/d__13_ DECAP_INV_G11
XG13047 XI11_1/XI0/XI0_52/d_12_ XI11_1/XI0/XI0_52/d__12_ DECAP_INV_G11
XG13048 XI11_1/XI0/XI0_52/d_11_ XI11_1/XI0/XI0_52/d__11_ DECAP_INV_G11
XG13049 XI11_1/XI0/XI0_52/d_10_ XI11_1/XI0/XI0_52/d__10_ DECAP_INV_G11
XG13050 XI11_1/XI0/XI0_52/d_9_ XI11_1/XI0/XI0_52/d__9_ DECAP_INV_G11
XG13051 XI11_1/XI0/XI0_52/d_8_ XI11_1/XI0/XI0_52/d__8_ DECAP_INV_G11
XG13052 XI11_1/XI0/XI0_52/d_7_ XI11_1/XI0/XI0_52/d__7_ DECAP_INV_G11
XG13053 XI11_1/XI0/XI0_52/d_6_ XI11_1/XI0/XI0_52/d__6_ DECAP_INV_G11
XG13054 XI11_1/XI0/XI0_52/d_5_ XI11_1/XI0/XI0_52/d__5_ DECAP_INV_G11
XG13055 XI11_1/XI0/XI0_52/d_4_ XI11_1/XI0/XI0_52/d__4_ DECAP_INV_G11
XG13056 XI11_1/XI0/XI0_52/d_3_ XI11_1/XI0/XI0_52/d__3_ DECAP_INV_G11
XG13057 XI11_1/XI0/XI0_52/d_2_ XI11_1/XI0/XI0_52/d__2_ DECAP_INV_G11
XG13058 XI11_1/XI0/XI0_52/d_1_ XI11_1/XI0/XI0_52/d__1_ DECAP_INV_G11
XG13059 XI11_1/XI0/XI0_52/d_0_ XI11_1/XI0/XI0_52/d__0_ DECAP_INV_G11
XG13060 XI11_1/XI0/XI0_51/d__15_ XI11_1/XI0/XI0_51/d_15_ DECAP_INV_G11
XG13061 XI11_1/XI0/XI0_51/d__14_ XI11_1/XI0/XI0_51/d_14_ DECAP_INV_G11
XG13062 XI11_1/XI0/XI0_51/d__13_ XI11_1/XI0/XI0_51/d_13_ DECAP_INV_G11
XG13063 XI11_1/XI0/XI0_51/d__12_ XI11_1/XI0/XI0_51/d_12_ DECAP_INV_G11
XG13064 XI11_1/XI0/XI0_51/d__11_ XI11_1/XI0/XI0_51/d_11_ DECAP_INV_G11
XG13065 XI11_1/XI0/XI0_51/d__10_ XI11_1/XI0/XI0_51/d_10_ DECAP_INV_G11
XG13066 XI11_1/XI0/XI0_51/d__9_ XI11_1/XI0/XI0_51/d_9_ DECAP_INV_G11
XG13067 XI11_1/XI0/XI0_51/d__8_ XI11_1/XI0/XI0_51/d_8_ DECAP_INV_G11
XG13068 XI11_1/XI0/XI0_51/d__7_ XI11_1/XI0/XI0_51/d_7_ DECAP_INV_G11
XG13069 XI11_1/XI0/XI0_51/d__6_ XI11_1/XI0/XI0_51/d_6_ DECAP_INV_G11
XG13070 XI11_1/XI0/XI0_51/d__5_ XI11_1/XI0/XI0_51/d_5_ DECAP_INV_G11
XG13071 XI11_1/XI0/XI0_51/d__4_ XI11_1/XI0/XI0_51/d_4_ DECAP_INV_G11
XG13072 XI11_1/XI0/XI0_51/d__3_ XI11_1/XI0/XI0_51/d_3_ DECAP_INV_G11
XG13073 XI11_1/XI0/XI0_51/d__2_ XI11_1/XI0/XI0_51/d_2_ DECAP_INV_G11
XG13074 XI11_1/XI0/XI0_51/d__1_ XI11_1/XI0/XI0_51/d_1_ DECAP_INV_G11
XG13075 XI11_1/XI0/XI0_51/d__0_ XI11_1/XI0/XI0_51/d_0_ DECAP_INV_G11
XG13076 XI11_1/XI0/XI0_51/d_15_ XI11_1/XI0/XI0_51/d__15_ DECAP_INV_G11
XG13077 XI11_1/XI0/XI0_51/d_14_ XI11_1/XI0/XI0_51/d__14_ DECAP_INV_G11
XG13078 XI11_1/XI0/XI0_51/d_13_ XI11_1/XI0/XI0_51/d__13_ DECAP_INV_G11
XG13079 XI11_1/XI0/XI0_51/d_12_ XI11_1/XI0/XI0_51/d__12_ DECAP_INV_G11
XG13080 XI11_1/XI0/XI0_51/d_11_ XI11_1/XI0/XI0_51/d__11_ DECAP_INV_G11
XG13081 XI11_1/XI0/XI0_51/d_10_ XI11_1/XI0/XI0_51/d__10_ DECAP_INV_G11
XG13082 XI11_1/XI0/XI0_51/d_9_ XI11_1/XI0/XI0_51/d__9_ DECAP_INV_G11
XG13083 XI11_1/XI0/XI0_51/d_8_ XI11_1/XI0/XI0_51/d__8_ DECAP_INV_G11
XG13084 XI11_1/XI0/XI0_51/d_7_ XI11_1/XI0/XI0_51/d__7_ DECAP_INV_G11
XG13085 XI11_1/XI0/XI0_51/d_6_ XI11_1/XI0/XI0_51/d__6_ DECAP_INV_G11
XG13086 XI11_1/XI0/XI0_51/d_5_ XI11_1/XI0/XI0_51/d__5_ DECAP_INV_G11
XG13087 XI11_1/XI0/XI0_51/d_4_ XI11_1/XI0/XI0_51/d__4_ DECAP_INV_G11
XG13088 XI11_1/XI0/XI0_51/d_3_ XI11_1/XI0/XI0_51/d__3_ DECAP_INV_G11
XG13089 XI11_1/XI0/XI0_51/d_2_ XI11_1/XI0/XI0_51/d__2_ DECAP_INV_G11
XG13090 XI11_1/XI0/XI0_51/d_1_ XI11_1/XI0/XI0_51/d__1_ DECAP_INV_G11
XG13091 XI11_1/XI0/XI0_51/d_0_ XI11_1/XI0/XI0_51/d__0_ DECAP_INV_G11
XG13092 XI11_1/XI0/XI0_50/d__15_ XI11_1/XI0/XI0_50/d_15_ DECAP_INV_G11
XG13093 XI11_1/XI0/XI0_50/d__14_ XI11_1/XI0/XI0_50/d_14_ DECAP_INV_G11
XG13094 XI11_1/XI0/XI0_50/d__13_ XI11_1/XI0/XI0_50/d_13_ DECAP_INV_G11
XG13095 XI11_1/XI0/XI0_50/d__12_ XI11_1/XI0/XI0_50/d_12_ DECAP_INV_G11
XG13096 XI11_1/XI0/XI0_50/d__11_ XI11_1/XI0/XI0_50/d_11_ DECAP_INV_G11
XG13097 XI11_1/XI0/XI0_50/d__10_ XI11_1/XI0/XI0_50/d_10_ DECAP_INV_G11
XG13098 XI11_1/XI0/XI0_50/d__9_ XI11_1/XI0/XI0_50/d_9_ DECAP_INV_G11
XG13099 XI11_1/XI0/XI0_50/d__8_ XI11_1/XI0/XI0_50/d_8_ DECAP_INV_G11
XG13100 XI11_1/XI0/XI0_50/d__7_ XI11_1/XI0/XI0_50/d_7_ DECAP_INV_G11
XG13101 XI11_1/XI0/XI0_50/d__6_ XI11_1/XI0/XI0_50/d_6_ DECAP_INV_G11
XG13102 XI11_1/XI0/XI0_50/d__5_ XI11_1/XI0/XI0_50/d_5_ DECAP_INV_G11
XG13103 XI11_1/XI0/XI0_50/d__4_ XI11_1/XI0/XI0_50/d_4_ DECAP_INV_G11
XG13104 XI11_1/XI0/XI0_50/d__3_ XI11_1/XI0/XI0_50/d_3_ DECAP_INV_G11
XG13105 XI11_1/XI0/XI0_50/d__2_ XI11_1/XI0/XI0_50/d_2_ DECAP_INV_G11
XG13106 XI11_1/XI0/XI0_50/d__1_ XI11_1/XI0/XI0_50/d_1_ DECAP_INV_G11
XG13107 XI11_1/XI0/XI0_50/d__0_ XI11_1/XI0/XI0_50/d_0_ DECAP_INV_G11
XG13108 XI11_1/XI0/XI0_50/d_15_ XI11_1/XI0/XI0_50/d__15_ DECAP_INV_G11
XG13109 XI11_1/XI0/XI0_50/d_14_ XI11_1/XI0/XI0_50/d__14_ DECAP_INV_G11
XG13110 XI11_1/XI0/XI0_50/d_13_ XI11_1/XI0/XI0_50/d__13_ DECAP_INV_G11
XG13111 XI11_1/XI0/XI0_50/d_12_ XI11_1/XI0/XI0_50/d__12_ DECAP_INV_G11
XG13112 XI11_1/XI0/XI0_50/d_11_ XI11_1/XI0/XI0_50/d__11_ DECAP_INV_G11
XG13113 XI11_1/XI0/XI0_50/d_10_ XI11_1/XI0/XI0_50/d__10_ DECAP_INV_G11
XG13114 XI11_1/XI0/XI0_50/d_9_ XI11_1/XI0/XI0_50/d__9_ DECAP_INV_G11
XG13115 XI11_1/XI0/XI0_50/d_8_ XI11_1/XI0/XI0_50/d__8_ DECAP_INV_G11
XG13116 XI11_1/XI0/XI0_50/d_7_ XI11_1/XI0/XI0_50/d__7_ DECAP_INV_G11
XG13117 XI11_1/XI0/XI0_50/d_6_ XI11_1/XI0/XI0_50/d__6_ DECAP_INV_G11
XG13118 XI11_1/XI0/XI0_50/d_5_ XI11_1/XI0/XI0_50/d__5_ DECAP_INV_G11
XG13119 XI11_1/XI0/XI0_50/d_4_ XI11_1/XI0/XI0_50/d__4_ DECAP_INV_G11
XG13120 XI11_1/XI0/XI0_50/d_3_ XI11_1/XI0/XI0_50/d__3_ DECAP_INV_G11
XG13121 XI11_1/XI0/XI0_50/d_2_ XI11_1/XI0/XI0_50/d__2_ DECAP_INV_G11
XG13122 XI11_1/XI0/XI0_50/d_1_ XI11_1/XI0/XI0_50/d__1_ DECAP_INV_G11
XG13123 XI11_1/XI0/XI0_50/d_0_ XI11_1/XI0/XI0_50/d__0_ DECAP_INV_G11
XG13124 XI11_1/XI0/XI0_49/d__15_ XI11_1/XI0/XI0_49/d_15_ DECAP_INV_G11
XG13125 XI11_1/XI0/XI0_49/d__14_ XI11_1/XI0/XI0_49/d_14_ DECAP_INV_G11
XG13126 XI11_1/XI0/XI0_49/d__13_ XI11_1/XI0/XI0_49/d_13_ DECAP_INV_G11
XG13127 XI11_1/XI0/XI0_49/d__12_ XI11_1/XI0/XI0_49/d_12_ DECAP_INV_G11
XG13128 XI11_1/XI0/XI0_49/d__11_ XI11_1/XI0/XI0_49/d_11_ DECAP_INV_G11
XG13129 XI11_1/XI0/XI0_49/d__10_ XI11_1/XI0/XI0_49/d_10_ DECAP_INV_G11
XG13130 XI11_1/XI0/XI0_49/d__9_ XI11_1/XI0/XI0_49/d_9_ DECAP_INV_G11
XG13131 XI11_1/XI0/XI0_49/d__8_ XI11_1/XI0/XI0_49/d_8_ DECAP_INV_G11
XG13132 XI11_1/XI0/XI0_49/d__7_ XI11_1/XI0/XI0_49/d_7_ DECAP_INV_G11
XG13133 XI11_1/XI0/XI0_49/d__6_ XI11_1/XI0/XI0_49/d_6_ DECAP_INV_G11
XG13134 XI11_1/XI0/XI0_49/d__5_ XI11_1/XI0/XI0_49/d_5_ DECAP_INV_G11
XG13135 XI11_1/XI0/XI0_49/d__4_ XI11_1/XI0/XI0_49/d_4_ DECAP_INV_G11
XG13136 XI11_1/XI0/XI0_49/d__3_ XI11_1/XI0/XI0_49/d_3_ DECAP_INV_G11
XG13137 XI11_1/XI0/XI0_49/d__2_ XI11_1/XI0/XI0_49/d_2_ DECAP_INV_G11
XG13138 XI11_1/XI0/XI0_49/d__1_ XI11_1/XI0/XI0_49/d_1_ DECAP_INV_G11
XG13139 XI11_1/XI0/XI0_49/d__0_ XI11_1/XI0/XI0_49/d_0_ DECAP_INV_G11
XG13140 XI11_1/XI0/XI0_49/d_15_ XI11_1/XI0/XI0_49/d__15_ DECAP_INV_G11
XG13141 XI11_1/XI0/XI0_49/d_14_ XI11_1/XI0/XI0_49/d__14_ DECAP_INV_G11
XG13142 XI11_1/XI0/XI0_49/d_13_ XI11_1/XI0/XI0_49/d__13_ DECAP_INV_G11
XG13143 XI11_1/XI0/XI0_49/d_12_ XI11_1/XI0/XI0_49/d__12_ DECAP_INV_G11
XG13144 XI11_1/XI0/XI0_49/d_11_ XI11_1/XI0/XI0_49/d__11_ DECAP_INV_G11
XG13145 XI11_1/XI0/XI0_49/d_10_ XI11_1/XI0/XI0_49/d__10_ DECAP_INV_G11
XG13146 XI11_1/XI0/XI0_49/d_9_ XI11_1/XI0/XI0_49/d__9_ DECAP_INV_G11
XG13147 XI11_1/XI0/XI0_49/d_8_ XI11_1/XI0/XI0_49/d__8_ DECAP_INV_G11
XG13148 XI11_1/XI0/XI0_49/d_7_ XI11_1/XI0/XI0_49/d__7_ DECAP_INV_G11
XG13149 XI11_1/XI0/XI0_49/d_6_ XI11_1/XI0/XI0_49/d__6_ DECAP_INV_G11
XG13150 XI11_1/XI0/XI0_49/d_5_ XI11_1/XI0/XI0_49/d__5_ DECAP_INV_G11
XG13151 XI11_1/XI0/XI0_49/d_4_ XI11_1/XI0/XI0_49/d__4_ DECAP_INV_G11
XG13152 XI11_1/XI0/XI0_49/d_3_ XI11_1/XI0/XI0_49/d__3_ DECAP_INV_G11
XG13153 XI11_1/XI0/XI0_49/d_2_ XI11_1/XI0/XI0_49/d__2_ DECAP_INV_G11
XG13154 XI11_1/XI0/XI0_49/d_1_ XI11_1/XI0/XI0_49/d__1_ DECAP_INV_G11
XG13155 XI11_1/XI0/XI0_49/d_0_ XI11_1/XI0/XI0_49/d__0_ DECAP_INV_G11
XG13156 XI11_1/XI0/XI0_48/d__15_ XI11_1/XI0/XI0_48/d_15_ DECAP_INV_G11
XG13157 XI11_1/XI0/XI0_48/d__14_ XI11_1/XI0/XI0_48/d_14_ DECAP_INV_G11
XG13158 XI11_1/XI0/XI0_48/d__13_ XI11_1/XI0/XI0_48/d_13_ DECAP_INV_G11
XG13159 XI11_1/XI0/XI0_48/d__12_ XI11_1/XI0/XI0_48/d_12_ DECAP_INV_G11
XG13160 XI11_1/XI0/XI0_48/d__11_ XI11_1/XI0/XI0_48/d_11_ DECAP_INV_G11
XG13161 XI11_1/XI0/XI0_48/d__10_ XI11_1/XI0/XI0_48/d_10_ DECAP_INV_G11
XG13162 XI11_1/XI0/XI0_48/d__9_ XI11_1/XI0/XI0_48/d_9_ DECAP_INV_G11
XG13163 XI11_1/XI0/XI0_48/d__8_ XI11_1/XI0/XI0_48/d_8_ DECAP_INV_G11
XG13164 XI11_1/XI0/XI0_48/d__7_ XI11_1/XI0/XI0_48/d_7_ DECAP_INV_G11
XG13165 XI11_1/XI0/XI0_48/d__6_ XI11_1/XI0/XI0_48/d_6_ DECAP_INV_G11
XG13166 XI11_1/XI0/XI0_48/d__5_ XI11_1/XI0/XI0_48/d_5_ DECAP_INV_G11
XG13167 XI11_1/XI0/XI0_48/d__4_ XI11_1/XI0/XI0_48/d_4_ DECAP_INV_G11
XG13168 XI11_1/XI0/XI0_48/d__3_ XI11_1/XI0/XI0_48/d_3_ DECAP_INV_G11
XG13169 XI11_1/XI0/XI0_48/d__2_ XI11_1/XI0/XI0_48/d_2_ DECAP_INV_G11
XG13170 XI11_1/XI0/XI0_48/d__1_ XI11_1/XI0/XI0_48/d_1_ DECAP_INV_G11
XG13171 XI11_1/XI0/XI0_48/d__0_ XI11_1/XI0/XI0_48/d_0_ DECAP_INV_G11
XG13172 XI11_1/XI0/XI0_48/d_15_ XI11_1/XI0/XI0_48/d__15_ DECAP_INV_G11
XG13173 XI11_1/XI0/XI0_48/d_14_ XI11_1/XI0/XI0_48/d__14_ DECAP_INV_G11
XG13174 XI11_1/XI0/XI0_48/d_13_ XI11_1/XI0/XI0_48/d__13_ DECAP_INV_G11
XG13175 XI11_1/XI0/XI0_48/d_12_ XI11_1/XI0/XI0_48/d__12_ DECAP_INV_G11
XG13176 XI11_1/XI0/XI0_48/d_11_ XI11_1/XI0/XI0_48/d__11_ DECAP_INV_G11
XG13177 XI11_1/XI0/XI0_48/d_10_ XI11_1/XI0/XI0_48/d__10_ DECAP_INV_G11
XG13178 XI11_1/XI0/XI0_48/d_9_ XI11_1/XI0/XI0_48/d__9_ DECAP_INV_G11
XG13179 XI11_1/XI0/XI0_48/d_8_ XI11_1/XI0/XI0_48/d__8_ DECAP_INV_G11
XG13180 XI11_1/XI0/XI0_48/d_7_ XI11_1/XI0/XI0_48/d__7_ DECAP_INV_G11
XG13181 XI11_1/XI0/XI0_48/d_6_ XI11_1/XI0/XI0_48/d__6_ DECAP_INV_G11
XG13182 XI11_1/XI0/XI0_48/d_5_ XI11_1/XI0/XI0_48/d__5_ DECAP_INV_G11
XG13183 XI11_1/XI0/XI0_48/d_4_ XI11_1/XI0/XI0_48/d__4_ DECAP_INV_G11
XG13184 XI11_1/XI0/XI0_48/d_3_ XI11_1/XI0/XI0_48/d__3_ DECAP_INV_G11
XG13185 XI11_1/XI0/XI0_48/d_2_ XI11_1/XI0/XI0_48/d__2_ DECAP_INV_G11
XG13186 XI11_1/XI0/XI0_48/d_1_ XI11_1/XI0/XI0_48/d__1_ DECAP_INV_G11
XG13187 XI11_1/XI0/XI0_48/d_0_ XI11_1/XI0/XI0_48/d__0_ DECAP_INV_G11
XG13188 XI11_1/XI0/XI0_47/d__15_ XI11_1/XI0/XI0_47/d_15_ DECAP_INV_G11
XG13189 XI11_1/XI0/XI0_47/d__14_ XI11_1/XI0/XI0_47/d_14_ DECAP_INV_G11
XG13190 XI11_1/XI0/XI0_47/d__13_ XI11_1/XI0/XI0_47/d_13_ DECAP_INV_G11
XG13191 XI11_1/XI0/XI0_47/d__12_ XI11_1/XI0/XI0_47/d_12_ DECAP_INV_G11
XG13192 XI11_1/XI0/XI0_47/d__11_ XI11_1/XI0/XI0_47/d_11_ DECAP_INV_G11
XG13193 XI11_1/XI0/XI0_47/d__10_ XI11_1/XI0/XI0_47/d_10_ DECAP_INV_G11
XG13194 XI11_1/XI0/XI0_47/d__9_ XI11_1/XI0/XI0_47/d_9_ DECAP_INV_G11
XG13195 XI11_1/XI0/XI0_47/d__8_ XI11_1/XI0/XI0_47/d_8_ DECAP_INV_G11
XG13196 XI11_1/XI0/XI0_47/d__7_ XI11_1/XI0/XI0_47/d_7_ DECAP_INV_G11
XG13197 XI11_1/XI0/XI0_47/d__6_ XI11_1/XI0/XI0_47/d_6_ DECAP_INV_G11
XG13198 XI11_1/XI0/XI0_47/d__5_ XI11_1/XI0/XI0_47/d_5_ DECAP_INV_G11
XG13199 XI11_1/XI0/XI0_47/d__4_ XI11_1/XI0/XI0_47/d_4_ DECAP_INV_G11
XG13200 XI11_1/XI0/XI0_47/d__3_ XI11_1/XI0/XI0_47/d_3_ DECAP_INV_G11
XG13201 XI11_1/XI0/XI0_47/d__2_ XI11_1/XI0/XI0_47/d_2_ DECAP_INV_G11
XG13202 XI11_1/XI0/XI0_47/d__1_ XI11_1/XI0/XI0_47/d_1_ DECAP_INV_G11
XG13203 XI11_1/XI0/XI0_47/d__0_ XI11_1/XI0/XI0_47/d_0_ DECAP_INV_G11
XG13204 XI11_1/XI0/XI0_47/d_15_ XI11_1/XI0/XI0_47/d__15_ DECAP_INV_G11
XG13205 XI11_1/XI0/XI0_47/d_14_ XI11_1/XI0/XI0_47/d__14_ DECAP_INV_G11
XG13206 XI11_1/XI0/XI0_47/d_13_ XI11_1/XI0/XI0_47/d__13_ DECAP_INV_G11
XG13207 XI11_1/XI0/XI0_47/d_12_ XI11_1/XI0/XI0_47/d__12_ DECAP_INV_G11
XG13208 XI11_1/XI0/XI0_47/d_11_ XI11_1/XI0/XI0_47/d__11_ DECAP_INV_G11
XG13209 XI11_1/XI0/XI0_47/d_10_ XI11_1/XI0/XI0_47/d__10_ DECAP_INV_G11
XG13210 XI11_1/XI0/XI0_47/d_9_ XI11_1/XI0/XI0_47/d__9_ DECAP_INV_G11
XG13211 XI11_1/XI0/XI0_47/d_8_ XI11_1/XI0/XI0_47/d__8_ DECAP_INV_G11
XG13212 XI11_1/XI0/XI0_47/d_7_ XI11_1/XI0/XI0_47/d__7_ DECAP_INV_G11
XG13213 XI11_1/XI0/XI0_47/d_6_ XI11_1/XI0/XI0_47/d__6_ DECAP_INV_G11
XG13214 XI11_1/XI0/XI0_47/d_5_ XI11_1/XI0/XI0_47/d__5_ DECAP_INV_G11
XG13215 XI11_1/XI0/XI0_47/d_4_ XI11_1/XI0/XI0_47/d__4_ DECAP_INV_G11
XG13216 XI11_1/XI0/XI0_47/d_3_ XI11_1/XI0/XI0_47/d__3_ DECAP_INV_G11
XG13217 XI11_1/XI0/XI0_47/d_2_ XI11_1/XI0/XI0_47/d__2_ DECAP_INV_G11
XG13218 XI11_1/XI0/XI0_47/d_1_ XI11_1/XI0/XI0_47/d__1_ DECAP_INV_G11
XG13219 XI11_1/XI0/XI0_47/d_0_ XI11_1/XI0/XI0_47/d__0_ DECAP_INV_G11
XG13220 XI11_1/XI0/XI0_46/d__15_ XI11_1/XI0/XI0_46/d_15_ DECAP_INV_G11
XG13221 XI11_1/XI0/XI0_46/d__14_ XI11_1/XI0/XI0_46/d_14_ DECAP_INV_G11
XG13222 XI11_1/XI0/XI0_46/d__13_ XI11_1/XI0/XI0_46/d_13_ DECAP_INV_G11
XG13223 XI11_1/XI0/XI0_46/d__12_ XI11_1/XI0/XI0_46/d_12_ DECAP_INV_G11
XG13224 XI11_1/XI0/XI0_46/d__11_ XI11_1/XI0/XI0_46/d_11_ DECAP_INV_G11
XG13225 XI11_1/XI0/XI0_46/d__10_ XI11_1/XI0/XI0_46/d_10_ DECAP_INV_G11
XG13226 XI11_1/XI0/XI0_46/d__9_ XI11_1/XI0/XI0_46/d_9_ DECAP_INV_G11
XG13227 XI11_1/XI0/XI0_46/d__8_ XI11_1/XI0/XI0_46/d_8_ DECAP_INV_G11
XG13228 XI11_1/XI0/XI0_46/d__7_ XI11_1/XI0/XI0_46/d_7_ DECAP_INV_G11
XG13229 XI11_1/XI0/XI0_46/d__6_ XI11_1/XI0/XI0_46/d_6_ DECAP_INV_G11
XG13230 XI11_1/XI0/XI0_46/d__5_ XI11_1/XI0/XI0_46/d_5_ DECAP_INV_G11
XG13231 XI11_1/XI0/XI0_46/d__4_ XI11_1/XI0/XI0_46/d_4_ DECAP_INV_G11
XG13232 XI11_1/XI0/XI0_46/d__3_ XI11_1/XI0/XI0_46/d_3_ DECAP_INV_G11
XG13233 XI11_1/XI0/XI0_46/d__2_ XI11_1/XI0/XI0_46/d_2_ DECAP_INV_G11
XG13234 XI11_1/XI0/XI0_46/d__1_ XI11_1/XI0/XI0_46/d_1_ DECAP_INV_G11
XG13235 XI11_1/XI0/XI0_46/d__0_ XI11_1/XI0/XI0_46/d_0_ DECAP_INV_G11
XG13236 XI11_1/XI0/XI0_46/d_15_ XI11_1/XI0/XI0_46/d__15_ DECAP_INV_G11
XG13237 XI11_1/XI0/XI0_46/d_14_ XI11_1/XI0/XI0_46/d__14_ DECAP_INV_G11
XG13238 XI11_1/XI0/XI0_46/d_13_ XI11_1/XI0/XI0_46/d__13_ DECAP_INV_G11
XG13239 XI11_1/XI0/XI0_46/d_12_ XI11_1/XI0/XI0_46/d__12_ DECAP_INV_G11
XG13240 XI11_1/XI0/XI0_46/d_11_ XI11_1/XI0/XI0_46/d__11_ DECAP_INV_G11
XG13241 XI11_1/XI0/XI0_46/d_10_ XI11_1/XI0/XI0_46/d__10_ DECAP_INV_G11
XG13242 XI11_1/XI0/XI0_46/d_9_ XI11_1/XI0/XI0_46/d__9_ DECAP_INV_G11
XG13243 XI11_1/XI0/XI0_46/d_8_ XI11_1/XI0/XI0_46/d__8_ DECAP_INV_G11
XG13244 XI11_1/XI0/XI0_46/d_7_ XI11_1/XI0/XI0_46/d__7_ DECAP_INV_G11
XG13245 XI11_1/XI0/XI0_46/d_6_ XI11_1/XI0/XI0_46/d__6_ DECAP_INV_G11
XG13246 XI11_1/XI0/XI0_46/d_5_ XI11_1/XI0/XI0_46/d__5_ DECAP_INV_G11
XG13247 XI11_1/XI0/XI0_46/d_4_ XI11_1/XI0/XI0_46/d__4_ DECAP_INV_G11
XG13248 XI11_1/XI0/XI0_46/d_3_ XI11_1/XI0/XI0_46/d__3_ DECAP_INV_G11
XG13249 XI11_1/XI0/XI0_46/d_2_ XI11_1/XI0/XI0_46/d__2_ DECAP_INV_G11
XG13250 XI11_1/XI0/XI0_46/d_1_ XI11_1/XI0/XI0_46/d__1_ DECAP_INV_G11
XG13251 XI11_1/XI0/XI0_46/d_0_ XI11_1/XI0/XI0_46/d__0_ DECAP_INV_G11
XG13252 XI11_1/XI0/XI0_45/d__15_ XI11_1/XI0/XI0_45/d_15_ DECAP_INV_G11
XG13253 XI11_1/XI0/XI0_45/d__14_ XI11_1/XI0/XI0_45/d_14_ DECAP_INV_G11
XG13254 XI11_1/XI0/XI0_45/d__13_ XI11_1/XI0/XI0_45/d_13_ DECAP_INV_G11
XG13255 XI11_1/XI0/XI0_45/d__12_ XI11_1/XI0/XI0_45/d_12_ DECAP_INV_G11
XG13256 XI11_1/XI0/XI0_45/d__11_ XI11_1/XI0/XI0_45/d_11_ DECAP_INV_G11
XG13257 XI11_1/XI0/XI0_45/d__10_ XI11_1/XI0/XI0_45/d_10_ DECAP_INV_G11
XG13258 XI11_1/XI0/XI0_45/d__9_ XI11_1/XI0/XI0_45/d_9_ DECAP_INV_G11
XG13259 XI11_1/XI0/XI0_45/d__8_ XI11_1/XI0/XI0_45/d_8_ DECAP_INV_G11
XG13260 XI11_1/XI0/XI0_45/d__7_ XI11_1/XI0/XI0_45/d_7_ DECAP_INV_G11
XG13261 XI11_1/XI0/XI0_45/d__6_ XI11_1/XI0/XI0_45/d_6_ DECAP_INV_G11
XG13262 XI11_1/XI0/XI0_45/d__5_ XI11_1/XI0/XI0_45/d_5_ DECAP_INV_G11
XG13263 XI11_1/XI0/XI0_45/d__4_ XI11_1/XI0/XI0_45/d_4_ DECAP_INV_G11
XG13264 XI11_1/XI0/XI0_45/d__3_ XI11_1/XI0/XI0_45/d_3_ DECAP_INV_G11
XG13265 XI11_1/XI0/XI0_45/d__2_ XI11_1/XI0/XI0_45/d_2_ DECAP_INV_G11
XG13266 XI11_1/XI0/XI0_45/d__1_ XI11_1/XI0/XI0_45/d_1_ DECAP_INV_G11
XG13267 XI11_1/XI0/XI0_45/d__0_ XI11_1/XI0/XI0_45/d_0_ DECAP_INV_G11
XG13268 XI11_1/XI0/XI0_45/d_15_ XI11_1/XI0/XI0_45/d__15_ DECAP_INV_G11
XG13269 XI11_1/XI0/XI0_45/d_14_ XI11_1/XI0/XI0_45/d__14_ DECAP_INV_G11
XG13270 XI11_1/XI0/XI0_45/d_13_ XI11_1/XI0/XI0_45/d__13_ DECAP_INV_G11
XG13271 XI11_1/XI0/XI0_45/d_12_ XI11_1/XI0/XI0_45/d__12_ DECAP_INV_G11
XG13272 XI11_1/XI0/XI0_45/d_11_ XI11_1/XI0/XI0_45/d__11_ DECAP_INV_G11
XG13273 XI11_1/XI0/XI0_45/d_10_ XI11_1/XI0/XI0_45/d__10_ DECAP_INV_G11
XG13274 XI11_1/XI0/XI0_45/d_9_ XI11_1/XI0/XI0_45/d__9_ DECAP_INV_G11
XG13275 XI11_1/XI0/XI0_45/d_8_ XI11_1/XI0/XI0_45/d__8_ DECAP_INV_G11
XG13276 XI11_1/XI0/XI0_45/d_7_ XI11_1/XI0/XI0_45/d__7_ DECAP_INV_G11
XG13277 XI11_1/XI0/XI0_45/d_6_ XI11_1/XI0/XI0_45/d__6_ DECAP_INV_G11
XG13278 XI11_1/XI0/XI0_45/d_5_ XI11_1/XI0/XI0_45/d__5_ DECAP_INV_G11
XG13279 XI11_1/XI0/XI0_45/d_4_ XI11_1/XI0/XI0_45/d__4_ DECAP_INV_G11
XG13280 XI11_1/XI0/XI0_45/d_3_ XI11_1/XI0/XI0_45/d__3_ DECAP_INV_G11
XG13281 XI11_1/XI0/XI0_45/d_2_ XI11_1/XI0/XI0_45/d__2_ DECAP_INV_G11
XG13282 XI11_1/XI0/XI0_45/d_1_ XI11_1/XI0/XI0_45/d__1_ DECAP_INV_G11
XG13283 XI11_1/XI0/XI0_45/d_0_ XI11_1/XI0/XI0_45/d__0_ DECAP_INV_G11
XG13284 XI11_1/XI0/XI0_44/d__15_ XI11_1/XI0/XI0_44/d_15_ DECAP_INV_G11
XG13285 XI11_1/XI0/XI0_44/d__14_ XI11_1/XI0/XI0_44/d_14_ DECAP_INV_G11
XG13286 XI11_1/XI0/XI0_44/d__13_ XI11_1/XI0/XI0_44/d_13_ DECAP_INV_G11
XG13287 XI11_1/XI0/XI0_44/d__12_ XI11_1/XI0/XI0_44/d_12_ DECAP_INV_G11
XG13288 XI11_1/XI0/XI0_44/d__11_ XI11_1/XI0/XI0_44/d_11_ DECAP_INV_G11
XG13289 XI11_1/XI0/XI0_44/d__10_ XI11_1/XI0/XI0_44/d_10_ DECAP_INV_G11
XG13290 XI11_1/XI0/XI0_44/d__9_ XI11_1/XI0/XI0_44/d_9_ DECAP_INV_G11
XG13291 XI11_1/XI0/XI0_44/d__8_ XI11_1/XI0/XI0_44/d_8_ DECAP_INV_G11
XG13292 XI11_1/XI0/XI0_44/d__7_ XI11_1/XI0/XI0_44/d_7_ DECAP_INV_G11
XG13293 XI11_1/XI0/XI0_44/d__6_ XI11_1/XI0/XI0_44/d_6_ DECAP_INV_G11
XG13294 XI11_1/XI0/XI0_44/d__5_ XI11_1/XI0/XI0_44/d_5_ DECAP_INV_G11
XG13295 XI11_1/XI0/XI0_44/d__4_ XI11_1/XI0/XI0_44/d_4_ DECAP_INV_G11
XG13296 XI11_1/XI0/XI0_44/d__3_ XI11_1/XI0/XI0_44/d_3_ DECAP_INV_G11
XG13297 XI11_1/XI0/XI0_44/d__2_ XI11_1/XI0/XI0_44/d_2_ DECAP_INV_G11
XG13298 XI11_1/XI0/XI0_44/d__1_ XI11_1/XI0/XI0_44/d_1_ DECAP_INV_G11
XG13299 XI11_1/XI0/XI0_44/d__0_ XI11_1/XI0/XI0_44/d_0_ DECAP_INV_G11
XG13300 XI11_1/XI0/XI0_44/d_15_ XI11_1/XI0/XI0_44/d__15_ DECAP_INV_G11
XG13301 XI11_1/XI0/XI0_44/d_14_ XI11_1/XI0/XI0_44/d__14_ DECAP_INV_G11
XG13302 XI11_1/XI0/XI0_44/d_13_ XI11_1/XI0/XI0_44/d__13_ DECAP_INV_G11
XG13303 XI11_1/XI0/XI0_44/d_12_ XI11_1/XI0/XI0_44/d__12_ DECAP_INV_G11
XG13304 XI11_1/XI0/XI0_44/d_11_ XI11_1/XI0/XI0_44/d__11_ DECAP_INV_G11
XG13305 XI11_1/XI0/XI0_44/d_10_ XI11_1/XI0/XI0_44/d__10_ DECAP_INV_G11
XG13306 XI11_1/XI0/XI0_44/d_9_ XI11_1/XI0/XI0_44/d__9_ DECAP_INV_G11
XG13307 XI11_1/XI0/XI0_44/d_8_ XI11_1/XI0/XI0_44/d__8_ DECAP_INV_G11
XG13308 XI11_1/XI0/XI0_44/d_7_ XI11_1/XI0/XI0_44/d__7_ DECAP_INV_G11
XG13309 XI11_1/XI0/XI0_44/d_6_ XI11_1/XI0/XI0_44/d__6_ DECAP_INV_G11
XG13310 XI11_1/XI0/XI0_44/d_5_ XI11_1/XI0/XI0_44/d__5_ DECAP_INV_G11
XG13311 XI11_1/XI0/XI0_44/d_4_ XI11_1/XI0/XI0_44/d__4_ DECAP_INV_G11
XG13312 XI11_1/XI0/XI0_44/d_3_ XI11_1/XI0/XI0_44/d__3_ DECAP_INV_G11
XG13313 XI11_1/XI0/XI0_44/d_2_ XI11_1/XI0/XI0_44/d__2_ DECAP_INV_G11
XG13314 XI11_1/XI0/XI0_44/d_1_ XI11_1/XI0/XI0_44/d__1_ DECAP_INV_G11
XG13315 XI11_1/XI0/XI0_44/d_0_ XI11_1/XI0/XI0_44/d__0_ DECAP_INV_G11
XG13316 XI11_1/XI0/XI0_43/d__15_ XI11_1/XI0/XI0_43/d_15_ DECAP_INV_G11
XG13317 XI11_1/XI0/XI0_43/d__14_ XI11_1/XI0/XI0_43/d_14_ DECAP_INV_G11
XG13318 XI11_1/XI0/XI0_43/d__13_ XI11_1/XI0/XI0_43/d_13_ DECAP_INV_G11
XG13319 XI11_1/XI0/XI0_43/d__12_ XI11_1/XI0/XI0_43/d_12_ DECAP_INV_G11
XG13320 XI11_1/XI0/XI0_43/d__11_ XI11_1/XI0/XI0_43/d_11_ DECAP_INV_G11
XG13321 XI11_1/XI0/XI0_43/d__10_ XI11_1/XI0/XI0_43/d_10_ DECAP_INV_G11
XG13322 XI11_1/XI0/XI0_43/d__9_ XI11_1/XI0/XI0_43/d_9_ DECAP_INV_G11
XG13323 XI11_1/XI0/XI0_43/d__8_ XI11_1/XI0/XI0_43/d_8_ DECAP_INV_G11
XG13324 XI11_1/XI0/XI0_43/d__7_ XI11_1/XI0/XI0_43/d_7_ DECAP_INV_G11
XG13325 XI11_1/XI0/XI0_43/d__6_ XI11_1/XI0/XI0_43/d_6_ DECAP_INV_G11
XG13326 XI11_1/XI0/XI0_43/d__5_ XI11_1/XI0/XI0_43/d_5_ DECAP_INV_G11
XG13327 XI11_1/XI0/XI0_43/d__4_ XI11_1/XI0/XI0_43/d_4_ DECAP_INV_G11
XG13328 XI11_1/XI0/XI0_43/d__3_ XI11_1/XI0/XI0_43/d_3_ DECAP_INV_G11
XG13329 XI11_1/XI0/XI0_43/d__2_ XI11_1/XI0/XI0_43/d_2_ DECAP_INV_G11
XG13330 XI11_1/XI0/XI0_43/d__1_ XI11_1/XI0/XI0_43/d_1_ DECAP_INV_G11
XG13331 XI11_1/XI0/XI0_43/d__0_ XI11_1/XI0/XI0_43/d_0_ DECAP_INV_G11
XG13332 XI11_1/XI0/XI0_43/d_15_ XI11_1/XI0/XI0_43/d__15_ DECAP_INV_G11
XG13333 XI11_1/XI0/XI0_43/d_14_ XI11_1/XI0/XI0_43/d__14_ DECAP_INV_G11
XG13334 XI11_1/XI0/XI0_43/d_13_ XI11_1/XI0/XI0_43/d__13_ DECAP_INV_G11
XG13335 XI11_1/XI0/XI0_43/d_12_ XI11_1/XI0/XI0_43/d__12_ DECAP_INV_G11
XG13336 XI11_1/XI0/XI0_43/d_11_ XI11_1/XI0/XI0_43/d__11_ DECAP_INV_G11
XG13337 XI11_1/XI0/XI0_43/d_10_ XI11_1/XI0/XI0_43/d__10_ DECAP_INV_G11
XG13338 XI11_1/XI0/XI0_43/d_9_ XI11_1/XI0/XI0_43/d__9_ DECAP_INV_G11
XG13339 XI11_1/XI0/XI0_43/d_8_ XI11_1/XI0/XI0_43/d__8_ DECAP_INV_G11
XG13340 XI11_1/XI0/XI0_43/d_7_ XI11_1/XI0/XI0_43/d__7_ DECAP_INV_G11
XG13341 XI11_1/XI0/XI0_43/d_6_ XI11_1/XI0/XI0_43/d__6_ DECAP_INV_G11
XG13342 XI11_1/XI0/XI0_43/d_5_ XI11_1/XI0/XI0_43/d__5_ DECAP_INV_G11
XG13343 XI11_1/XI0/XI0_43/d_4_ XI11_1/XI0/XI0_43/d__4_ DECAP_INV_G11
XG13344 XI11_1/XI0/XI0_43/d_3_ XI11_1/XI0/XI0_43/d__3_ DECAP_INV_G11
XG13345 XI11_1/XI0/XI0_43/d_2_ XI11_1/XI0/XI0_43/d__2_ DECAP_INV_G11
XG13346 XI11_1/XI0/XI0_43/d_1_ XI11_1/XI0/XI0_43/d__1_ DECAP_INV_G11
XG13347 XI11_1/XI0/XI0_43/d_0_ XI11_1/XI0/XI0_43/d__0_ DECAP_INV_G11
XG13348 XI11_1/XI0/XI0_42/d__15_ XI11_1/XI0/XI0_42/d_15_ DECAP_INV_G11
XG13349 XI11_1/XI0/XI0_42/d__14_ XI11_1/XI0/XI0_42/d_14_ DECAP_INV_G11
XG13350 XI11_1/XI0/XI0_42/d__13_ XI11_1/XI0/XI0_42/d_13_ DECAP_INV_G11
XG13351 XI11_1/XI0/XI0_42/d__12_ XI11_1/XI0/XI0_42/d_12_ DECAP_INV_G11
XG13352 XI11_1/XI0/XI0_42/d__11_ XI11_1/XI0/XI0_42/d_11_ DECAP_INV_G11
XG13353 XI11_1/XI0/XI0_42/d__10_ XI11_1/XI0/XI0_42/d_10_ DECAP_INV_G11
XG13354 XI11_1/XI0/XI0_42/d__9_ XI11_1/XI0/XI0_42/d_9_ DECAP_INV_G11
XG13355 XI11_1/XI0/XI0_42/d__8_ XI11_1/XI0/XI0_42/d_8_ DECAP_INV_G11
XG13356 XI11_1/XI0/XI0_42/d__7_ XI11_1/XI0/XI0_42/d_7_ DECAP_INV_G11
XG13357 XI11_1/XI0/XI0_42/d__6_ XI11_1/XI0/XI0_42/d_6_ DECAP_INV_G11
XG13358 XI11_1/XI0/XI0_42/d__5_ XI11_1/XI0/XI0_42/d_5_ DECAP_INV_G11
XG13359 XI11_1/XI0/XI0_42/d__4_ XI11_1/XI0/XI0_42/d_4_ DECAP_INV_G11
XG13360 XI11_1/XI0/XI0_42/d__3_ XI11_1/XI0/XI0_42/d_3_ DECAP_INV_G11
XG13361 XI11_1/XI0/XI0_42/d__2_ XI11_1/XI0/XI0_42/d_2_ DECAP_INV_G11
XG13362 XI11_1/XI0/XI0_42/d__1_ XI11_1/XI0/XI0_42/d_1_ DECAP_INV_G11
XG13363 XI11_1/XI0/XI0_42/d__0_ XI11_1/XI0/XI0_42/d_0_ DECAP_INV_G11
XG13364 XI11_1/XI0/XI0_42/d_15_ XI11_1/XI0/XI0_42/d__15_ DECAP_INV_G11
XG13365 XI11_1/XI0/XI0_42/d_14_ XI11_1/XI0/XI0_42/d__14_ DECAP_INV_G11
XG13366 XI11_1/XI0/XI0_42/d_13_ XI11_1/XI0/XI0_42/d__13_ DECAP_INV_G11
XG13367 XI11_1/XI0/XI0_42/d_12_ XI11_1/XI0/XI0_42/d__12_ DECAP_INV_G11
XG13368 XI11_1/XI0/XI0_42/d_11_ XI11_1/XI0/XI0_42/d__11_ DECAP_INV_G11
XG13369 XI11_1/XI0/XI0_42/d_10_ XI11_1/XI0/XI0_42/d__10_ DECAP_INV_G11
XG13370 XI11_1/XI0/XI0_42/d_9_ XI11_1/XI0/XI0_42/d__9_ DECAP_INV_G11
XG13371 XI11_1/XI0/XI0_42/d_8_ XI11_1/XI0/XI0_42/d__8_ DECAP_INV_G11
XG13372 XI11_1/XI0/XI0_42/d_7_ XI11_1/XI0/XI0_42/d__7_ DECAP_INV_G11
XG13373 XI11_1/XI0/XI0_42/d_6_ XI11_1/XI0/XI0_42/d__6_ DECAP_INV_G11
XG13374 XI11_1/XI0/XI0_42/d_5_ XI11_1/XI0/XI0_42/d__5_ DECAP_INV_G11
XG13375 XI11_1/XI0/XI0_42/d_4_ XI11_1/XI0/XI0_42/d__4_ DECAP_INV_G11
XG13376 XI11_1/XI0/XI0_42/d_3_ XI11_1/XI0/XI0_42/d__3_ DECAP_INV_G11
XG13377 XI11_1/XI0/XI0_42/d_2_ XI11_1/XI0/XI0_42/d__2_ DECAP_INV_G11
XG13378 XI11_1/XI0/XI0_42/d_1_ XI11_1/XI0/XI0_42/d__1_ DECAP_INV_G11
XG13379 XI11_1/XI0/XI0_42/d_0_ XI11_1/XI0/XI0_42/d__0_ DECAP_INV_G11
XG13380 XI11_1/XI0/XI0_41/d__15_ XI11_1/XI0/XI0_41/d_15_ DECAP_INV_G11
XG13381 XI11_1/XI0/XI0_41/d__14_ XI11_1/XI0/XI0_41/d_14_ DECAP_INV_G11
XG13382 XI11_1/XI0/XI0_41/d__13_ XI11_1/XI0/XI0_41/d_13_ DECAP_INV_G11
XG13383 XI11_1/XI0/XI0_41/d__12_ XI11_1/XI0/XI0_41/d_12_ DECAP_INV_G11
XG13384 XI11_1/XI0/XI0_41/d__11_ XI11_1/XI0/XI0_41/d_11_ DECAP_INV_G11
XG13385 XI11_1/XI0/XI0_41/d__10_ XI11_1/XI0/XI0_41/d_10_ DECAP_INV_G11
XG13386 XI11_1/XI0/XI0_41/d__9_ XI11_1/XI0/XI0_41/d_9_ DECAP_INV_G11
XG13387 XI11_1/XI0/XI0_41/d__8_ XI11_1/XI0/XI0_41/d_8_ DECAP_INV_G11
XG13388 XI11_1/XI0/XI0_41/d__7_ XI11_1/XI0/XI0_41/d_7_ DECAP_INV_G11
XG13389 XI11_1/XI0/XI0_41/d__6_ XI11_1/XI0/XI0_41/d_6_ DECAP_INV_G11
XG13390 XI11_1/XI0/XI0_41/d__5_ XI11_1/XI0/XI0_41/d_5_ DECAP_INV_G11
XG13391 XI11_1/XI0/XI0_41/d__4_ XI11_1/XI0/XI0_41/d_4_ DECAP_INV_G11
XG13392 XI11_1/XI0/XI0_41/d__3_ XI11_1/XI0/XI0_41/d_3_ DECAP_INV_G11
XG13393 XI11_1/XI0/XI0_41/d__2_ XI11_1/XI0/XI0_41/d_2_ DECAP_INV_G11
XG13394 XI11_1/XI0/XI0_41/d__1_ XI11_1/XI0/XI0_41/d_1_ DECAP_INV_G11
XG13395 XI11_1/XI0/XI0_41/d__0_ XI11_1/XI0/XI0_41/d_0_ DECAP_INV_G11
XG13396 XI11_1/XI0/XI0_41/d_15_ XI11_1/XI0/XI0_41/d__15_ DECAP_INV_G11
XG13397 XI11_1/XI0/XI0_41/d_14_ XI11_1/XI0/XI0_41/d__14_ DECAP_INV_G11
XG13398 XI11_1/XI0/XI0_41/d_13_ XI11_1/XI0/XI0_41/d__13_ DECAP_INV_G11
XG13399 XI11_1/XI0/XI0_41/d_12_ XI11_1/XI0/XI0_41/d__12_ DECAP_INV_G11
XG13400 XI11_1/XI0/XI0_41/d_11_ XI11_1/XI0/XI0_41/d__11_ DECAP_INV_G11
XG13401 XI11_1/XI0/XI0_41/d_10_ XI11_1/XI0/XI0_41/d__10_ DECAP_INV_G11
XG13402 XI11_1/XI0/XI0_41/d_9_ XI11_1/XI0/XI0_41/d__9_ DECAP_INV_G11
XG13403 XI11_1/XI0/XI0_41/d_8_ XI11_1/XI0/XI0_41/d__8_ DECAP_INV_G11
XG13404 XI11_1/XI0/XI0_41/d_7_ XI11_1/XI0/XI0_41/d__7_ DECAP_INV_G11
XG13405 XI11_1/XI0/XI0_41/d_6_ XI11_1/XI0/XI0_41/d__6_ DECAP_INV_G11
XG13406 XI11_1/XI0/XI0_41/d_5_ XI11_1/XI0/XI0_41/d__5_ DECAP_INV_G11
XG13407 XI11_1/XI0/XI0_41/d_4_ XI11_1/XI0/XI0_41/d__4_ DECAP_INV_G11
XG13408 XI11_1/XI0/XI0_41/d_3_ XI11_1/XI0/XI0_41/d__3_ DECAP_INV_G11
XG13409 XI11_1/XI0/XI0_41/d_2_ XI11_1/XI0/XI0_41/d__2_ DECAP_INV_G11
XG13410 XI11_1/XI0/XI0_41/d_1_ XI11_1/XI0/XI0_41/d__1_ DECAP_INV_G11
XG13411 XI11_1/XI0/XI0_41/d_0_ XI11_1/XI0/XI0_41/d__0_ DECAP_INV_G11
XG13412 XI11_1/XI0/XI0_40/d__15_ XI11_1/XI0/XI0_40/d_15_ DECAP_INV_G11
XG13413 XI11_1/XI0/XI0_40/d__14_ XI11_1/XI0/XI0_40/d_14_ DECAP_INV_G11
XG13414 XI11_1/XI0/XI0_40/d__13_ XI11_1/XI0/XI0_40/d_13_ DECAP_INV_G11
XG13415 XI11_1/XI0/XI0_40/d__12_ XI11_1/XI0/XI0_40/d_12_ DECAP_INV_G11
XG13416 XI11_1/XI0/XI0_40/d__11_ XI11_1/XI0/XI0_40/d_11_ DECAP_INV_G11
XG13417 XI11_1/XI0/XI0_40/d__10_ XI11_1/XI0/XI0_40/d_10_ DECAP_INV_G11
XG13418 XI11_1/XI0/XI0_40/d__9_ XI11_1/XI0/XI0_40/d_9_ DECAP_INV_G11
XG13419 XI11_1/XI0/XI0_40/d__8_ XI11_1/XI0/XI0_40/d_8_ DECAP_INV_G11
XG13420 XI11_1/XI0/XI0_40/d__7_ XI11_1/XI0/XI0_40/d_7_ DECAP_INV_G11
XG13421 XI11_1/XI0/XI0_40/d__6_ XI11_1/XI0/XI0_40/d_6_ DECAP_INV_G11
XG13422 XI11_1/XI0/XI0_40/d__5_ XI11_1/XI0/XI0_40/d_5_ DECAP_INV_G11
XG13423 XI11_1/XI0/XI0_40/d__4_ XI11_1/XI0/XI0_40/d_4_ DECAP_INV_G11
XG13424 XI11_1/XI0/XI0_40/d__3_ XI11_1/XI0/XI0_40/d_3_ DECAP_INV_G11
XG13425 XI11_1/XI0/XI0_40/d__2_ XI11_1/XI0/XI0_40/d_2_ DECAP_INV_G11
XG13426 XI11_1/XI0/XI0_40/d__1_ XI11_1/XI0/XI0_40/d_1_ DECAP_INV_G11
XG13427 XI11_1/XI0/XI0_40/d__0_ XI11_1/XI0/XI0_40/d_0_ DECAP_INV_G11
XG13428 XI11_1/XI0/XI0_40/d_15_ XI11_1/XI0/XI0_40/d__15_ DECAP_INV_G11
XG13429 XI11_1/XI0/XI0_40/d_14_ XI11_1/XI0/XI0_40/d__14_ DECAP_INV_G11
XG13430 XI11_1/XI0/XI0_40/d_13_ XI11_1/XI0/XI0_40/d__13_ DECAP_INV_G11
XG13431 XI11_1/XI0/XI0_40/d_12_ XI11_1/XI0/XI0_40/d__12_ DECAP_INV_G11
XG13432 XI11_1/XI0/XI0_40/d_11_ XI11_1/XI0/XI0_40/d__11_ DECAP_INV_G11
XG13433 XI11_1/XI0/XI0_40/d_10_ XI11_1/XI0/XI0_40/d__10_ DECAP_INV_G11
XG13434 XI11_1/XI0/XI0_40/d_9_ XI11_1/XI0/XI0_40/d__9_ DECAP_INV_G11
XG13435 XI11_1/XI0/XI0_40/d_8_ XI11_1/XI0/XI0_40/d__8_ DECAP_INV_G11
XG13436 XI11_1/XI0/XI0_40/d_7_ XI11_1/XI0/XI0_40/d__7_ DECAP_INV_G11
XG13437 XI11_1/XI0/XI0_40/d_6_ XI11_1/XI0/XI0_40/d__6_ DECAP_INV_G11
XG13438 XI11_1/XI0/XI0_40/d_5_ XI11_1/XI0/XI0_40/d__5_ DECAP_INV_G11
XG13439 XI11_1/XI0/XI0_40/d_4_ XI11_1/XI0/XI0_40/d__4_ DECAP_INV_G11
XG13440 XI11_1/XI0/XI0_40/d_3_ XI11_1/XI0/XI0_40/d__3_ DECAP_INV_G11
XG13441 XI11_1/XI0/XI0_40/d_2_ XI11_1/XI0/XI0_40/d__2_ DECAP_INV_G11
XG13442 XI11_1/XI0/XI0_40/d_1_ XI11_1/XI0/XI0_40/d__1_ DECAP_INV_G11
XG13443 XI11_1/XI0/XI0_40/d_0_ XI11_1/XI0/XI0_40/d__0_ DECAP_INV_G11
XG13444 XI11_1/XI0/XI0_39/d__15_ XI11_1/XI0/XI0_39/d_15_ DECAP_INV_G11
XG13445 XI11_1/XI0/XI0_39/d__14_ XI11_1/XI0/XI0_39/d_14_ DECAP_INV_G11
XG13446 XI11_1/XI0/XI0_39/d__13_ XI11_1/XI0/XI0_39/d_13_ DECAP_INV_G11
XG13447 XI11_1/XI0/XI0_39/d__12_ XI11_1/XI0/XI0_39/d_12_ DECAP_INV_G11
XG13448 XI11_1/XI0/XI0_39/d__11_ XI11_1/XI0/XI0_39/d_11_ DECAP_INV_G11
XG13449 XI11_1/XI0/XI0_39/d__10_ XI11_1/XI0/XI0_39/d_10_ DECAP_INV_G11
XG13450 XI11_1/XI0/XI0_39/d__9_ XI11_1/XI0/XI0_39/d_9_ DECAP_INV_G11
XG13451 XI11_1/XI0/XI0_39/d__8_ XI11_1/XI0/XI0_39/d_8_ DECAP_INV_G11
XG13452 XI11_1/XI0/XI0_39/d__7_ XI11_1/XI0/XI0_39/d_7_ DECAP_INV_G11
XG13453 XI11_1/XI0/XI0_39/d__6_ XI11_1/XI0/XI0_39/d_6_ DECAP_INV_G11
XG13454 XI11_1/XI0/XI0_39/d__5_ XI11_1/XI0/XI0_39/d_5_ DECAP_INV_G11
XG13455 XI11_1/XI0/XI0_39/d__4_ XI11_1/XI0/XI0_39/d_4_ DECAP_INV_G11
XG13456 XI11_1/XI0/XI0_39/d__3_ XI11_1/XI0/XI0_39/d_3_ DECAP_INV_G11
XG13457 XI11_1/XI0/XI0_39/d__2_ XI11_1/XI0/XI0_39/d_2_ DECAP_INV_G11
XG13458 XI11_1/XI0/XI0_39/d__1_ XI11_1/XI0/XI0_39/d_1_ DECAP_INV_G11
XG13459 XI11_1/XI0/XI0_39/d__0_ XI11_1/XI0/XI0_39/d_0_ DECAP_INV_G11
XG13460 XI11_1/XI0/XI0_39/d_15_ XI11_1/XI0/XI0_39/d__15_ DECAP_INV_G11
XG13461 XI11_1/XI0/XI0_39/d_14_ XI11_1/XI0/XI0_39/d__14_ DECAP_INV_G11
XG13462 XI11_1/XI0/XI0_39/d_13_ XI11_1/XI0/XI0_39/d__13_ DECAP_INV_G11
XG13463 XI11_1/XI0/XI0_39/d_12_ XI11_1/XI0/XI0_39/d__12_ DECAP_INV_G11
XG13464 XI11_1/XI0/XI0_39/d_11_ XI11_1/XI0/XI0_39/d__11_ DECAP_INV_G11
XG13465 XI11_1/XI0/XI0_39/d_10_ XI11_1/XI0/XI0_39/d__10_ DECAP_INV_G11
XG13466 XI11_1/XI0/XI0_39/d_9_ XI11_1/XI0/XI0_39/d__9_ DECAP_INV_G11
XG13467 XI11_1/XI0/XI0_39/d_8_ XI11_1/XI0/XI0_39/d__8_ DECAP_INV_G11
XG13468 XI11_1/XI0/XI0_39/d_7_ XI11_1/XI0/XI0_39/d__7_ DECAP_INV_G11
XG13469 XI11_1/XI0/XI0_39/d_6_ XI11_1/XI0/XI0_39/d__6_ DECAP_INV_G11
XG13470 XI11_1/XI0/XI0_39/d_5_ XI11_1/XI0/XI0_39/d__5_ DECAP_INV_G11
XG13471 XI11_1/XI0/XI0_39/d_4_ XI11_1/XI0/XI0_39/d__4_ DECAP_INV_G11
XG13472 XI11_1/XI0/XI0_39/d_3_ XI11_1/XI0/XI0_39/d__3_ DECAP_INV_G11
XG13473 XI11_1/XI0/XI0_39/d_2_ XI11_1/XI0/XI0_39/d__2_ DECAP_INV_G11
XG13474 XI11_1/XI0/XI0_39/d_1_ XI11_1/XI0/XI0_39/d__1_ DECAP_INV_G11
XG13475 XI11_1/XI0/XI0_39/d_0_ XI11_1/XI0/XI0_39/d__0_ DECAP_INV_G11
XG13476 XI11_1/XI0/XI0_38/d__15_ XI11_1/XI0/XI0_38/d_15_ DECAP_INV_G11
XG13477 XI11_1/XI0/XI0_38/d__14_ XI11_1/XI0/XI0_38/d_14_ DECAP_INV_G11
XG13478 XI11_1/XI0/XI0_38/d__13_ XI11_1/XI0/XI0_38/d_13_ DECAP_INV_G11
XG13479 XI11_1/XI0/XI0_38/d__12_ XI11_1/XI0/XI0_38/d_12_ DECAP_INV_G11
XG13480 XI11_1/XI0/XI0_38/d__11_ XI11_1/XI0/XI0_38/d_11_ DECAP_INV_G11
XG13481 XI11_1/XI0/XI0_38/d__10_ XI11_1/XI0/XI0_38/d_10_ DECAP_INV_G11
XG13482 XI11_1/XI0/XI0_38/d__9_ XI11_1/XI0/XI0_38/d_9_ DECAP_INV_G11
XG13483 XI11_1/XI0/XI0_38/d__8_ XI11_1/XI0/XI0_38/d_8_ DECAP_INV_G11
XG13484 XI11_1/XI0/XI0_38/d__7_ XI11_1/XI0/XI0_38/d_7_ DECAP_INV_G11
XG13485 XI11_1/XI0/XI0_38/d__6_ XI11_1/XI0/XI0_38/d_6_ DECAP_INV_G11
XG13486 XI11_1/XI0/XI0_38/d__5_ XI11_1/XI0/XI0_38/d_5_ DECAP_INV_G11
XG13487 XI11_1/XI0/XI0_38/d__4_ XI11_1/XI0/XI0_38/d_4_ DECAP_INV_G11
XG13488 XI11_1/XI0/XI0_38/d__3_ XI11_1/XI0/XI0_38/d_3_ DECAP_INV_G11
XG13489 XI11_1/XI0/XI0_38/d__2_ XI11_1/XI0/XI0_38/d_2_ DECAP_INV_G11
XG13490 XI11_1/XI0/XI0_38/d__1_ XI11_1/XI0/XI0_38/d_1_ DECAP_INV_G11
XG13491 XI11_1/XI0/XI0_38/d__0_ XI11_1/XI0/XI0_38/d_0_ DECAP_INV_G11
XG13492 XI11_1/XI0/XI0_38/d_15_ XI11_1/XI0/XI0_38/d__15_ DECAP_INV_G11
XG13493 XI11_1/XI0/XI0_38/d_14_ XI11_1/XI0/XI0_38/d__14_ DECAP_INV_G11
XG13494 XI11_1/XI0/XI0_38/d_13_ XI11_1/XI0/XI0_38/d__13_ DECAP_INV_G11
XG13495 XI11_1/XI0/XI0_38/d_12_ XI11_1/XI0/XI0_38/d__12_ DECAP_INV_G11
XG13496 XI11_1/XI0/XI0_38/d_11_ XI11_1/XI0/XI0_38/d__11_ DECAP_INV_G11
XG13497 XI11_1/XI0/XI0_38/d_10_ XI11_1/XI0/XI0_38/d__10_ DECAP_INV_G11
XG13498 XI11_1/XI0/XI0_38/d_9_ XI11_1/XI0/XI0_38/d__9_ DECAP_INV_G11
XG13499 XI11_1/XI0/XI0_38/d_8_ XI11_1/XI0/XI0_38/d__8_ DECAP_INV_G11
XG13500 XI11_1/XI0/XI0_38/d_7_ XI11_1/XI0/XI0_38/d__7_ DECAP_INV_G11
XG13501 XI11_1/XI0/XI0_38/d_6_ XI11_1/XI0/XI0_38/d__6_ DECAP_INV_G11
XG13502 XI11_1/XI0/XI0_38/d_5_ XI11_1/XI0/XI0_38/d__5_ DECAP_INV_G11
XG13503 XI11_1/XI0/XI0_38/d_4_ XI11_1/XI0/XI0_38/d__4_ DECAP_INV_G11
XG13504 XI11_1/XI0/XI0_38/d_3_ XI11_1/XI0/XI0_38/d__3_ DECAP_INV_G11
XG13505 XI11_1/XI0/XI0_38/d_2_ XI11_1/XI0/XI0_38/d__2_ DECAP_INV_G11
XG13506 XI11_1/XI0/XI0_38/d_1_ XI11_1/XI0/XI0_38/d__1_ DECAP_INV_G11
XG13507 XI11_1/XI0/XI0_38/d_0_ XI11_1/XI0/XI0_38/d__0_ DECAP_INV_G11
XG13508 XI11_1/XI0/XI0_37/d__15_ XI11_1/XI0/XI0_37/d_15_ DECAP_INV_G11
XG13509 XI11_1/XI0/XI0_37/d__14_ XI11_1/XI0/XI0_37/d_14_ DECAP_INV_G11
XG13510 XI11_1/XI0/XI0_37/d__13_ XI11_1/XI0/XI0_37/d_13_ DECAP_INV_G11
XG13511 XI11_1/XI0/XI0_37/d__12_ XI11_1/XI0/XI0_37/d_12_ DECAP_INV_G11
XG13512 XI11_1/XI0/XI0_37/d__11_ XI11_1/XI0/XI0_37/d_11_ DECAP_INV_G11
XG13513 XI11_1/XI0/XI0_37/d__10_ XI11_1/XI0/XI0_37/d_10_ DECAP_INV_G11
XG13514 XI11_1/XI0/XI0_37/d__9_ XI11_1/XI0/XI0_37/d_9_ DECAP_INV_G11
XG13515 XI11_1/XI0/XI0_37/d__8_ XI11_1/XI0/XI0_37/d_8_ DECAP_INV_G11
XG13516 XI11_1/XI0/XI0_37/d__7_ XI11_1/XI0/XI0_37/d_7_ DECAP_INV_G11
XG13517 XI11_1/XI0/XI0_37/d__6_ XI11_1/XI0/XI0_37/d_6_ DECAP_INV_G11
XG13518 XI11_1/XI0/XI0_37/d__5_ XI11_1/XI0/XI0_37/d_5_ DECAP_INV_G11
XG13519 XI11_1/XI0/XI0_37/d__4_ XI11_1/XI0/XI0_37/d_4_ DECAP_INV_G11
XG13520 XI11_1/XI0/XI0_37/d__3_ XI11_1/XI0/XI0_37/d_3_ DECAP_INV_G11
XG13521 XI11_1/XI0/XI0_37/d__2_ XI11_1/XI0/XI0_37/d_2_ DECAP_INV_G11
XG13522 XI11_1/XI0/XI0_37/d__1_ XI11_1/XI0/XI0_37/d_1_ DECAP_INV_G11
XG13523 XI11_1/XI0/XI0_37/d__0_ XI11_1/XI0/XI0_37/d_0_ DECAP_INV_G11
XG13524 XI11_1/XI0/XI0_37/d_15_ XI11_1/XI0/XI0_37/d__15_ DECAP_INV_G11
XG13525 XI11_1/XI0/XI0_37/d_14_ XI11_1/XI0/XI0_37/d__14_ DECAP_INV_G11
XG13526 XI11_1/XI0/XI0_37/d_13_ XI11_1/XI0/XI0_37/d__13_ DECAP_INV_G11
XG13527 XI11_1/XI0/XI0_37/d_12_ XI11_1/XI0/XI0_37/d__12_ DECAP_INV_G11
XG13528 XI11_1/XI0/XI0_37/d_11_ XI11_1/XI0/XI0_37/d__11_ DECAP_INV_G11
XG13529 XI11_1/XI0/XI0_37/d_10_ XI11_1/XI0/XI0_37/d__10_ DECAP_INV_G11
XG13530 XI11_1/XI0/XI0_37/d_9_ XI11_1/XI0/XI0_37/d__9_ DECAP_INV_G11
XG13531 XI11_1/XI0/XI0_37/d_8_ XI11_1/XI0/XI0_37/d__8_ DECAP_INV_G11
XG13532 XI11_1/XI0/XI0_37/d_7_ XI11_1/XI0/XI0_37/d__7_ DECAP_INV_G11
XG13533 XI11_1/XI0/XI0_37/d_6_ XI11_1/XI0/XI0_37/d__6_ DECAP_INV_G11
XG13534 XI11_1/XI0/XI0_37/d_5_ XI11_1/XI0/XI0_37/d__5_ DECAP_INV_G11
XG13535 XI11_1/XI0/XI0_37/d_4_ XI11_1/XI0/XI0_37/d__4_ DECAP_INV_G11
XG13536 XI11_1/XI0/XI0_37/d_3_ XI11_1/XI0/XI0_37/d__3_ DECAP_INV_G11
XG13537 XI11_1/XI0/XI0_37/d_2_ XI11_1/XI0/XI0_37/d__2_ DECAP_INV_G11
XG13538 XI11_1/XI0/XI0_37/d_1_ XI11_1/XI0/XI0_37/d__1_ DECAP_INV_G11
XG13539 XI11_1/XI0/XI0_37/d_0_ XI11_1/XI0/XI0_37/d__0_ DECAP_INV_G11
XG13540 XI11_1/XI0/XI0_36/d__15_ XI11_1/XI0/XI0_36/d_15_ DECAP_INV_G11
XG13541 XI11_1/XI0/XI0_36/d__14_ XI11_1/XI0/XI0_36/d_14_ DECAP_INV_G11
XG13542 XI11_1/XI0/XI0_36/d__13_ XI11_1/XI0/XI0_36/d_13_ DECAP_INV_G11
XG13543 XI11_1/XI0/XI0_36/d__12_ XI11_1/XI0/XI0_36/d_12_ DECAP_INV_G11
XG13544 XI11_1/XI0/XI0_36/d__11_ XI11_1/XI0/XI0_36/d_11_ DECAP_INV_G11
XG13545 XI11_1/XI0/XI0_36/d__10_ XI11_1/XI0/XI0_36/d_10_ DECAP_INV_G11
XG13546 XI11_1/XI0/XI0_36/d__9_ XI11_1/XI0/XI0_36/d_9_ DECAP_INV_G11
XG13547 XI11_1/XI0/XI0_36/d__8_ XI11_1/XI0/XI0_36/d_8_ DECAP_INV_G11
XG13548 XI11_1/XI0/XI0_36/d__7_ XI11_1/XI0/XI0_36/d_7_ DECAP_INV_G11
XG13549 XI11_1/XI0/XI0_36/d__6_ XI11_1/XI0/XI0_36/d_6_ DECAP_INV_G11
XG13550 XI11_1/XI0/XI0_36/d__5_ XI11_1/XI0/XI0_36/d_5_ DECAP_INV_G11
XG13551 XI11_1/XI0/XI0_36/d__4_ XI11_1/XI0/XI0_36/d_4_ DECAP_INV_G11
XG13552 XI11_1/XI0/XI0_36/d__3_ XI11_1/XI0/XI0_36/d_3_ DECAP_INV_G11
XG13553 XI11_1/XI0/XI0_36/d__2_ XI11_1/XI0/XI0_36/d_2_ DECAP_INV_G11
XG13554 XI11_1/XI0/XI0_36/d__1_ XI11_1/XI0/XI0_36/d_1_ DECAP_INV_G11
XG13555 XI11_1/XI0/XI0_36/d__0_ XI11_1/XI0/XI0_36/d_0_ DECAP_INV_G11
XG13556 XI11_1/XI0/XI0_36/d_15_ XI11_1/XI0/XI0_36/d__15_ DECAP_INV_G11
XG13557 XI11_1/XI0/XI0_36/d_14_ XI11_1/XI0/XI0_36/d__14_ DECAP_INV_G11
XG13558 XI11_1/XI0/XI0_36/d_13_ XI11_1/XI0/XI0_36/d__13_ DECAP_INV_G11
XG13559 XI11_1/XI0/XI0_36/d_12_ XI11_1/XI0/XI0_36/d__12_ DECAP_INV_G11
XG13560 XI11_1/XI0/XI0_36/d_11_ XI11_1/XI0/XI0_36/d__11_ DECAP_INV_G11
XG13561 XI11_1/XI0/XI0_36/d_10_ XI11_1/XI0/XI0_36/d__10_ DECAP_INV_G11
XG13562 XI11_1/XI0/XI0_36/d_9_ XI11_1/XI0/XI0_36/d__9_ DECAP_INV_G11
XG13563 XI11_1/XI0/XI0_36/d_8_ XI11_1/XI0/XI0_36/d__8_ DECAP_INV_G11
XG13564 XI11_1/XI0/XI0_36/d_7_ XI11_1/XI0/XI0_36/d__7_ DECAP_INV_G11
XG13565 XI11_1/XI0/XI0_36/d_6_ XI11_1/XI0/XI0_36/d__6_ DECAP_INV_G11
XG13566 XI11_1/XI0/XI0_36/d_5_ XI11_1/XI0/XI0_36/d__5_ DECAP_INV_G11
XG13567 XI11_1/XI0/XI0_36/d_4_ XI11_1/XI0/XI0_36/d__4_ DECAP_INV_G11
XG13568 XI11_1/XI0/XI0_36/d_3_ XI11_1/XI0/XI0_36/d__3_ DECAP_INV_G11
XG13569 XI11_1/XI0/XI0_36/d_2_ XI11_1/XI0/XI0_36/d__2_ DECAP_INV_G11
XG13570 XI11_1/XI0/XI0_36/d_1_ XI11_1/XI0/XI0_36/d__1_ DECAP_INV_G11
XG13571 XI11_1/XI0/XI0_36/d_0_ XI11_1/XI0/XI0_36/d__0_ DECAP_INV_G11
XG13572 XI11_1/XI0/XI0_35/d__15_ XI11_1/XI0/XI0_35/d_15_ DECAP_INV_G11
XG13573 XI11_1/XI0/XI0_35/d__14_ XI11_1/XI0/XI0_35/d_14_ DECAP_INV_G11
XG13574 XI11_1/XI0/XI0_35/d__13_ XI11_1/XI0/XI0_35/d_13_ DECAP_INV_G11
XG13575 XI11_1/XI0/XI0_35/d__12_ XI11_1/XI0/XI0_35/d_12_ DECAP_INV_G11
XG13576 XI11_1/XI0/XI0_35/d__11_ XI11_1/XI0/XI0_35/d_11_ DECAP_INV_G11
XG13577 XI11_1/XI0/XI0_35/d__10_ XI11_1/XI0/XI0_35/d_10_ DECAP_INV_G11
XG13578 XI11_1/XI0/XI0_35/d__9_ XI11_1/XI0/XI0_35/d_9_ DECAP_INV_G11
XG13579 XI11_1/XI0/XI0_35/d__8_ XI11_1/XI0/XI0_35/d_8_ DECAP_INV_G11
XG13580 XI11_1/XI0/XI0_35/d__7_ XI11_1/XI0/XI0_35/d_7_ DECAP_INV_G11
XG13581 XI11_1/XI0/XI0_35/d__6_ XI11_1/XI0/XI0_35/d_6_ DECAP_INV_G11
XG13582 XI11_1/XI0/XI0_35/d__5_ XI11_1/XI0/XI0_35/d_5_ DECAP_INV_G11
XG13583 XI11_1/XI0/XI0_35/d__4_ XI11_1/XI0/XI0_35/d_4_ DECAP_INV_G11
XG13584 XI11_1/XI0/XI0_35/d__3_ XI11_1/XI0/XI0_35/d_3_ DECAP_INV_G11
XG13585 XI11_1/XI0/XI0_35/d__2_ XI11_1/XI0/XI0_35/d_2_ DECAP_INV_G11
XG13586 XI11_1/XI0/XI0_35/d__1_ XI11_1/XI0/XI0_35/d_1_ DECAP_INV_G11
XG13587 XI11_1/XI0/XI0_35/d__0_ XI11_1/XI0/XI0_35/d_0_ DECAP_INV_G11
XG13588 XI11_1/XI0/XI0_35/d_15_ XI11_1/XI0/XI0_35/d__15_ DECAP_INV_G11
XG13589 XI11_1/XI0/XI0_35/d_14_ XI11_1/XI0/XI0_35/d__14_ DECAP_INV_G11
XG13590 XI11_1/XI0/XI0_35/d_13_ XI11_1/XI0/XI0_35/d__13_ DECAP_INV_G11
XG13591 XI11_1/XI0/XI0_35/d_12_ XI11_1/XI0/XI0_35/d__12_ DECAP_INV_G11
XG13592 XI11_1/XI0/XI0_35/d_11_ XI11_1/XI0/XI0_35/d__11_ DECAP_INV_G11
XG13593 XI11_1/XI0/XI0_35/d_10_ XI11_1/XI0/XI0_35/d__10_ DECAP_INV_G11
XG13594 XI11_1/XI0/XI0_35/d_9_ XI11_1/XI0/XI0_35/d__9_ DECAP_INV_G11
XG13595 XI11_1/XI0/XI0_35/d_8_ XI11_1/XI0/XI0_35/d__8_ DECAP_INV_G11
XG13596 XI11_1/XI0/XI0_35/d_7_ XI11_1/XI0/XI0_35/d__7_ DECAP_INV_G11
XG13597 XI11_1/XI0/XI0_35/d_6_ XI11_1/XI0/XI0_35/d__6_ DECAP_INV_G11
XG13598 XI11_1/XI0/XI0_35/d_5_ XI11_1/XI0/XI0_35/d__5_ DECAP_INV_G11
XG13599 XI11_1/XI0/XI0_35/d_4_ XI11_1/XI0/XI0_35/d__4_ DECAP_INV_G11
XG13600 XI11_1/XI0/XI0_35/d_3_ XI11_1/XI0/XI0_35/d__3_ DECAP_INV_G11
XG13601 XI11_1/XI0/XI0_35/d_2_ XI11_1/XI0/XI0_35/d__2_ DECAP_INV_G11
XG13602 XI11_1/XI0/XI0_35/d_1_ XI11_1/XI0/XI0_35/d__1_ DECAP_INV_G11
XG13603 XI11_1/XI0/XI0_35/d_0_ XI11_1/XI0/XI0_35/d__0_ DECAP_INV_G11
XG13604 XI11_1/XI0/XI0_34/d__15_ XI11_1/XI0/XI0_34/d_15_ DECAP_INV_G11
XG13605 XI11_1/XI0/XI0_34/d__14_ XI11_1/XI0/XI0_34/d_14_ DECAP_INV_G11
XG13606 XI11_1/XI0/XI0_34/d__13_ XI11_1/XI0/XI0_34/d_13_ DECAP_INV_G11
XG13607 XI11_1/XI0/XI0_34/d__12_ XI11_1/XI0/XI0_34/d_12_ DECAP_INV_G11
XG13608 XI11_1/XI0/XI0_34/d__11_ XI11_1/XI0/XI0_34/d_11_ DECAP_INV_G11
XG13609 XI11_1/XI0/XI0_34/d__10_ XI11_1/XI0/XI0_34/d_10_ DECAP_INV_G11
XG13610 XI11_1/XI0/XI0_34/d__9_ XI11_1/XI0/XI0_34/d_9_ DECAP_INV_G11
XG13611 XI11_1/XI0/XI0_34/d__8_ XI11_1/XI0/XI0_34/d_8_ DECAP_INV_G11
XG13612 XI11_1/XI0/XI0_34/d__7_ XI11_1/XI0/XI0_34/d_7_ DECAP_INV_G11
XG13613 XI11_1/XI0/XI0_34/d__6_ XI11_1/XI0/XI0_34/d_6_ DECAP_INV_G11
XG13614 XI11_1/XI0/XI0_34/d__5_ XI11_1/XI0/XI0_34/d_5_ DECAP_INV_G11
XG13615 XI11_1/XI0/XI0_34/d__4_ XI11_1/XI0/XI0_34/d_4_ DECAP_INV_G11
XG13616 XI11_1/XI0/XI0_34/d__3_ XI11_1/XI0/XI0_34/d_3_ DECAP_INV_G11
XG13617 XI11_1/XI0/XI0_34/d__2_ XI11_1/XI0/XI0_34/d_2_ DECAP_INV_G11
XG13618 XI11_1/XI0/XI0_34/d__1_ XI11_1/XI0/XI0_34/d_1_ DECAP_INV_G11
XG13619 XI11_1/XI0/XI0_34/d__0_ XI11_1/XI0/XI0_34/d_0_ DECAP_INV_G11
XG13620 XI11_1/XI0/XI0_34/d_15_ XI11_1/XI0/XI0_34/d__15_ DECAP_INV_G11
XG13621 XI11_1/XI0/XI0_34/d_14_ XI11_1/XI0/XI0_34/d__14_ DECAP_INV_G11
XG13622 XI11_1/XI0/XI0_34/d_13_ XI11_1/XI0/XI0_34/d__13_ DECAP_INV_G11
XG13623 XI11_1/XI0/XI0_34/d_12_ XI11_1/XI0/XI0_34/d__12_ DECAP_INV_G11
XG13624 XI11_1/XI0/XI0_34/d_11_ XI11_1/XI0/XI0_34/d__11_ DECAP_INV_G11
XG13625 XI11_1/XI0/XI0_34/d_10_ XI11_1/XI0/XI0_34/d__10_ DECAP_INV_G11
XG13626 XI11_1/XI0/XI0_34/d_9_ XI11_1/XI0/XI0_34/d__9_ DECAP_INV_G11
XG13627 XI11_1/XI0/XI0_34/d_8_ XI11_1/XI0/XI0_34/d__8_ DECAP_INV_G11
XG13628 XI11_1/XI0/XI0_34/d_7_ XI11_1/XI0/XI0_34/d__7_ DECAP_INV_G11
XG13629 XI11_1/XI0/XI0_34/d_6_ XI11_1/XI0/XI0_34/d__6_ DECAP_INV_G11
XG13630 XI11_1/XI0/XI0_34/d_5_ XI11_1/XI0/XI0_34/d__5_ DECAP_INV_G11
XG13631 XI11_1/XI0/XI0_34/d_4_ XI11_1/XI0/XI0_34/d__4_ DECAP_INV_G11
XG13632 XI11_1/XI0/XI0_34/d_3_ XI11_1/XI0/XI0_34/d__3_ DECAP_INV_G11
XG13633 XI11_1/XI0/XI0_34/d_2_ XI11_1/XI0/XI0_34/d__2_ DECAP_INV_G11
XG13634 XI11_1/XI0/XI0_34/d_1_ XI11_1/XI0/XI0_34/d__1_ DECAP_INV_G11
XG13635 XI11_1/XI0/XI0_34/d_0_ XI11_1/XI0/XI0_34/d__0_ DECAP_INV_G11
XG13636 XI11_1/XI0/XI0_33/d__15_ XI11_1/XI0/XI0_33/d_15_ DECAP_INV_G11
XG13637 XI11_1/XI0/XI0_33/d__14_ XI11_1/XI0/XI0_33/d_14_ DECAP_INV_G11
XG13638 XI11_1/XI0/XI0_33/d__13_ XI11_1/XI0/XI0_33/d_13_ DECAP_INV_G11
XG13639 XI11_1/XI0/XI0_33/d__12_ XI11_1/XI0/XI0_33/d_12_ DECAP_INV_G11
XG13640 XI11_1/XI0/XI0_33/d__11_ XI11_1/XI0/XI0_33/d_11_ DECAP_INV_G11
XG13641 XI11_1/XI0/XI0_33/d__10_ XI11_1/XI0/XI0_33/d_10_ DECAP_INV_G11
XG13642 XI11_1/XI0/XI0_33/d__9_ XI11_1/XI0/XI0_33/d_9_ DECAP_INV_G11
XG13643 XI11_1/XI0/XI0_33/d__8_ XI11_1/XI0/XI0_33/d_8_ DECAP_INV_G11
XG13644 XI11_1/XI0/XI0_33/d__7_ XI11_1/XI0/XI0_33/d_7_ DECAP_INV_G11
XG13645 XI11_1/XI0/XI0_33/d__6_ XI11_1/XI0/XI0_33/d_6_ DECAP_INV_G11
XG13646 XI11_1/XI0/XI0_33/d__5_ XI11_1/XI0/XI0_33/d_5_ DECAP_INV_G11
XG13647 XI11_1/XI0/XI0_33/d__4_ XI11_1/XI0/XI0_33/d_4_ DECAP_INV_G11
XG13648 XI11_1/XI0/XI0_33/d__3_ XI11_1/XI0/XI0_33/d_3_ DECAP_INV_G11
XG13649 XI11_1/XI0/XI0_33/d__2_ XI11_1/XI0/XI0_33/d_2_ DECAP_INV_G11
XG13650 XI11_1/XI0/XI0_33/d__1_ XI11_1/XI0/XI0_33/d_1_ DECAP_INV_G11
XG13651 XI11_1/XI0/XI0_33/d__0_ XI11_1/XI0/XI0_33/d_0_ DECAP_INV_G11
XG13652 XI11_1/XI0/XI0_33/d_15_ XI11_1/XI0/XI0_33/d__15_ DECAP_INV_G11
XG13653 XI11_1/XI0/XI0_33/d_14_ XI11_1/XI0/XI0_33/d__14_ DECAP_INV_G11
XG13654 XI11_1/XI0/XI0_33/d_13_ XI11_1/XI0/XI0_33/d__13_ DECAP_INV_G11
XG13655 XI11_1/XI0/XI0_33/d_12_ XI11_1/XI0/XI0_33/d__12_ DECAP_INV_G11
XG13656 XI11_1/XI0/XI0_33/d_11_ XI11_1/XI0/XI0_33/d__11_ DECAP_INV_G11
XG13657 XI11_1/XI0/XI0_33/d_10_ XI11_1/XI0/XI0_33/d__10_ DECAP_INV_G11
XG13658 XI11_1/XI0/XI0_33/d_9_ XI11_1/XI0/XI0_33/d__9_ DECAP_INV_G11
XG13659 XI11_1/XI0/XI0_33/d_8_ XI11_1/XI0/XI0_33/d__8_ DECAP_INV_G11
XG13660 XI11_1/XI0/XI0_33/d_7_ XI11_1/XI0/XI0_33/d__7_ DECAP_INV_G11
XG13661 XI11_1/XI0/XI0_33/d_6_ XI11_1/XI0/XI0_33/d__6_ DECAP_INV_G11
XG13662 XI11_1/XI0/XI0_33/d_5_ XI11_1/XI0/XI0_33/d__5_ DECAP_INV_G11
XG13663 XI11_1/XI0/XI0_33/d_4_ XI11_1/XI0/XI0_33/d__4_ DECAP_INV_G11
XG13664 XI11_1/XI0/XI0_33/d_3_ XI11_1/XI0/XI0_33/d__3_ DECAP_INV_G11
XG13665 XI11_1/XI0/XI0_33/d_2_ XI11_1/XI0/XI0_33/d__2_ DECAP_INV_G11
XG13666 XI11_1/XI0/XI0_33/d_1_ XI11_1/XI0/XI0_33/d__1_ DECAP_INV_G11
XG13667 XI11_1/XI0/XI0_33/d_0_ XI11_1/XI0/XI0_33/d__0_ DECAP_INV_G11
XG13668 XI11_1/XI0/XI0_32/d__15_ XI11_1/XI0/XI0_32/d_15_ DECAP_INV_G11
XG13669 XI11_1/XI0/XI0_32/d__14_ XI11_1/XI0/XI0_32/d_14_ DECAP_INV_G11
XG13670 XI11_1/XI0/XI0_32/d__13_ XI11_1/XI0/XI0_32/d_13_ DECAP_INV_G11
XG13671 XI11_1/XI0/XI0_32/d__12_ XI11_1/XI0/XI0_32/d_12_ DECAP_INV_G11
XG13672 XI11_1/XI0/XI0_32/d__11_ XI11_1/XI0/XI0_32/d_11_ DECAP_INV_G11
XG13673 XI11_1/XI0/XI0_32/d__10_ XI11_1/XI0/XI0_32/d_10_ DECAP_INV_G11
XG13674 XI11_1/XI0/XI0_32/d__9_ XI11_1/XI0/XI0_32/d_9_ DECAP_INV_G11
XG13675 XI11_1/XI0/XI0_32/d__8_ XI11_1/XI0/XI0_32/d_8_ DECAP_INV_G11
XG13676 XI11_1/XI0/XI0_32/d__7_ XI11_1/XI0/XI0_32/d_7_ DECAP_INV_G11
XG13677 XI11_1/XI0/XI0_32/d__6_ XI11_1/XI0/XI0_32/d_6_ DECAP_INV_G11
XG13678 XI11_1/XI0/XI0_32/d__5_ XI11_1/XI0/XI0_32/d_5_ DECAP_INV_G11
XG13679 XI11_1/XI0/XI0_32/d__4_ XI11_1/XI0/XI0_32/d_4_ DECAP_INV_G11
XG13680 XI11_1/XI0/XI0_32/d__3_ XI11_1/XI0/XI0_32/d_3_ DECAP_INV_G11
XG13681 XI11_1/XI0/XI0_32/d__2_ XI11_1/XI0/XI0_32/d_2_ DECAP_INV_G11
XG13682 XI11_1/XI0/XI0_32/d__1_ XI11_1/XI0/XI0_32/d_1_ DECAP_INV_G11
XG13683 XI11_1/XI0/XI0_32/d__0_ XI11_1/XI0/XI0_32/d_0_ DECAP_INV_G11
XG13684 XI11_1/XI0/XI0_32/d_15_ XI11_1/XI0/XI0_32/d__15_ DECAP_INV_G11
XG13685 XI11_1/XI0/XI0_32/d_14_ XI11_1/XI0/XI0_32/d__14_ DECAP_INV_G11
XG13686 XI11_1/XI0/XI0_32/d_13_ XI11_1/XI0/XI0_32/d__13_ DECAP_INV_G11
XG13687 XI11_1/XI0/XI0_32/d_12_ XI11_1/XI0/XI0_32/d__12_ DECAP_INV_G11
XG13688 XI11_1/XI0/XI0_32/d_11_ XI11_1/XI0/XI0_32/d__11_ DECAP_INV_G11
XG13689 XI11_1/XI0/XI0_32/d_10_ XI11_1/XI0/XI0_32/d__10_ DECAP_INV_G11
XG13690 XI11_1/XI0/XI0_32/d_9_ XI11_1/XI0/XI0_32/d__9_ DECAP_INV_G11
XG13691 XI11_1/XI0/XI0_32/d_8_ XI11_1/XI0/XI0_32/d__8_ DECAP_INV_G11
XG13692 XI11_1/XI0/XI0_32/d_7_ XI11_1/XI0/XI0_32/d__7_ DECAP_INV_G11
XG13693 XI11_1/XI0/XI0_32/d_6_ XI11_1/XI0/XI0_32/d__6_ DECAP_INV_G11
XG13694 XI11_1/XI0/XI0_32/d_5_ XI11_1/XI0/XI0_32/d__5_ DECAP_INV_G11
XG13695 XI11_1/XI0/XI0_32/d_4_ XI11_1/XI0/XI0_32/d__4_ DECAP_INV_G11
XG13696 XI11_1/XI0/XI0_32/d_3_ XI11_1/XI0/XI0_32/d__3_ DECAP_INV_G11
XG13697 XI11_1/XI0/XI0_32/d_2_ XI11_1/XI0/XI0_32/d__2_ DECAP_INV_G11
XG13698 XI11_1/XI0/XI0_32/d_1_ XI11_1/XI0/XI0_32/d__1_ DECAP_INV_G11
XG13699 XI11_1/XI0/XI0_32/d_0_ XI11_1/XI0/XI0_32/d__0_ DECAP_INV_G11
XG13700 XI11_1/XI0/XI0_31/d__15_ XI11_1/XI0/XI0_31/d_15_ DECAP_INV_G11
XG13701 XI11_1/XI0/XI0_31/d__14_ XI11_1/XI0/XI0_31/d_14_ DECAP_INV_G11
XG13702 XI11_1/XI0/XI0_31/d__13_ XI11_1/XI0/XI0_31/d_13_ DECAP_INV_G11
XG13703 XI11_1/XI0/XI0_31/d__12_ XI11_1/XI0/XI0_31/d_12_ DECAP_INV_G11
XG13704 XI11_1/XI0/XI0_31/d__11_ XI11_1/XI0/XI0_31/d_11_ DECAP_INV_G11
XG13705 XI11_1/XI0/XI0_31/d__10_ XI11_1/XI0/XI0_31/d_10_ DECAP_INV_G11
XG13706 XI11_1/XI0/XI0_31/d__9_ XI11_1/XI0/XI0_31/d_9_ DECAP_INV_G11
XG13707 XI11_1/XI0/XI0_31/d__8_ XI11_1/XI0/XI0_31/d_8_ DECAP_INV_G11
XG13708 XI11_1/XI0/XI0_31/d__7_ XI11_1/XI0/XI0_31/d_7_ DECAP_INV_G11
XG13709 XI11_1/XI0/XI0_31/d__6_ XI11_1/XI0/XI0_31/d_6_ DECAP_INV_G11
XG13710 XI11_1/XI0/XI0_31/d__5_ XI11_1/XI0/XI0_31/d_5_ DECAP_INV_G11
XG13711 XI11_1/XI0/XI0_31/d__4_ XI11_1/XI0/XI0_31/d_4_ DECAP_INV_G11
XG13712 XI11_1/XI0/XI0_31/d__3_ XI11_1/XI0/XI0_31/d_3_ DECAP_INV_G11
XG13713 XI11_1/XI0/XI0_31/d__2_ XI11_1/XI0/XI0_31/d_2_ DECAP_INV_G11
XG13714 XI11_1/XI0/XI0_31/d__1_ XI11_1/XI0/XI0_31/d_1_ DECAP_INV_G11
XG13715 XI11_1/XI0/XI0_31/d__0_ XI11_1/XI0/XI0_31/d_0_ DECAP_INV_G11
XG13716 XI11_1/XI0/XI0_31/d_15_ XI11_1/XI0/XI0_31/d__15_ DECAP_INV_G11
XG13717 XI11_1/XI0/XI0_31/d_14_ XI11_1/XI0/XI0_31/d__14_ DECAP_INV_G11
XG13718 XI11_1/XI0/XI0_31/d_13_ XI11_1/XI0/XI0_31/d__13_ DECAP_INV_G11
XG13719 XI11_1/XI0/XI0_31/d_12_ XI11_1/XI0/XI0_31/d__12_ DECAP_INV_G11
XG13720 XI11_1/XI0/XI0_31/d_11_ XI11_1/XI0/XI0_31/d__11_ DECAP_INV_G11
XG13721 XI11_1/XI0/XI0_31/d_10_ XI11_1/XI0/XI0_31/d__10_ DECAP_INV_G11
XG13722 XI11_1/XI0/XI0_31/d_9_ XI11_1/XI0/XI0_31/d__9_ DECAP_INV_G11
XG13723 XI11_1/XI0/XI0_31/d_8_ XI11_1/XI0/XI0_31/d__8_ DECAP_INV_G11
XG13724 XI11_1/XI0/XI0_31/d_7_ XI11_1/XI0/XI0_31/d__7_ DECAP_INV_G11
XG13725 XI11_1/XI0/XI0_31/d_6_ XI11_1/XI0/XI0_31/d__6_ DECAP_INV_G11
XG13726 XI11_1/XI0/XI0_31/d_5_ XI11_1/XI0/XI0_31/d__5_ DECAP_INV_G11
XG13727 XI11_1/XI0/XI0_31/d_4_ XI11_1/XI0/XI0_31/d__4_ DECAP_INV_G11
XG13728 XI11_1/XI0/XI0_31/d_3_ XI11_1/XI0/XI0_31/d__3_ DECAP_INV_G11
XG13729 XI11_1/XI0/XI0_31/d_2_ XI11_1/XI0/XI0_31/d__2_ DECAP_INV_G11
XG13730 XI11_1/XI0/XI0_31/d_1_ XI11_1/XI0/XI0_31/d__1_ DECAP_INV_G11
XG13731 XI11_1/XI0/XI0_31/d_0_ XI11_1/XI0/XI0_31/d__0_ DECAP_INV_G11
XG13732 XI11_1/XI0/XI0_30/d__15_ XI11_1/XI0/XI0_30/d_15_ DECAP_INV_G11
XG13733 XI11_1/XI0/XI0_30/d__14_ XI11_1/XI0/XI0_30/d_14_ DECAP_INV_G11
XG13734 XI11_1/XI0/XI0_30/d__13_ XI11_1/XI0/XI0_30/d_13_ DECAP_INV_G11
XG13735 XI11_1/XI0/XI0_30/d__12_ XI11_1/XI0/XI0_30/d_12_ DECAP_INV_G11
XG13736 XI11_1/XI0/XI0_30/d__11_ XI11_1/XI0/XI0_30/d_11_ DECAP_INV_G11
XG13737 XI11_1/XI0/XI0_30/d__10_ XI11_1/XI0/XI0_30/d_10_ DECAP_INV_G11
XG13738 XI11_1/XI0/XI0_30/d__9_ XI11_1/XI0/XI0_30/d_9_ DECAP_INV_G11
XG13739 XI11_1/XI0/XI0_30/d__8_ XI11_1/XI0/XI0_30/d_8_ DECAP_INV_G11
XG13740 XI11_1/XI0/XI0_30/d__7_ XI11_1/XI0/XI0_30/d_7_ DECAP_INV_G11
XG13741 XI11_1/XI0/XI0_30/d__6_ XI11_1/XI0/XI0_30/d_6_ DECAP_INV_G11
XG13742 XI11_1/XI0/XI0_30/d__5_ XI11_1/XI0/XI0_30/d_5_ DECAP_INV_G11
XG13743 XI11_1/XI0/XI0_30/d__4_ XI11_1/XI0/XI0_30/d_4_ DECAP_INV_G11
XG13744 XI11_1/XI0/XI0_30/d__3_ XI11_1/XI0/XI0_30/d_3_ DECAP_INV_G11
XG13745 XI11_1/XI0/XI0_30/d__2_ XI11_1/XI0/XI0_30/d_2_ DECAP_INV_G11
XG13746 XI11_1/XI0/XI0_30/d__1_ XI11_1/XI0/XI0_30/d_1_ DECAP_INV_G11
XG13747 XI11_1/XI0/XI0_30/d__0_ XI11_1/XI0/XI0_30/d_0_ DECAP_INV_G11
XG13748 XI11_1/XI0/XI0_30/d_15_ XI11_1/XI0/XI0_30/d__15_ DECAP_INV_G11
XG13749 XI11_1/XI0/XI0_30/d_14_ XI11_1/XI0/XI0_30/d__14_ DECAP_INV_G11
XG13750 XI11_1/XI0/XI0_30/d_13_ XI11_1/XI0/XI0_30/d__13_ DECAP_INV_G11
XG13751 XI11_1/XI0/XI0_30/d_12_ XI11_1/XI0/XI0_30/d__12_ DECAP_INV_G11
XG13752 XI11_1/XI0/XI0_30/d_11_ XI11_1/XI0/XI0_30/d__11_ DECAP_INV_G11
XG13753 XI11_1/XI0/XI0_30/d_10_ XI11_1/XI0/XI0_30/d__10_ DECAP_INV_G11
XG13754 XI11_1/XI0/XI0_30/d_9_ XI11_1/XI0/XI0_30/d__9_ DECAP_INV_G11
XG13755 XI11_1/XI0/XI0_30/d_8_ XI11_1/XI0/XI0_30/d__8_ DECAP_INV_G11
XG13756 XI11_1/XI0/XI0_30/d_7_ XI11_1/XI0/XI0_30/d__7_ DECAP_INV_G11
XG13757 XI11_1/XI0/XI0_30/d_6_ XI11_1/XI0/XI0_30/d__6_ DECAP_INV_G11
XG13758 XI11_1/XI0/XI0_30/d_5_ XI11_1/XI0/XI0_30/d__5_ DECAP_INV_G11
XG13759 XI11_1/XI0/XI0_30/d_4_ XI11_1/XI0/XI0_30/d__4_ DECAP_INV_G11
XG13760 XI11_1/XI0/XI0_30/d_3_ XI11_1/XI0/XI0_30/d__3_ DECAP_INV_G11
XG13761 XI11_1/XI0/XI0_30/d_2_ XI11_1/XI0/XI0_30/d__2_ DECAP_INV_G11
XG13762 XI11_1/XI0/XI0_30/d_1_ XI11_1/XI0/XI0_30/d__1_ DECAP_INV_G11
XG13763 XI11_1/XI0/XI0_30/d_0_ XI11_1/XI0/XI0_30/d__0_ DECAP_INV_G11
XG13764 XI11_1/XI0/XI0_29/d__15_ XI11_1/XI0/XI0_29/d_15_ DECAP_INV_G11
XG13765 XI11_1/XI0/XI0_29/d__14_ XI11_1/XI0/XI0_29/d_14_ DECAP_INV_G11
XG13766 XI11_1/XI0/XI0_29/d__13_ XI11_1/XI0/XI0_29/d_13_ DECAP_INV_G11
XG13767 XI11_1/XI0/XI0_29/d__12_ XI11_1/XI0/XI0_29/d_12_ DECAP_INV_G11
XG13768 XI11_1/XI0/XI0_29/d__11_ XI11_1/XI0/XI0_29/d_11_ DECAP_INV_G11
XG13769 XI11_1/XI0/XI0_29/d__10_ XI11_1/XI0/XI0_29/d_10_ DECAP_INV_G11
XG13770 XI11_1/XI0/XI0_29/d__9_ XI11_1/XI0/XI0_29/d_9_ DECAP_INV_G11
XG13771 XI11_1/XI0/XI0_29/d__8_ XI11_1/XI0/XI0_29/d_8_ DECAP_INV_G11
XG13772 XI11_1/XI0/XI0_29/d__7_ XI11_1/XI0/XI0_29/d_7_ DECAP_INV_G11
XG13773 XI11_1/XI0/XI0_29/d__6_ XI11_1/XI0/XI0_29/d_6_ DECAP_INV_G11
XG13774 XI11_1/XI0/XI0_29/d__5_ XI11_1/XI0/XI0_29/d_5_ DECAP_INV_G11
XG13775 XI11_1/XI0/XI0_29/d__4_ XI11_1/XI0/XI0_29/d_4_ DECAP_INV_G11
XG13776 XI11_1/XI0/XI0_29/d__3_ XI11_1/XI0/XI0_29/d_3_ DECAP_INV_G11
XG13777 XI11_1/XI0/XI0_29/d__2_ XI11_1/XI0/XI0_29/d_2_ DECAP_INV_G11
XG13778 XI11_1/XI0/XI0_29/d__1_ XI11_1/XI0/XI0_29/d_1_ DECAP_INV_G11
XG13779 XI11_1/XI0/XI0_29/d__0_ XI11_1/XI0/XI0_29/d_0_ DECAP_INV_G11
XG13780 XI11_1/XI0/XI0_29/d_15_ XI11_1/XI0/XI0_29/d__15_ DECAP_INV_G11
XG13781 XI11_1/XI0/XI0_29/d_14_ XI11_1/XI0/XI0_29/d__14_ DECAP_INV_G11
XG13782 XI11_1/XI0/XI0_29/d_13_ XI11_1/XI0/XI0_29/d__13_ DECAP_INV_G11
XG13783 XI11_1/XI0/XI0_29/d_12_ XI11_1/XI0/XI0_29/d__12_ DECAP_INV_G11
XG13784 XI11_1/XI0/XI0_29/d_11_ XI11_1/XI0/XI0_29/d__11_ DECAP_INV_G11
XG13785 XI11_1/XI0/XI0_29/d_10_ XI11_1/XI0/XI0_29/d__10_ DECAP_INV_G11
XG13786 XI11_1/XI0/XI0_29/d_9_ XI11_1/XI0/XI0_29/d__9_ DECAP_INV_G11
XG13787 XI11_1/XI0/XI0_29/d_8_ XI11_1/XI0/XI0_29/d__8_ DECAP_INV_G11
XG13788 XI11_1/XI0/XI0_29/d_7_ XI11_1/XI0/XI0_29/d__7_ DECAP_INV_G11
XG13789 XI11_1/XI0/XI0_29/d_6_ XI11_1/XI0/XI0_29/d__6_ DECAP_INV_G11
XG13790 XI11_1/XI0/XI0_29/d_5_ XI11_1/XI0/XI0_29/d__5_ DECAP_INV_G11
XG13791 XI11_1/XI0/XI0_29/d_4_ XI11_1/XI0/XI0_29/d__4_ DECAP_INV_G11
XG13792 XI11_1/XI0/XI0_29/d_3_ XI11_1/XI0/XI0_29/d__3_ DECAP_INV_G11
XG13793 XI11_1/XI0/XI0_29/d_2_ XI11_1/XI0/XI0_29/d__2_ DECAP_INV_G11
XG13794 XI11_1/XI0/XI0_29/d_1_ XI11_1/XI0/XI0_29/d__1_ DECAP_INV_G11
XG13795 XI11_1/XI0/XI0_29/d_0_ XI11_1/XI0/XI0_29/d__0_ DECAP_INV_G11
XG13796 XI11_1/XI0/XI0_28/d__15_ XI11_1/XI0/XI0_28/d_15_ DECAP_INV_G11
XG13797 XI11_1/XI0/XI0_28/d__14_ XI11_1/XI0/XI0_28/d_14_ DECAP_INV_G11
XG13798 XI11_1/XI0/XI0_28/d__13_ XI11_1/XI0/XI0_28/d_13_ DECAP_INV_G11
XG13799 XI11_1/XI0/XI0_28/d__12_ XI11_1/XI0/XI0_28/d_12_ DECAP_INV_G11
XG13800 XI11_1/XI0/XI0_28/d__11_ XI11_1/XI0/XI0_28/d_11_ DECAP_INV_G11
XG13801 XI11_1/XI0/XI0_28/d__10_ XI11_1/XI0/XI0_28/d_10_ DECAP_INV_G11
XG13802 XI11_1/XI0/XI0_28/d__9_ XI11_1/XI0/XI0_28/d_9_ DECAP_INV_G11
XG13803 XI11_1/XI0/XI0_28/d__8_ XI11_1/XI0/XI0_28/d_8_ DECAP_INV_G11
XG13804 XI11_1/XI0/XI0_28/d__7_ XI11_1/XI0/XI0_28/d_7_ DECAP_INV_G11
XG13805 XI11_1/XI0/XI0_28/d__6_ XI11_1/XI0/XI0_28/d_6_ DECAP_INV_G11
XG13806 XI11_1/XI0/XI0_28/d__5_ XI11_1/XI0/XI0_28/d_5_ DECAP_INV_G11
XG13807 XI11_1/XI0/XI0_28/d__4_ XI11_1/XI0/XI0_28/d_4_ DECAP_INV_G11
XG13808 XI11_1/XI0/XI0_28/d__3_ XI11_1/XI0/XI0_28/d_3_ DECAP_INV_G11
XG13809 XI11_1/XI0/XI0_28/d__2_ XI11_1/XI0/XI0_28/d_2_ DECAP_INV_G11
XG13810 XI11_1/XI0/XI0_28/d__1_ XI11_1/XI0/XI0_28/d_1_ DECAP_INV_G11
XG13811 XI11_1/XI0/XI0_28/d__0_ XI11_1/XI0/XI0_28/d_0_ DECAP_INV_G11
XG13812 XI11_1/XI0/XI0_28/d_15_ XI11_1/XI0/XI0_28/d__15_ DECAP_INV_G11
XG13813 XI11_1/XI0/XI0_28/d_14_ XI11_1/XI0/XI0_28/d__14_ DECAP_INV_G11
XG13814 XI11_1/XI0/XI0_28/d_13_ XI11_1/XI0/XI0_28/d__13_ DECAP_INV_G11
XG13815 XI11_1/XI0/XI0_28/d_12_ XI11_1/XI0/XI0_28/d__12_ DECAP_INV_G11
XG13816 XI11_1/XI0/XI0_28/d_11_ XI11_1/XI0/XI0_28/d__11_ DECAP_INV_G11
XG13817 XI11_1/XI0/XI0_28/d_10_ XI11_1/XI0/XI0_28/d__10_ DECAP_INV_G11
XG13818 XI11_1/XI0/XI0_28/d_9_ XI11_1/XI0/XI0_28/d__9_ DECAP_INV_G11
XG13819 XI11_1/XI0/XI0_28/d_8_ XI11_1/XI0/XI0_28/d__8_ DECAP_INV_G11
XG13820 XI11_1/XI0/XI0_28/d_7_ XI11_1/XI0/XI0_28/d__7_ DECAP_INV_G11
XG13821 XI11_1/XI0/XI0_28/d_6_ XI11_1/XI0/XI0_28/d__6_ DECAP_INV_G11
XG13822 XI11_1/XI0/XI0_28/d_5_ XI11_1/XI0/XI0_28/d__5_ DECAP_INV_G11
XG13823 XI11_1/XI0/XI0_28/d_4_ XI11_1/XI0/XI0_28/d__4_ DECAP_INV_G11
XG13824 XI11_1/XI0/XI0_28/d_3_ XI11_1/XI0/XI0_28/d__3_ DECAP_INV_G11
XG13825 XI11_1/XI0/XI0_28/d_2_ XI11_1/XI0/XI0_28/d__2_ DECAP_INV_G11
XG13826 XI11_1/XI0/XI0_28/d_1_ XI11_1/XI0/XI0_28/d__1_ DECAP_INV_G11
XG13827 XI11_1/XI0/XI0_28/d_0_ XI11_1/XI0/XI0_28/d__0_ DECAP_INV_G11
XG13828 XI11_1/XI0/XI0_27/d__15_ XI11_1/XI0/XI0_27/d_15_ DECAP_INV_G11
XG13829 XI11_1/XI0/XI0_27/d__14_ XI11_1/XI0/XI0_27/d_14_ DECAP_INV_G11
XG13830 XI11_1/XI0/XI0_27/d__13_ XI11_1/XI0/XI0_27/d_13_ DECAP_INV_G11
XG13831 XI11_1/XI0/XI0_27/d__12_ XI11_1/XI0/XI0_27/d_12_ DECAP_INV_G11
XG13832 XI11_1/XI0/XI0_27/d__11_ XI11_1/XI0/XI0_27/d_11_ DECAP_INV_G11
XG13833 XI11_1/XI0/XI0_27/d__10_ XI11_1/XI0/XI0_27/d_10_ DECAP_INV_G11
XG13834 XI11_1/XI0/XI0_27/d__9_ XI11_1/XI0/XI0_27/d_9_ DECAP_INV_G11
XG13835 XI11_1/XI0/XI0_27/d__8_ XI11_1/XI0/XI0_27/d_8_ DECAP_INV_G11
XG13836 XI11_1/XI0/XI0_27/d__7_ XI11_1/XI0/XI0_27/d_7_ DECAP_INV_G11
XG13837 XI11_1/XI0/XI0_27/d__6_ XI11_1/XI0/XI0_27/d_6_ DECAP_INV_G11
XG13838 XI11_1/XI0/XI0_27/d__5_ XI11_1/XI0/XI0_27/d_5_ DECAP_INV_G11
XG13839 XI11_1/XI0/XI0_27/d__4_ XI11_1/XI0/XI0_27/d_4_ DECAP_INV_G11
XG13840 XI11_1/XI0/XI0_27/d__3_ XI11_1/XI0/XI0_27/d_3_ DECAP_INV_G11
XG13841 XI11_1/XI0/XI0_27/d__2_ XI11_1/XI0/XI0_27/d_2_ DECAP_INV_G11
XG13842 XI11_1/XI0/XI0_27/d__1_ XI11_1/XI0/XI0_27/d_1_ DECAP_INV_G11
XG13843 XI11_1/XI0/XI0_27/d__0_ XI11_1/XI0/XI0_27/d_0_ DECAP_INV_G11
XG13844 XI11_1/XI0/XI0_27/d_15_ XI11_1/XI0/XI0_27/d__15_ DECAP_INV_G11
XG13845 XI11_1/XI0/XI0_27/d_14_ XI11_1/XI0/XI0_27/d__14_ DECAP_INV_G11
XG13846 XI11_1/XI0/XI0_27/d_13_ XI11_1/XI0/XI0_27/d__13_ DECAP_INV_G11
XG13847 XI11_1/XI0/XI0_27/d_12_ XI11_1/XI0/XI0_27/d__12_ DECAP_INV_G11
XG13848 XI11_1/XI0/XI0_27/d_11_ XI11_1/XI0/XI0_27/d__11_ DECAP_INV_G11
XG13849 XI11_1/XI0/XI0_27/d_10_ XI11_1/XI0/XI0_27/d__10_ DECAP_INV_G11
XG13850 XI11_1/XI0/XI0_27/d_9_ XI11_1/XI0/XI0_27/d__9_ DECAP_INV_G11
XG13851 XI11_1/XI0/XI0_27/d_8_ XI11_1/XI0/XI0_27/d__8_ DECAP_INV_G11
XG13852 XI11_1/XI0/XI0_27/d_7_ XI11_1/XI0/XI0_27/d__7_ DECAP_INV_G11
XG13853 XI11_1/XI0/XI0_27/d_6_ XI11_1/XI0/XI0_27/d__6_ DECAP_INV_G11
XG13854 XI11_1/XI0/XI0_27/d_5_ XI11_1/XI0/XI0_27/d__5_ DECAP_INV_G11
XG13855 XI11_1/XI0/XI0_27/d_4_ XI11_1/XI0/XI0_27/d__4_ DECAP_INV_G11
XG13856 XI11_1/XI0/XI0_27/d_3_ XI11_1/XI0/XI0_27/d__3_ DECAP_INV_G11
XG13857 XI11_1/XI0/XI0_27/d_2_ XI11_1/XI0/XI0_27/d__2_ DECAP_INV_G11
XG13858 XI11_1/XI0/XI0_27/d_1_ XI11_1/XI0/XI0_27/d__1_ DECAP_INV_G11
XG13859 XI11_1/XI0/XI0_27/d_0_ XI11_1/XI0/XI0_27/d__0_ DECAP_INV_G11
XG13860 XI11_1/XI0/XI0_26/d__15_ XI11_1/XI0/XI0_26/d_15_ DECAP_INV_G11
XG13861 XI11_1/XI0/XI0_26/d__14_ XI11_1/XI0/XI0_26/d_14_ DECAP_INV_G11
XG13862 XI11_1/XI0/XI0_26/d__13_ XI11_1/XI0/XI0_26/d_13_ DECAP_INV_G11
XG13863 XI11_1/XI0/XI0_26/d__12_ XI11_1/XI0/XI0_26/d_12_ DECAP_INV_G11
XG13864 XI11_1/XI0/XI0_26/d__11_ XI11_1/XI0/XI0_26/d_11_ DECAP_INV_G11
XG13865 XI11_1/XI0/XI0_26/d__10_ XI11_1/XI0/XI0_26/d_10_ DECAP_INV_G11
XG13866 XI11_1/XI0/XI0_26/d__9_ XI11_1/XI0/XI0_26/d_9_ DECAP_INV_G11
XG13867 XI11_1/XI0/XI0_26/d__8_ XI11_1/XI0/XI0_26/d_8_ DECAP_INV_G11
XG13868 XI11_1/XI0/XI0_26/d__7_ XI11_1/XI0/XI0_26/d_7_ DECAP_INV_G11
XG13869 XI11_1/XI0/XI0_26/d__6_ XI11_1/XI0/XI0_26/d_6_ DECAP_INV_G11
XG13870 XI11_1/XI0/XI0_26/d__5_ XI11_1/XI0/XI0_26/d_5_ DECAP_INV_G11
XG13871 XI11_1/XI0/XI0_26/d__4_ XI11_1/XI0/XI0_26/d_4_ DECAP_INV_G11
XG13872 XI11_1/XI0/XI0_26/d__3_ XI11_1/XI0/XI0_26/d_3_ DECAP_INV_G11
XG13873 XI11_1/XI0/XI0_26/d__2_ XI11_1/XI0/XI0_26/d_2_ DECAP_INV_G11
XG13874 XI11_1/XI0/XI0_26/d__1_ XI11_1/XI0/XI0_26/d_1_ DECAP_INV_G11
XG13875 XI11_1/XI0/XI0_26/d__0_ XI11_1/XI0/XI0_26/d_0_ DECAP_INV_G11
XG13876 XI11_1/XI0/XI0_26/d_15_ XI11_1/XI0/XI0_26/d__15_ DECAP_INV_G11
XG13877 XI11_1/XI0/XI0_26/d_14_ XI11_1/XI0/XI0_26/d__14_ DECAP_INV_G11
XG13878 XI11_1/XI0/XI0_26/d_13_ XI11_1/XI0/XI0_26/d__13_ DECAP_INV_G11
XG13879 XI11_1/XI0/XI0_26/d_12_ XI11_1/XI0/XI0_26/d__12_ DECAP_INV_G11
XG13880 XI11_1/XI0/XI0_26/d_11_ XI11_1/XI0/XI0_26/d__11_ DECAP_INV_G11
XG13881 XI11_1/XI0/XI0_26/d_10_ XI11_1/XI0/XI0_26/d__10_ DECAP_INV_G11
XG13882 XI11_1/XI0/XI0_26/d_9_ XI11_1/XI0/XI0_26/d__9_ DECAP_INV_G11
XG13883 XI11_1/XI0/XI0_26/d_8_ XI11_1/XI0/XI0_26/d__8_ DECAP_INV_G11
XG13884 XI11_1/XI0/XI0_26/d_7_ XI11_1/XI0/XI0_26/d__7_ DECAP_INV_G11
XG13885 XI11_1/XI0/XI0_26/d_6_ XI11_1/XI0/XI0_26/d__6_ DECAP_INV_G11
XG13886 XI11_1/XI0/XI0_26/d_5_ XI11_1/XI0/XI0_26/d__5_ DECAP_INV_G11
XG13887 XI11_1/XI0/XI0_26/d_4_ XI11_1/XI0/XI0_26/d__4_ DECAP_INV_G11
XG13888 XI11_1/XI0/XI0_26/d_3_ XI11_1/XI0/XI0_26/d__3_ DECAP_INV_G11
XG13889 XI11_1/XI0/XI0_26/d_2_ XI11_1/XI0/XI0_26/d__2_ DECAP_INV_G11
XG13890 XI11_1/XI0/XI0_26/d_1_ XI11_1/XI0/XI0_26/d__1_ DECAP_INV_G11
XG13891 XI11_1/XI0/XI0_26/d_0_ XI11_1/XI0/XI0_26/d__0_ DECAP_INV_G11
XG13892 XI11_1/XI0/XI0_25/d__15_ XI11_1/XI0/XI0_25/d_15_ DECAP_INV_G11
XG13893 XI11_1/XI0/XI0_25/d__14_ XI11_1/XI0/XI0_25/d_14_ DECAP_INV_G11
XG13894 XI11_1/XI0/XI0_25/d__13_ XI11_1/XI0/XI0_25/d_13_ DECAP_INV_G11
XG13895 XI11_1/XI0/XI0_25/d__12_ XI11_1/XI0/XI0_25/d_12_ DECAP_INV_G11
XG13896 XI11_1/XI0/XI0_25/d__11_ XI11_1/XI0/XI0_25/d_11_ DECAP_INV_G11
XG13897 XI11_1/XI0/XI0_25/d__10_ XI11_1/XI0/XI0_25/d_10_ DECAP_INV_G11
XG13898 XI11_1/XI0/XI0_25/d__9_ XI11_1/XI0/XI0_25/d_9_ DECAP_INV_G11
XG13899 XI11_1/XI0/XI0_25/d__8_ XI11_1/XI0/XI0_25/d_8_ DECAP_INV_G11
XG13900 XI11_1/XI0/XI0_25/d__7_ XI11_1/XI0/XI0_25/d_7_ DECAP_INV_G11
XG13901 XI11_1/XI0/XI0_25/d__6_ XI11_1/XI0/XI0_25/d_6_ DECAP_INV_G11
XG13902 XI11_1/XI0/XI0_25/d__5_ XI11_1/XI0/XI0_25/d_5_ DECAP_INV_G11
XG13903 XI11_1/XI0/XI0_25/d__4_ XI11_1/XI0/XI0_25/d_4_ DECAP_INV_G11
XG13904 XI11_1/XI0/XI0_25/d__3_ XI11_1/XI0/XI0_25/d_3_ DECAP_INV_G11
XG13905 XI11_1/XI0/XI0_25/d__2_ XI11_1/XI0/XI0_25/d_2_ DECAP_INV_G11
XG13906 XI11_1/XI0/XI0_25/d__1_ XI11_1/XI0/XI0_25/d_1_ DECAP_INV_G11
XG13907 XI11_1/XI0/XI0_25/d__0_ XI11_1/XI0/XI0_25/d_0_ DECAP_INV_G11
XG13908 XI11_1/XI0/XI0_25/d_15_ XI11_1/XI0/XI0_25/d__15_ DECAP_INV_G11
XG13909 XI11_1/XI0/XI0_25/d_14_ XI11_1/XI0/XI0_25/d__14_ DECAP_INV_G11
XG13910 XI11_1/XI0/XI0_25/d_13_ XI11_1/XI0/XI0_25/d__13_ DECAP_INV_G11
XG13911 XI11_1/XI0/XI0_25/d_12_ XI11_1/XI0/XI0_25/d__12_ DECAP_INV_G11
XG13912 XI11_1/XI0/XI0_25/d_11_ XI11_1/XI0/XI0_25/d__11_ DECAP_INV_G11
XG13913 XI11_1/XI0/XI0_25/d_10_ XI11_1/XI0/XI0_25/d__10_ DECAP_INV_G11
XG13914 XI11_1/XI0/XI0_25/d_9_ XI11_1/XI0/XI0_25/d__9_ DECAP_INV_G11
XG13915 XI11_1/XI0/XI0_25/d_8_ XI11_1/XI0/XI0_25/d__8_ DECAP_INV_G11
XG13916 XI11_1/XI0/XI0_25/d_7_ XI11_1/XI0/XI0_25/d__7_ DECAP_INV_G11
XG13917 XI11_1/XI0/XI0_25/d_6_ XI11_1/XI0/XI0_25/d__6_ DECAP_INV_G11
XG13918 XI11_1/XI0/XI0_25/d_5_ XI11_1/XI0/XI0_25/d__5_ DECAP_INV_G11
XG13919 XI11_1/XI0/XI0_25/d_4_ XI11_1/XI0/XI0_25/d__4_ DECAP_INV_G11
XG13920 XI11_1/XI0/XI0_25/d_3_ XI11_1/XI0/XI0_25/d__3_ DECAP_INV_G11
XG13921 XI11_1/XI0/XI0_25/d_2_ XI11_1/XI0/XI0_25/d__2_ DECAP_INV_G11
XG13922 XI11_1/XI0/XI0_25/d_1_ XI11_1/XI0/XI0_25/d__1_ DECAP_INV_G11
XG13923 XI11_1/XI0/XI0_25/d_0_ XI11_1/XI0/XI0_25/d__0_ DECAP_INV_G11
XG13924 XI11_1/XI0/XI0_24/d__15_ XI11_1/XI0/XI0_24/d_15_ DECAP_INV_G11
XG13925 XI11_1/XI0/XI0_24/d__14_ XI11_1/XI0/XI0_24/d_14_ DECAP_INV_G11
XG13926 XI11_1/XI0/XI0_24/d__13_ XI11_1/XI0/XI0_24/d_13_ DECAP_INV_G11
XG13927 XI11_1/XI0/XI0_24/d__12_ XI11_1/XI0/XI0_24/d_12_ DECAP_INV_G11
XG13928 XI11_1/XI0/XI0_24/d__11_ XI11_1/XI0/XI0_24/d_11_ DECAP_INV_G11
XG13929 XI11_1/XI0/XI0_24/d__10_ XI11_1/XI0/XI0_24/d_10_ DECAP_INV_G11
XG13930 XI11_1/XI0/XI0_24/d__9_ XI11_1/XI0/XI0_24/d_9_ DECAP_INV_G11
XG13931 XI11_1/XI0/XI0_24/d__8_ XI11_1/XI0/XI0_24/d_8_ DECAP_INV_G11
XG13932 XI11_1/XI0/XI0_24/d__7_ XI11_1/XI0/XI0_24/d_7_ DECAP_INV_G11
XG13933 XI11_1/XI0/XI0_24/d__6_ XI11_1/XI0/XI0_24/d_6_ DECAP_INV_G11
XG13934 XI11_1/XI0/XI0_24/d__5_ XI11_1/XI0/XI0_24/d_5_ DECAP_INV_G11
XG13935 XI11_1/XI0/XI0_24/d__4_ XI11_1/XI0/XI0_24/d_4_ DECAP_INV_G11
XG13936 XI11_1/XI0/XI0_24/d__3_ XI11_1/XI0/XI0_24/d_3_ DECAP_INV_G11
XG13937 XI11_1/XI0/XI0_24/d__2_ XI11_1/XI0/XI0_24/d_2_ DECAP_INV_G11
XG13938 XI11_1/XI0/XI0_24/d__1_ XI11_1/XI0/XI0_24/d_1_ DECAP_INV_G11
XG13939 XI11_1/XI0/XI0_24/d__0_ XI11_1/XI0/XI0_24/d_0_ DECAP_INV_G11
XG13940 XI11_1/XI0/XI0_24/d_15_ XI11_1/XI0/XI0_24/d__15_ DECAP_INV_G11
XG13941 XI11_1/XI0/XI0_24/d_14_ XI11_1/XI0/XI0_24/d__14_ DECAP_INV_G11
XG13942 XI11_1/XI0/XI0_24/d_13_ XI11_1/XI0/XI0_24/d__13_ DECAP_INV_G11
XG13943 XI11_1/XI0/XI0_24/d_12_ XI11_1/XI0/XI0_24/d__12_ DECAP_INV_G11
XG13944 XI11_1/XI0/XI0_24/d_11_ XI11_1/XI0/XI0_24/d__11_ DECAP_INV_G11
XG13945 XI11_1/XI0/XI0_24/d_10_ XI11_1/XI0/XI0_24/d__10_ DECAP_INV_G11
XG13946 XI11_1/XI0/XI0_24/d_9_ XI11_1/XI0/XI0_24/d__9_ DECAP_INV_G11
XG13947 XI11_1/XI0/XI0_24/d_8_ XI11_1/XI0/XI0_24/d__8_ DECAP_INV_G11
XG13948 XI11_1/XI0/XI0_24/d_7_ XI11_1/XI0/XI0_24/d__7_ DECAP_INV_G11
XG13949 XI11_1/XI0/XI0_24/d_6_ XI11_1/XI0/XI0_24/d__6_ DECAP_INV_G11
XG13950 XI11_1/XI0/XI0_24/d_5_ XI11_1/XI0/XI0_24/d__5_ DECAP_INV_G11
XG13951 XI11_1/XI0/XI0_24/d_4_ XI11_1/XI0/XI0_24/d__4_ DECAP_INV_G11
XG13952 XI11_1/XI0/XI0_24/d_3_ XI11_1/XI0/XI0_24/d__3_ DECAP_INV_G11
XG13953 XI11_1/XI0/XI0_24/d_2_ XI11_1/XI0/XI0_24/d__2_ DECAP_INV_G11
XG13954 XI11_1/XI0/XI0_24/d_1_ XI11_1/XI0/XI0_24/d__1_ DECAP_INV_G11
XG13955 XI11_1/XI0/XI0_24/d_0_ XI11_1/XI0/XI0_24/d__0_ DECAP_INV_G11
XG13956 XI11_1/XI0/XI0_23/d__15_ XI11_1/XI0/XI0_23/d_15_ DECAP_INV_G11
XG13957 XI11_1/XI0/XI0_23/d__14_ XI11_1/XI0/XI0_23/d_14_ DECAP_INV_G11
XG13958 XI11_1/XI0/XI0_23/d__13_ XI11_1/XI0/XI0_23/d_13_ DECAP_INV_G11
XG13959 XI11_1/XI0/XI0_23/d__12_ XI11_1/XI0/XI0_23/d_12_ DECAP_INV_G11
XG13960 XI11_1/XI0/XI0_23/d__11_ XI11_1/XI0/XI0_23/d_11_ DECAP_INV_G11
XG13961 XI11_1/XI0/XI0_23/d__10_ XI11_1/XI0/XI0_23/d_10_ DECAP_INV_G11
XG13962 XI11_1/XI0/XI0_23/d__9_ XI11_1/XI0/XI0_23/d_9_ DECAP_INV_G11
XG13963 XI11_1/XI0/XI0_23/d__8_ XI11_1/XI0/XI0_23/d_8_ DECAP_INV_G11
XG13964 XI11_1/XI0/XI0_23/d__7_ XI11_1/XI0/XI0_23/d_7_ DECAP_INV_G11
XG13965 XI11_1/XI0/XI0_23/d__6_ XI11_1/XI0/XI0_23/d_6_ DECAP_INV_G11
XG13966 XI11_1/XI0/XI0_23/d__5_ XI11_1/XI0/XI0_23/d_5_ DECAP_INV_G11
XG13967 XI11_1/XI0/XI0_23/d__4_ XI11_1/XI0/XI0_23/d_4_ DECAP_INV_G11
XG13968 XI11_1/XI0/XI0_23/d__3_ XI11_1/XI0/XI0_23/d_3_ DECAP_INV_G11
XG13969 XI11_1/XI0/XI0_23/d__2_ XI11_1/XI0/XI0_23/d_2_ DECAP_INV_G11
XG13970 XI11_1/XI0/XI0_23/d__1_ XI11_1/XI0/XI0_23/d_1_ DECAP_INV_G11
XG13971 XI11_1/XI0/XI0_23/d__0_ XI11_1/XI0/XI0_23/d_0_ DECAP_INV_G11
XG13972 XI11_1/XI0/XI0_23/d_15_ XI11_1/XI0/XI0_23/d__15_ DECAP_INV_G11
XG13973 XI11_1/XI0/XI0_23/d_14_ XI11_1/XI0/XI0_23/d__14_ DECAP_INV_G11
XG13974 XI11_1/XI0/XI0_23/d_13_ XI11_1/XI0/XI0_23/d__13_ DECAP_INV_G11
XG13975 XI11_1/XI0/XI0_23/d_12_ XI11_1/XI0/XI0_23/d__12_ DECAP_INV_G11
XG13976 XI11_1/XI0/XI0_23/d_11_ XI11_1/XI0/XI0_23/d__11_ DECAP_INV_G11
XG13977 XI11_1/XI0/XI0_23/d_10_ XI11_1/XI0/XI0_23/d__10_ DECAP_INV_G11
XG13978 XI11_1/XI0/XI0_23/d_9_ XI11_1/XI0/XI0_23/d__9_ DECAP_INV_G11
XG13979 XI11_1/XI0/XI0_23/d_8_ XI11_1/XI0/XI0_23/d__8_ DECAP_INV_G11
XG13980 XI11_1/XI0/XI0_23/d_7_ XI11_1/XI0/XI0_23/d__7_ DECAP_INV_G11
XG13981 XI11_1/XI0/XI0_23/d_6_ XI11_1/XI0/XI0_23/d__6_ DECAP_INV_G11
XG13982 XI11_1/XI0/XI0_23/d_5_ XI11_1/XI0/XI0_23/d__5_ DECAP_INV_G11
XG13983 XI11_1/XI0/XI0_23/d_4_ XI11_1/XI0/XI0_23/d__4_ DECAP_INV_G11
XG13984 XI11_1/XI0/XI0_23/d_3_ XI11_1/XI0/XI0_23/d__3_ DECAP_INV_G11
XG13985 XI11_1/XI0/XI0_23/d_2_ XI11_1/XI0/XI0_23/d__2_ DECAP_INV_G11
XG13986 XI11_1/XI0/XI0_23/d_1_ XI11_1/XI0/XI0_23/d__1_ DECAP_INV_G11
XG13987 XI11_1/XI0/XI0_23/d_0_ XI11_1/XI0/XI0_23/d__0_ DECAP_INV_G11
XG13988 XI11_1/XI0/XI0_22/d__15_ XI11_1/XI0/XI0_22/d_15_ DECAP_INV_G11
XG13989 XI11_1/XI0/XI0_22/d__14_ XI11_1/XI0/XI0_22/d_14_ DECAP_INV_G11
XG13990 XI11_1/XI0/XI0_22/d__13_ XI11_1/XI0/XI0_22/d_13_ DECAP_INV_G11
XG13991 XI11_1/XI0/XI0_22/d__12_ XI11_1/XI0/XI0_22/d_12_ DECAP_INV_G11
XG13992 XI11_1/XI0/XI0_22/d__11_ XI11_1/XI0/XI0_22/d_11_ DECAP_INV_G11
XG13993 XI11_1/XI0/XI0_22/d__10_ XI11_1/XI0/XI0_22/d_10_ DECAP_INV_G11
XG13994 XI11_1/XI0/XI0_22/d__9_ XI11_1/XI0/XI0_22/d_9_ DECAP_INV_G11
XG13995 XI11_1/XI0/XI0_22/d__8_ XI11_1/XI0/XI0_22/d_8_ DECAP_INV_G11
XG13996 XI11_1/XI0/XI0_22/d__7_ XI11_1/XI0/XI0_22/d_7_ DECAP_INV_G11
XG13997 XI11_1/XI0/XI0_22/d__6_ XI11_1/XI0/XI0_22/d_6_ DECAP_INV_G11
XG13998 XI11_1/XI0/XI0_22/d__5_ XI11_1/XI0/XI0_22/d_5_ DECAP_INV_G11
XG13999 XI11_1/XI0/XI0_22/d__4_ XI11_1/XI0/XI0_22/d_4_ DECAP_INV_G11
XG14000 XI11_1/XI0/XI0_22/d__3_ XI11_1/XI0/XI0_22/d_3_ DECAP_INV_G11
XG14001 XI11_1/XI0/XI0_22/d__2_ XI11_1/XI0/XI0_22/d_2_ DECAP_INV_G11
XG14002 XI11_1/XI0/XI0_22/d__1_ XI11_1/XI0/XI0_22/d_1_ DECAP_INV_G11
XG14003 XI11_1/XI0/XI0_22/d__0_ XI11_1/XI0/XI0_22/d_0_ DECAP_INV_G11
XG14004 XI11_1/XI0/XI0_22/d_15_ XI11_1/XI0/XI0_22/d__15_ DECAP_INV_G11
XG14005 XI11_1/XI0/XI0_22/d_14_ XI11_1/XI0/XI0_22/d__14_ DECAP_INV_G11
XG14006 XI11_1/XI0/XI0_22/d_13_ XI11_1/XI0/XI0_22/d__13_ DECAP_INV_G11
XG14007 XI11_1/XI0/XI0_22/d_12_ XI11_1/XI0/XI0_22/d__12_ DECAP_INV_G11
XG14008 XI11_1/XI0/XI0_22/d_11_ XI11_1/XI0/XI0_22/d__11_ DECAP_INV_G11
XG14009 XI11_1/XI0/XI0_22/d_10_ XI11_1/XI0/XI0_22/d__10_ DECAP_INV_G11
XG14010 XI11_1/XI0/XI0_22/d_9_ XI11_1/XI0/XI0_22/d__9_ DECAP_INV_G11
XG14011 XI11_1/XI0/XI0_22/d_8_ XI11_1/XI0/XI0_22/d__8_ DECAP_INV_G11
XG14012 XI11_1/XI0/XI0_22/d_7_ XI11_1/XI0/XI0_22/d__7_ DECAP_INV_G11
XG14013 XI11_1/XI0/XI0_22/d_6_ XI11_1/XI0/XI0_22/d__6_ DECAP_INV_G11
XG14014 XI11_1/XI0/XI0_22/d_5_ XI11_1/XI0/XI0_22/d__5_ DECAP_INV_G11
XG14015 XI11_1/XI0/XI0_22/d_4_ XI11_1/XI0/XI0_22/d__4_ DECAP_INV_G11
XG14016 XI11_1/XI0/XI0_22/d_3_ XI11_1/XI0/XI0_22/d__3_ DECAP_INV_G11
XG14017 XI11_1/XI0/XI0_22/d_2_ XI11_1/XI0/XI0_22/d__2_ DECAP_INV_G11
XG14018 XI11_1/XI0/XI0_22/d_1_ XI11_1/XI0/XI0_22/d__1_ DECAP_INV_G11
XG14019 XI11_1/XI0/XI0_22/d_0_ XI11_1/XI0/XI0_22/d__0_ DECAP_INV_G11
XG14020 XI11_1/XI0/XI0_21/d__15_ XI11_1/XI0/XI0_21/d_15_ DECAP_INV_G11
XG14021 XI11_1/XI0/XI0_21/d__14_ XI11_1/XI0/XI0_21/d_14_ DECAP_INV_G11
XG14022 XI11_1/XI0/XI0_21/d__13_ XI11_1/XI0/XI0_21/d_13_ DECAP_INV_G11
XG14023 XI11_1/XI0/XI0_21/d__12_ XI11_1/XI0/XI0_21/d_12_ DECAP_INV_G11
XG14024 XI11_1/XI0/XI0_21/d__11_ XI11_1/XI0/XI0_21/d_11_ DECAP_INV_G11
XG14025 XI11_1/XI0/XI0_21/d__10_ XI11_1/XI0/XI0_21/d_10_ DECAP_INV_G11
XG14026 XI11_1/XI0/XI0_21/d__9_ XI11_1/XI0/XI0_21/d_9_ DECAP_INV_G11
XG14027 XI11_1/XI0/XI0_21/d__8_ XI11_1/XI0/XI0_21/d_8_ DECAP_INV_G11
XG14028 XI11_1/XI0/XI0_21/d__7_ XI11_1/XI0/XI0_21/d_7_ DECAP_INV_G11
XG14029 XI11_1/XI0/XI0_21/d__6_ XI11_1/XI0/XI0_21/d_6_ DECAP_INV_G11
XG14030 XI11_1/XI0/XI0_21/d__5_ XI11_1/XI0/XI0_21/d_5_ DECAP_INV_G11
XG14031 XI11_1/XI0/XI0_21/d__4_ XI11_1/XI0/XI0_21/d_4_ DECAP_INV_G11
XG14032 XI11_1/XI0/XI0_21/d__3_ XI11_1/XI0/XI0_21/d_3_ DECAP_INV_G11
XG14033 XI11_1/XI0/XI0_21/d__2_ XI11_1/XI0/XI0_21/d_2_ DECAP_INV_G11
XG14034 XI11_1/XI0/XI0_21/d__1_ XI11_1/XI0/XI0_21/d_1_ DECAP_INV_G11
XG14035 XI11_1/XI0/XI0_21/d__0_ XI11_1/XI0/XI0_21/d_0_ DECAP_INV_G11
XG14036 XI11_1/XI0/XI0_21/d_15_ XI11_1/XI0/XI0_21/d__15_ DECAP_INV_G11
XG14037 XI11_1/XI0/XI0_21/d_14_ XI11_1/XI0/XI0_21/d__14_ DECAP_INV_G11
XG14038 XI11_1/XI0/XI0_21/d_13_ XI11_1/XI0/XI0_21/d__13_ DECAP_INV_G11
XG14039 XI11_1/XI0/XI0_21/d_12_ XI11_1/XI0/XI0_21/d__12_ DECAP_INV_G11
XG14040 XI11_1/XI0/XI0_21/d_11_ XI11_1/XI0/XI0_21/d__11_ DECAP_INV_G11
XG14041 XI11_1/XI0/XI0_21/d_10_ XI11_1/XI0/XI0_21/d__10_ DECAP_INV_G11
XG14042 XI11_1/XI0/XI0_21/d_9_ XI11_1/XI0/XI0_21/d__9_ DECAP_INV_G11
XG14043 XI11_1/XI0/XI0_21/d_8_ XI11_1/XI0/XI0_21/d__8_ DECAP_INV_G11
XG14044 XI11_1/XI0/XI0_21/d_7_ XI11_1/XI0/XI0_21/d__7_ DECAP_INV_G11
XG14045 XI11_1/XI0/XI0_21/d_6_ XI11_1/XI0/XI0_21/d__6_ DECAP_INV_G11
XG14046 XI11_1/XI0/XI0_21/d_5_ XI11_1/XI0/XI0_21/d__5_ DECAP_INV_G11
XG14047 XI11_1/XI0/XI0_21/d_4_ XI11_1/XI0/XI0_21/d__4_ DECAP_INV_G11
XG14048 XI11_1/XI0/XI0_21/d_3_ XI11_1/XI0/XI0_21/d__3_ DECAP_INV_G11
XG14049 XI11_1/XI0/XI0_21/d_2_ XI11_1/XI0/XI0_21/d__2_ DECAP_INV_G11
XG14050 XI11_1/XI0/XI0_21/d_1_ XI11_1/XI0/XI0_21/d__1_ DECAP_INV_G11
XG14051 XI11_1/XI0/XI0_21/d_0_ XI11_1/XI0/XI0_21/d__0_ DECAP_INV_G11
XG14052 XI11_1/XI0/XI0_20/d__15_ XI11_1/XI0/XI0_20/d_15_ DECAP_INV_G11
XG14053 XI11_1/XI0/XI0_20/d__14_ XI11_1/XI0/XI0_20/d_14_ DECAP_INV_G11
XG14054 XI11_1/XI0/XI0_20/d__13_ XI11_1/XI0/XI0_20/d_13_ DECAP_INV_G11
XG14055 XI11_1/XI0/XI0_20/d__12_ XI11_1/XI0/XI0_20/d_12_ DECAP_INV_G11
XG14056 XI11_1/XI0/XI0_20/d__11_ XI11_1/XI0/XI0_20/d_11_ DECAP_INV_G11
XG14057 XI11_1/XI0/XI0_20/d__10_ XI11_1/XI0/XI0_20/d_10_ DECAP_INV_G11
XG14058 XI11_1/XI0/XI0_20/d__9_ XI11_1/XI0/XI0_20/d_9_ DECAP_INV_G11
XG14059 XI11_1/XI0/XI0_20/d__8_ XI11_1/XI0/XI0_20/d_8_ DECAP_INV_G11
XG14060 XI11_1/XI0/XI0_20/d__7_ XI11_1/XI0/XI0_20/d_7_ DECAP_INV_G11
XG14061 XI11_1/XI0/XI0_20/d__6_ XI11_1/XI0/XI0_20/d_6_ DECAP_INV_G11
XG14062 XI11_1/XI0/XI0_20/d__5_ XI11_1/XI0/XI0_20/d_5_ DECAP_INV_G11
XG14063 XI11_1/XI0/XI0_20/d__4_ XI11_1/XI0/XI0_20/d_4_ DECAP_INV_G11
XG14064 XI11_1/XI0/XI0_20/d__3_ XI11_1/XI0/XI0_20/d_3_ DECAP_INV_G11
XG14065 XI11_1/XI0/XI0_20/d__2_ XI11_1/XI0/XI0_20/d_2_ DECAP_INV_G11
XG14066 XI11_1/XI0/XI0_20/d__1_ XI11_1/XI0/XI0_20/d_1_ DECAP_INV_G11
XG14067 XI11_1/XI0/XI0_20/d__0_ XI11_1/XI0/XI0_20/d_0_ DECAP_INV_G11
XG14068 XI11_1/XI0/XI0_20/d_15_ XI11_1/XI0/XI0_20/d__15_ DECAP_INV_G11
XG14069 XI11_1/XI0/XI0_20/d_14_ XI11_1/XI0/XI0_20/d__14_ DECAP_INV_G11
XG14070 XI11_1/XI0/XI0_20/d_13_ XI11_1/XI0/XI0_20/d__13_ DECAP_INV_G11
XG14071 XI11_1/XI0/XI0_20/d_12_ XI11_1/XI0/XI0_20/d__12_ DECAP_INV_G11
XG14072 XI11_1/XI0/XI0_20/d_11_ XI11_1/XI0/XI0_20/d__11_ DECAP_INV_G11
XG14073 XI11_1/XI0/XI0_20/d_10_ XI11_1/XI0/XI0_20/d__10_ DECAP_INV_G11
XG14074 XI11_1/XI0/XI0_20/d_9_ XI11_1/XI0/XI0_20/d__9_ DECAP_INV_G11
XG14075 XI11_1/XI0/XI0_20/d_8_ XI11_1/XI0/XI0_20/d__8_ DECAP_INV_G11
XG14076 XI11_1/XI0/XI0_20/d_7_ XI11_1/XI0/XI0_20/d__7_ DECAP_INV_G11
XG14077 XI11_1/XI0/XI0_20/d_6_ XI11_1/XI0/XI0_20/d__6_ DECAP_INV_G11
XG14078 XI11_1/XI0/XI0_20/d_5_ XI11_1/XI0/XI0_20/d__5_ DECAP_INV_G11
XG14079 XI11_1/XI0/XI0_20/d_4_ XI11_1/XI0/XI0_20/d__4_ DECAP_INV_G11
XG14080 XI11_1/XI0/XI0_20/d_3_ XI11_1/XI0/XI0_20/d__3_ DECAP_INV_G11
XG14081 XI11_1/XI0/XI0_20/d_2_ XI11_1/XI0/XI0_20/d__2_ DECAP_INV_G11
XG14082 XI11_1/XI0/XI0_20/d_1_ XI11_1/XI0/XI0_20/d__1_ DECAP_INV_G11
XG14083 XI11_1/XI0/XI0_20/d_0_ XI11_1/XI0/XI0_20/d__0_ DECAP_INV_G11
XG14084 XI11_1/XI0/XI0_19/d__15_ XI11_1/XI0/XI0_19/d_15_ DECAP_INV_G11
XG14085 XI11_1/XI0/XI0_19/d__14_ XI11_1/XI0/XI0_19/d_14_ DECAP_INV_G11
XG14086 XI11_1/XI0/XI0_19/d__13_ XI11_1/XI0/XI0_19/d_13_ DECAP_INV_G11
XG14087 XI11_1/XI0/XI0_19/d__12_ XI11_1/XI0/XI0_19/d_12_ DECAP_INV_G11
XG14088 XI11_1/XI0/XI0_19/d__11_ XI11_1/XI0/XI0_19/d_11_ DECAP_INV_G11
XG14089 XI11_1/XI0/XI0_19/d__10_ XI11_1/XI0/XI0_19/d_10_ DECAP_INV_G11
XG14090 XI11_1/XI0/XI0_19/d__9_ XI11_1/XI0/XI0_19/d_9_ DECAP_INV_G11
XG14091 XI11_1/XI0/XI0_19/d__8_ XI11_1/XI0/XI0_19/d_8_ DECAP_INV_G11
XG14092 XI11_1/XI0/XI0_19/d__7_ XI11_1/XI0/XI0_19/d_7_ DECAP_INV_G11
XG14093 XI11_1/XI0/XI0_19/d__6_ XI11_1/XI0/XI0_19/d_6_ DECAP_INV_G11
XG14094 XI11_1/XI0/XI0_19/d__5_ XI11_1/XI0/XI0_19/d_5_ DECAP_INV_G11
XG14095 XI11_1/XI0/XI0_19/d__4_ XI11_1/XI0/XI0_19/d_4_ DECAP_INV_G11
XG14096 XI11_1/XI0/XI0_19/d__3_ XI11_1/XI0/XI0_19/d_3_ DECAP_INV_G11
XG14097 XI11_1/XI0/XI0_19/d__2_ XI11_1/XI0/XI0_19/d_2_ DECAP_INV_G11
XG14098 XI11_1/XI0/XI0_19/d__1_ XI11_1/XI0/XI0_19/d_1_ DECAP_INV_G11
XG14099 XI11_1/XI0/XI0_19/d__0_ XI11_1/XI0/XI0_19/d_0_ DECAP_INV_G11
XG14100 XI11_1/XI0/XI0_19/d_15_ XI11_1/XI0/XI0_19/d__15_ DECAP_INV_G11
XG14101 XI11_1/XI0/XI0_19/d_14_ XI11_1/XI0/XI0_19/d__14_ DECAP_INV_G11
XG14102 XI11_1/XI0/XI0_19/d_13_ XI11_1/XI0/XI0_19/d__13_ DECAP_INV_G11
XG14103 XI11_1/XI0/XI0_19/d_12_ XI11_1/XI0/XI0_19/d__12_ DECAP_INV_G11
XG14104 XI11_1/XI0/XI0_19/d_11_ XI11_1/XI0/XI0_19/d__11_ DECAP_INV_G11
XG14105 XI11_1/XI0/XI0_19/d_10_ XI11_1/XI0/XI0_19/d__10_ DECAP_INV_G11
XG14106 XI11_1/XI0/XI0_19/d_9_ XI11_1/XI0/XI0_19/d__9_ DECAP_INV_G11
XG14107 XI11_1/XI0/XI0_19/d_8_ XI11_1/XI0/XI0_19/d__8_ DECAP_INV_G11
XG14108 XI11_1/XI0/XI0_19/d_7_ XI11_1/XI0/XI0_19/d__7_ DECAP_INV_G11
XG14109 XI11_1/XI0/XI0_19/d_6_ XI11_1/XI0/XI0_19/d__6_ DECAP_INV_G11
XG14110 XI11_1/XI0/XI0_19/d_5_ XI11_1/XI0/XI0_19/d__5_ DECAP_INV_G11
XG14111 XI11_1/XI0/XI0_19/d_4_ XI11_1/XI0/XI0_19/d__4_ DECAP_INV_G11
XG14112 XI11_1/XI0/XI0_19/d_3_ XI11_1/XI0/XI0_19/d__3_ DECAP_INV_G11
XG14113 XI11_1/XI0/XI0_19/d_2_ XI11_1/XI0/XI0_19/d__2_ DECAP_INV_G11
XG14114 XI11_1/XI0/XI0_19/d_1_ XI11_1/XI0/XI0_19/d__1_ DECAP_INV_G11
XG14115 XI11_1/XI0/XI0_19/d_0_ XI11_1/XI0/XI0_19/d__0_ DECAP_INV_G11
XG14116 XI11_1/XI0/XI0_18/d__15_ XI11_1/XI0/XI0_18/d_15_ DECAP_INV_G11
XG14117 XI11_1/XI0/XI0_18/d__14_ XI11_1/XI0/XI0_18/d_14_ DECAP_INV_G11
XG14118 XI11_1/XI0/XI0_18/d__13_ XI11_1/XI0/XI0_18/d_13_ DECAP_INV_G11
XG14119 XI11_1/XI0/XI0_18/d__12_ XI11_1/XI0/XI0_18/d_12_ DECAP_INV_G11
XG14120 XI11_1/XI0/XI0_18/d__11_ XI11_1/XI0/XI0_18/d_11_ DECAP_INV_G11
XG14121 XI11_1/XI0/XI0_18/d__10_ XI11_1/XI0/XI0_18/d_10_ DECAP_INV_G11
XG14122 XI11_1/XI0/XI0_18/d__9_ XI11_1/XI0/XI0_18/d_9_ DECAP_INV_G11
XG14123 XI11_1/XI0/XI0_18/d__8_ XI11_1/XI0/XI0_18/d_8_ DECAP_INV_G11
XG14124 XI11_1/XI0/XI0_18/d__7_ XI11_1/XI0/XI0_18/d_7_ DECAP_INV_G11
XG14125 XI11_1/XI0/XI0_18/d__6_ XI11_1/XI0/XI0_18/d_6_ DECAP_INV_G11
XG14126 XI11_1/XI0/XI0_18/d__5_ XI11_1/XI0/XI0_18/d_5_ DECAP_INV_G11
XG14127 XI11_1/XI0/XI0_18/d__4_ XI11_1/XI0/XI0_18/d_4_ DECAP_INV_G11
XG14128 XI11_1/XI0/XI0_18/d__3_ XI11_1/XI0/XI0_18/d_3_ DECAP_INV_G11
XG14129 XI11_1/XI0/XI0_18/d__2_ XI11_1/XI0/XI0_18/d_2_ DECAP_INV_G11
XG14130 XI11_1/XI0/XI0_18/d__1_ XI11_1/XI0/XI0_18/d_1_ DECAP_INV_G11
XG14131 XI11_1/XI0/XI0_18/d__0_ XI11_1/XI0/XI0_18/d_0_ DECAP_INV_G11
XG14132 XI11_1/XI0/XI0_18/d_15_ XI11_1/XI0/XI0_18/d__15_ DECAP_INV_G11
XG14133 XI11_1/XI0/XI0_18/d_14_ XI11_1/XI0/XI0_18/d__14_ DECAP_INV_G11
XG14134 XI11_1/XI0/XI0_18/d_13_ XI11_1/XI0/XI0_18/d__13_ DECAP_INV_G11
XG14135 XI11_1/XI0/XI0_18/d_12_ XI11_1/XI0/XI0_18/d__12_ DECAP_INV_G11
XG14136 XI11_1/XI0/XI0_18/d_11_ XI11_1/XI0/XI0_18/d__11_ DECAP_INV_G11
XG14137 XI11_1/XI0/XI0_18/d_10_ XI11_1/XI0/XI0_18/d__10_ DECAP_INV_G11
XG14138 XI11_1/XI0/XI0_18/d_9_ XI11_1/XI0/XI0_18/d__9_ DECAP_INV_G11
XG14139 XI11_1/XI0/XI0_18/d_8_ XI11_1/XI0/XI0_18/d__8_ DECAP_INV_G11
XG14140 XI11_1/XI0/XI0_18/d_7_ XI11_1/XI0/XI0_18/d__7_ DECAP_INV_G11
XG14141 XI11_1/XI0/XI0_18/d_6_ XI11_1/XI0/XI0_18/d__6_ DECAP_INV_G11
XG14142 XI11_1/XI0/XI0_18/d_5_ XI11_1/XI0/XI0_18/d__5_ DECAP_INV_G11
XG14143 XI11_1/XI0/XI0_18/d_4_ XI11_1/XI0/XI0_18/d__4_ DECAP_INV_G11
XG14144 XI11_1/XI0/XI0_18/d_3_ XI11_1/XI0/XI0_18/d__3_ DECAP_INV_G11
XG14145 XI11_1/XI0/XI0_18/d_2_ XI11_1/XI0/XI0_18/d__2_ DECAP_INV_G11
XG14146 XI11_1/XI0/XI0_18/d_1_ XI11_1/XI0/XI0_18/d__1_ DECAP_INV_G11
XG14147 XI11_1/XI0/XI0_18/d_0_ XI11_1/XI0/XI0_18/d__0_ DECAP_INV_G11
XG14148 XI11_1/XI0/XI0_17/d__15_ XI11_1/XI0/XI0_17/d_15_ DECAP_INV_G11
XG14149 XI11_1/XI0/XI0_17/d__14_ XI11_1/XI0/XI0_17/d_14_ DECAP_INV_G11
XG14150 XI11_1/XI0/XI0_17/d__13_ XI11_1/XI0/XI0_17/d_13_ DECAP_INV_G11
XG14151 XI11_1/XI0/XI0_17/d__12_ XI11_1/XI0/XI0_17/d_12_ DECAP_INV_G11
XG14152 XI11_1/XI0/XI0_17/d__11_ XI11_1/XI0/XI0_17/d_11_ DECAP_INV_G11
XG14153 XI11_1/XI0/XI0_17/d__10_ XI11_1/XI0/XI0_17/d_10_ DECAP_INV_G11
XG14154 XI11_1/XI0/XI0_17/d__9_ XI11_1/XI0/XI0_17/d_9_ DECAP_INV_G11
XG14155 XI11_1/XI0/XI0_17/d__8_ XI11_1/XI0/XI0_17/d_8_ DECAP_INV_G11
XG14156 XI11_1/XI0/XI0_17/d__7_ XI11_1/XI0/XI0_17/d_7_ DECAP_INV_G11
XG14157 XI11_1/XI0/XI0_17/d__6_ XI11_1/XI0/XI0_17/d_6_ DECAP_INV_G11
XG14158 XI11_1/XI0/XI0_17/d__5_ XI11_1/XI0/XI0_17/d_5_ DECAP_INV_G11
XG14159 XI11_1/XI0/XI0_17/d__4_ XI11_1/XI0/XI0_17/d_4_ DECAP_INV_G11
XG14160 XI11_1/XI0/XI0_17/d__3_ XI11_1/XI0/XI0_17/d_3_ DECAP_INV_G11
XG14161 XI11_1/XI0/XI0_17/d__2_ XI11_1/XI0/XI0_17/d_2_ DECAP_INV_G11
XG14162 XI11_1/XI0/XI0_17/d__1_ XI11_1/XI0/XI0_17/d_1_ DECAP_INV_G11
XG14163 XI11_1/XI0/XI0_17/d__0_ XI11_1/XI0/XI0_17/d_0_ DECAP_INV_G11
XG14164 XI11_1/XI0/XI0_17/d_15_ XI11_1/XI0/XI0_17/d__15_ DECAP_INV_G11
XG14165 XI11_1/XI0/XI0_17/d_14_ XI11_1/XI0/XI0_17/d__14_ DECAP_INV_G11
XG14166 XI11_1/XI0/XI0_17/d_13_ XI11_1/XI0/XI0_17/d__13_ DECAP_INV_G11
XG14167 XI11_1/XI0/XI0_17/d_12_ XI11_1/XI0/XI0_17/d__12_ DECAP_INV_G11
XG14168 XI11_1/XI0/XI0_17/d_11_ XI11_1/XI0/XI0_17/d__11_ DECAP_INV_G11
XG14169 XI11_1/XI0/XI0_17/d_10_ XI11_1/XI0/XI0_17/d__10_ DECAP_INV_G11
XG14170 XI11_1/XI0/XI0_17/d_9_ XI11_1/XI0/XI0_17/d__9_ DECAP_INV_G11
XG14171 XI11_1/XI0/XI0_17/d_8_ XI11_1/XI0/XI0_17/d__8_ DECAP_INV_G11
XG14172 XI11_1/XI0/XI0_17/d_7_ XI11_1/XI0/XI0_17/d__7_ DECAP_INV_G11
XG14173 XI11_1/XI0/XI0_17/d_6_ XI11_1/XI0/XI0_17/d__6_ DECAP_INV_G11
XG14174 XI11_1/XI0/XI0_17/d_5_ XI11_1/XI0/XI0_17/d__5_ DECAP_INV_G11
XG14175 XI11_1/XI0/XI0_17/d_4_ XI11_1/XI0/XI0_17/d__4_ DECAP_INV_G11
XG14176 XI11_1/XI0/XI0_17/d_3_ XI11_1/XI0/XI0_17/d__3_ DECAP_INV_G11
XG14177 XI11_1/XI0/XI0_17/d_2_ XI11_1/XI0/XI0_17/d__2_ DECAP_INV_G11
XG14178 XI11_1/XI0/XI0_17/d_1_ XI11_1/XI0/XI0_17/d__1_ DECAP_INV_G11
XG14179 XI11_1/XI0/XI0_17/d_0_ XI11_1/XI0/XI0_17/d__0_ DECAP_INV_G11
XG14180 XI11_1/XI0/XI0_16/d__15_ XI11_1/XI0/XI0_16/d_15_ DECAP_INV_G11
XG14181 XI11_1/XI0/XI0_16/d__14_ XI11_1/XI0/XI0_16/d_14_ DECAP_INV_G11
XG14182 XI11_1/XI0/XI0_16/d__13_ XI11_1/XI0/XI0_16/d_13_ DECAP_INV_G11
XG14183 XI11_1/XI0/XI0_16/d__12_ XI11_1/XI0/XI0_16/d_12_ DECAP_INV_G11
XG14184 XI11_1/XI0/XI0_16/d__11_ XI11_1/XI0/XI0_16/d_11_ DECAP_INV_G11
XG14185 XI11_1/XI0/XI0_16/d__10_ XI11_1/XI0/XI0_16/d_10_ DECAP_INV_G11
XG14186 XI11_1/XI0/XI0_16/d__9_ XI11_1/XI0/XI0_16/d_9_ DECAP_INV_G11
XG14187 XI11_1/XI0/XI0_16/d__8_ XI11_1/XI0/XI0_16/d_8_ DECAP_INV_G11
XG14188 XI11_1/XI0/XI0_16/d__7_ XI11_1/XI0/XI0_16/d_7_ DECAP_INV_G11
XG14189 XI11_1/XI0/XI0_16/d__6_ XI11_1/XI0/XI0_16/d_6_ DECAP_INV_G11
XG14190 XI11_1/XI0/XI0_16/d__5_ XI11_1/XI0/XI0_16/d_5_ DECAP_INV_G11
XG14191 XI11_1/XI0/XI0_16/d__4_ XI11_1/XI0/XI0_16/d_4_ DECAP_INV_G11
XG14192 XI11_1/XI0/XI0_16/d__3_ XI11_1/XI0/XI0_16/d_3_ DECAP_INV_G11
XG14193 XI11_1/XI0/XI0_16/d__2_ XI11_1/XI0/XI0_16/d_2_ DECAP_INV_G11
XG14194 XI11_1/XI0/XI0_16/d__1_ XI11_1/XI0/XI0_16/d_1_ DECAP_INV_G11
XG14195 XI11_1/XI0/XI0_16/d__0_ XI11_1/XI0/XI0_16/d_0_ DECAP_INV_G11
XG14196 XI11_1/XI0/XI0_16/d_15_ XI11_1/XI0/XI0_16/d__15_ DECAP_INV_G11
XG14197 XI11_1/XI0/XI0_16/d_14_ XI11_1/XI0/XI0_16/d__14_ DECAP_INV_G11
XG14198 XI11_1/XI0/XI0_16/d_13_ XI11_1/XI0/XI0_16/d__13_ DECAP_INV_G11
XG14199 XI11_1/XI0/XI0_16/d_12_ XI11_1/XI0/XI0_16/d__12_ DECAP_INV_G11
XG14200 XI11_1/XI0/XI0_16/d_11_ XI11_1/XI0/XI0_16/d__11_ DECAP_INV_G11
XG14201 XI11_1/XI0/XI0_16/d_10_ XI11_1/XI0/XI0_16/d__10_ DECAP_INV_G11
XG14202 XI11_1/XI0/XI0_16/d_9_ XI11_1/XI0/XI0_16/d__9_ DECAP_INV_G11
XG14203 XI11_1/XI0/XI0_16/d_8_ XI11_1/XI0/XI0_16/d__8_ DECAP_INV_G11
XG14204 XI11_1/XI0/XI0_16/d_7_ XI11_1/XI0/XI0_16/d__7_ DECAP_INV_G11
XG14205 XI11_1/XI0/XI0_16/d_6_ XI11_1/XI0/XI0_16/d__6_ DECAP_INV_G11
XG14206 XI11_1/XI0/XI0_16/d_5_ XI11_1/XI0/XI0_16/d__5_ DECAP_INV_G11
XG14207 XI11_1/XI0/XI0_16/d_4_ XI11_1/XI0/XI0_16/d__4_ DECAP_INV_G11
XG14208 XI11_1/XI0/XI0_16/d_3_ XI11_1/XI0/XI0_16/d__3_ DECAP_INV_G11
XG14209 XI11_1/XI0/XI0_16/d_2_ XI11_1/XI0/XI0_16/d__2_ DECAP_INV_G11
XG14210 XI11_1/XI0/XI0_16/d_1_ XI11_1/XI0/XI0_16/d__1_ DECAP_INV_G11
XG14211 XI11_1/XI0/XI0_16/d_0_ XI11_1/XI0/XI0_16/d__0_ DECAP_INV_G11
XG14212 XI11_1/XI0/XI0_15/d__15_ XI11_1/XI0/XI0_15/d_15_ DECAP_INV_G11
XG14213 XI11_1/XI0/XI0_15/d__14_ XI11_1/XI0/XI0_15/d_14_ DECAP_INV_G11
XG14214 XI11_1/XI0/XI0_15/d__13_ XI11_1/XI0/XI0_15/d_13_ DECAP_INV_G11
XG14215 XI11_1/XI0/XI0_15/d__12_ XI11_1/XI0/XI0_15/d_12_ DECAP_INV_G11
XG14216 XI11_1/XI0/XI0_15/d__11_ XI11_1/XI0/XI0_15/d_11_ DECAP_INV_G11
XG14217 XI11_1/XI0/XI0_15/d__10_ XI11_1/XI0/XI0_15/d_10_ DECAP_INV_G11
XG14218 XI11_1/XI0/XI0_15/d__9_ XI11_1/XI0/XI0_15/d_9_ DECAP_INV_G11
XG14219 XI11_1/XI0/XI0_15/d__8_ XI11_1/XI0/XI0_15/d_8_ DECAP_INV_G11
XG14220 XI11_1/XI0/XI0_15/d__7_ XI11_1/XI0/XI0_15/d_7_ DECAP_INV_G11
XG14221 XI11_1/XI0/XI0_15/d__6_ XI11_1/XI0/XI0_15/d_6_ DECAP_INV_G11
XG14222 XI11_1/XI0/XI0_15/d__5_ XI11_1/XI0/XI0_15/d_5_ DECAP_INV_G11
XG14223 XI11_1/XI0/XI0_15/d__4_ XI11_1/XI0/XI0_15/d_4_ DECAP_INV_G11
XG14224 XI11_1/XI0/XI0_15/d__3_ XI11_1/XI0/XI0_15/d_3_ DECAP_INV_G11
XG14225 XI11_1/XI0/XI0_15/d__2_ XI11_1/XI0/XI0_15/d_2_ DECAP_INV_G11
XG14226 XI11_1/XI0/XI0_15/d__1_ XI11_1/XI0/XI0_15/d_1_ DECAP_INV_G11
XG14227 XI11_1/XI0/XI0_15/d__0_ XI11_1/XI0/XI0_15/d_0_ DECAP_INV_G11
XG14228 XI11_1/XI0/XI0_15/d_15_ XI11_1/XI0/XI0_15/d__15_ DECAP_INV_G11
XG14229 XI11_1/XI0/XI0_15/d_14_ XI11_1/XI0/XI0_15/d__14_ DECAP_INV_G11
XG14230 XI11_1/XI0/XI0_15/d_13_ XI11_1/XI0/XI0_15/d__13_ DECAP_INV_G11
XG14231 XI11_1/XI0/XI0_15/d_12_ XI11_1/XI0/XI0_15/d__12_ DECAP_INV_G11
XG14232 XI11_1/XI0/XI0_15/d_11_ XI11_1/XI0/XI0_15/d__11_ DECAP_INV_G11
XG14233 XI11_1/XI0/XI0_15/d_10_ XI11_1/XI0/XI0_15/d__10_ DECAP_INV_G11
XG14234 XI11_1/XI0/XI0_15/d_9_ XI11_1/XI0/XI0_15/d__9_ DECAP_INV_G11
XG14235 XI11_1/XI0/XI0_15/d_8_ XI11_1/XI0/XI0_15/d__8_ DECAP_INV_G11
XG14236 XI11_1/XI0/XI0_15/d_7_ XI11_1/XI0/XI0_15/d__7_ DECAP_INV_G11
XG14237 XI11_1/XI0/XI0_15/d_6_ XI11_1/XI0/XI0_15/d__6_ DECAP_INV_G11
XG14238 XI11_1/XI0/XI0_15/d_5_ XI11_1/XI0/XI0_15/d__5_ DECAP_INV_G11
XG14239 XI11_1/XI0/XI0_15/d_4_ XI11_1/XI0/XI0_15/d__4_ DECAP_INV_G11
XG14240 XI11_1/XI0/XI0_15/d_3_ XI11_1/XI0/XI0_15/d__3_ DECAP_INV_G11
XG14241 XI11_1/XI0/XI0_15/d_2_ XI11_1/XI0/XI0_15/d__2_ DECAP_INV_G11
XG14242 XI11_1/XI0/XI0_15/d_1_ XI11_1/XI0/XI0_15/d__1_ DECAP_INV_G11
XG14243 XI11_1/XI0/XI0_15/d_0_ XI11_1/XI0/XI0_15/d__0_ DECAP_INV_G11
XG14244 XI11_1/XI0/XI0_14/d__15_ XI11_1/XI0/XI0_14/d_15_ DECAP_INV_G11
XG14245 XI11_1/XI0/XI0_14/d__14_ XI11_1/XI0/XI0_14/d_14_ DECAP_INV_G11
XG14246 XI11_1/XI0/XI0_14/d__13_ XI11_1/XI0/XI0_14/d_13_ DECAP_INV_G11
XG14247 XI11_1/XI0/XI0_14/d__12_ XI11_1/XI0/XI0_14/d_12_ DECAP_INV_G11
XG14248 XI11_1/XI0/XI0_14/d__11_ XI11_1/XI0/XI0_14/d_11_ DECAP_INV_G11
XG14249 XI11_1/XI0/XI0_14/d__10_ XI11_1/XI0/XI0_14/d_10_ DECAP_INV_G11
XG14250 XI11_1/XI0/XI0_14/d__9_ XI11_1/XI0/XI0_14/d_9_ DECAP_INV_G11
XG14251 XI11_1/XI0/XI0_14/d__8_ XI11_1/XI0/XI0_14/d_8_ DECAP_INV_G11
XG14252 XI11_1/XI0/XI0_14/d__7_ XI11_1/XI0/XI0_14/d_7_ DECAP_INV_G11
XG14253 XI11_1/XI0/XI0_14/d__6_ XI11_1/XI0/XI0_14/d_6_ DECAP_INV_G11
XG14254 XI11_1/XI0/XI0_14/d__5_ XI11_1/XI0/XI0_14/d_5_ DECAP_INV_G11
XG14255 XI11_1/XI0/XI0_14/d__4_ XI11_1/XI0/XI0_14/d_4_ DECAP_INV_G11
XG14256 XI11_1/XI0/XI0_14/d__3_ XI11_1/XI0/XI0_14/d_3_ DECAP_INV_G11
XG14257 XI11_1/XI0/XI0_14/d__2_ XI11_1/XI0/XI0_14/d_2_ DECAP_INV_G11
XG14258 XI11_1/XI0/XI0_14/d__1_ XI11_1/XI0/XI0_14/d_1_ DECAP_INV_G11
XG14259 XI11_1/XI0/XI0_14/d__0_ XI11_1/XI0/XI0_14/d_0_ DECAP_INV_G11
XG14260 XI11_1/XI0/XI0_14/d_15_ XI11_1/XI0/XI0_14/d__15_ DECAP_INV_G11
XG14261 XI11_1/XI0/XI0_14/d_14_ XI11_1/XI0/XI0_14/d__14_ DECAP_INV_G11
XG14262 XI11_1/XI0/XI0_14/d_13_ XI11_1/XI0/XI0_14/d__13_ DECAP_INV_G11
XG14263 XI11_1/XI0/XI0_14/d_12_ XI11_1/XI0/XI0_14/d__12_ DECAP_INV_G11
XG14264 XI11_1/XI0/XI0_14/d_11_ XI11_1/XI0/XI0_14/d__11_ DECAP_INV_G11
XG14265 XI11_1/XI0/XI0_14/d_10_ XI11_1/XI0/XI0_14/d__10_ DECAP_INV_G11
XG14266 XI11_1/XI0/XI0_14/d_9_ XI11_1/XI0/XI0_14/d__9_ DECAP_INV_G11
XG14267 XI11_1/XI0/XI0_14/d_8_ XI11_1/XI0/XI0_14/d__8_ DECAP_INV_G11
XG14268 XI11_1/XI0/XI0_14/d_7_ XI11_1/XI0/XI0_14/d__7_ DECAP_INV_G11
XG14269 XI11_1/XI0/XI0_14/d_6_ XI11_1/XI0/XI0_14/d__6_ DECAP_INV_G11
XG14270 XI11_1/XI0/XI0_14/d_5_ XI11_1/XI0/XI0_14/d__5_ DECAP_INV_G11
XG14271 XI11_1/XI0/XI0_14/d_4_ XI11_1/XI0/XI0_14/d__4_ DECAP_INV_G11
XG14272 XI11_1/XI0/XI0_14/d_3_ XI11_1/XI0/XI0_14/d__3_ DECAP_INV_G11
XG14273 XI11_1/XI0/XI0_14/d_2_ XI11_1/XI0/XI0_14/d__2_ DECAP_INV_G11
XG14274 XI11_1/XI0/XI0_14/d_1_ XI11_1/XI0/XI0_14/d__1_ DECAP_INV_G11
XG14275 XI11_1/XI0/XI0_14/d_0_ XI11_1/XI0/XI0_14/d__0_ DECAP_INV_G11
XG14276 XI11_1/XI0/XI0_13/d__15_ XI11_1/XI0/XI0_13/d_15_ DECAP_INV_G11
XG14277 XI11_1/XI0/XI0_13/d__14_ XI11_1/XI0/XI0_13/d_14_ DECAP_INV_G11
XG14278 XI11_1/XI0/XI0_13/d__13_ XI11_1/XI0/XI0_13/d_13_ DECAP_INV_G11
XG14279 XI11_1/XI0/XI0_13/d__12_ XI11_1/XI0/XI0_13/d_12_ DECAP_INV_G11
XG14280 XI11_1/XI0/XI0_13/d__11_ XI11_1/XI0/XI0_13/d_11_ DECAP_INV_G11
XG14281 XI11_1/XI0/XI0_13/d__10_ XI11_1/XI0/XI0_13/d_10_ DECAP_INV_G11
XG14282 XI11_1/XI0/XI0_13/d__9_ XI11_1/XI0/XI0_13/d_9_ DECAP_INV_G11
XG14283 XI11_1/XI0/XI0_13/d__8_ XI11_1/XI0/XI0_13/d_8_ DECAP_INV_G11
XG14284 XI11_1/XI0/XI0_13/d__7_ XI11_1/XI0/XI0_13/d_7_ DECAP_INV_G11
XG14285 XI11_1/XI0/XI0_13/d__6_ XI11_1/XI0/XI0_13/d_6_ DECAP_INV_G11
XG14286 XI11_1/XI0/XI0_13/d__5_ XI11_1/XI0/XI0_13/d_5_ DECAP_INV_G11
XG14287 XI11_1/XI0/XI0_13/d__4_ XI11_1/XI0/XI0_13/d_4_ DECAP_INV_G11
XG14288 XI11_1/XI0/XI0_13/d__3_ XI11_1/XI0/XI0_13/d_3_ DECAP_INV_G11
XG14289 XI11_1/XI0/XI0_13/d__2_ XI11_1/XI0/XI0_13/d_2_ DECAP_INV_G11
XG14290 XI11_1/XI0/XI0_13/d__1_ XI11_1/XI0/XI0_13/d_1_ DECAP_INV_G11
XG14291 XI11_1/XI0/XI0_13/d__0_ XI11_1/XI0/XI0_13/d_0_ DECAP_INV_G11
XG14292 XI11_1/XI0/XI0_13/d_15_ XI11_1/XI0/XI0_13/d__15_ DECAP_INV_G11
XG14293 XI11_1/XI0/XI0_13/d_14_ XI11_1/XI0/XI0_13/d__14_ DECAP_INV_G11
XG14294 XI11_1/XI0/XI0_13/d_13_ XI11_1/XI0/XI0_13/d__13_ DECAP_INV_G11
XG14295 XI11_1/XI0/XI0_13/d_12_ XI11_1/XI0/XI0_13/d__12_ DECAP_INV_G11
XG14296 XI11_1/XI0/XI0_13/d_11_ XI11_1/XI0/XI0_13/d__11_ DECAP_INV_G11
XG14297 XI11_1/XI0/XI0_13/d_10_ XI11_1/XI0/XI0_13/d__10_ DECAP_INV_G11
XG14298 XI11_1/XI0/XI0_13/d_9_ XI11_1/XI0/XI0_13/d__9_ DECAP_INV_G11
XG14299 XI11_1/XI0/XI0_13/d_8_ XI11_1/XI0/XI0_13/d__8_ DECAP_INV_G11
XG14300 XI11_1/XI0/XI0_13/d_7_ XI11_1/XI0/XI0_13/d__7_ DECAP_INV_G11
XG14301 XI11_1/XI0/XI0_13/d_6_ XI11_1/XI0/XI0_13/d__6_ DECAP_INV_G11
XG14302 XI11_1/XI0/XI0_13/d_5_ XI11_1/XI0/XI0_13/d__5_ DECAP_INV_G11
XG14303 XI11_1/XI0/XI0_13/d_4_ XI11_1/XI0/XI0_13/d__4_ DECAP_INV_G11
XG14304 XI11_1/XI0/XI0_13/d_3_ XI11_1/XI0/XI0_13/d__3_ DECAP_INV_G11
XG14305 XI11_1/XI0/XI0_13/d_2_ XI11_1/XI0/XI0_13/d__2_ DECAP_INV_G11
XG14306 XI11_1/XI0/XI0_13/d_1_ XI11_1/XI0/XI0_13/d__1_ DECAP_INV_G11
XG14307 XI11_1/XI0/XI0_13/d_0_ XI11_1/XI0/XI0_13/d__0_ DECAP_INV_G11
XG14308 XI11_1/XI0/XI0_12/d__15_ XI11_1/XI0/XI0_12/d_15_ DECAP_INV_G11
XG14309 XI11_1/XI0/XI0_12/d__14_ XI11_1/XI0/XI0_12/d_14_ DECAP_INV_G11
XG14310 XI11_1/XI0/XI0_12/d__13_ XI11_1/XI0/XI0_12/d_13_ DECAP_INV_G11
XG14311 XI11_1/XI0/XI0_12/d__12_ XI11_1/XI0/XI0_12/d_12_ DECAP_INV_G11
XG14312 XI11_1/XI0/XI0_12/d__11_ XI11_1/XI0/XI0_12/d_11_ DECAP_INV_G11
XG14313 XI11_1/XI0/XI0_12/d__10_ XI11_1/XI0/XI0_12/d_10_ DECAP_INV_G11
XG14314 XI11_1/XI0/XI0_12/d__9_ XI11_1/XI0/XI0_12/d_9_ DECAP_INV_G11
XG14315 XI11_1/XI0/XI0_12/d__8_ XI11_1/XI0/XI0_12/d_8_ DECAP_INV_G11
XG14316 XI11_1/XI0/XI0_12/d__7_ XI11_1/XI0/XI0_12/d_7_ DECAP_INV_G11
XG14317 XI11_1/XI0/XI0_12/d__6_ XI11_1/XI0/XI0_12/d_6_ DECAP_INV_G11
XG14318 XI11_1/XI0/XI0_12/d__5_ XI11_1/XI0/XI0_12/d_5_ DECAP_INV_G11
XG14319 XI11_1/XI0/XI0_12/d__4_ XI11_1/XI0/XI0_12/d_4_ DECAP_INV_G11
XG14320 XI11_1/XI0/XI0_12/d__3_ XI11_1/XI0/XI0_12/d_3_ DECAP_INV_G11
XG14321 XI11_1/XI0/XI0_12/d__2_ XI11_1/XI0/XI0_12/d_2_ DECAP_INV_G11
XG14322 XI11_1/XI0/XI0_12/d__1_ XI11_1/XI0/XI0_12/d_1_ DECAP_INV_G11
XG14323 XI11_1/XI0/XI0_12/d__0_ XI11_1/XI0/XI0_12/d_0_ DECAP_INV_G11
XG14324 XI11_1/XI0/XI0_12/d_15_ XI11_1/XI0/XI0_12/d__15_ DECAP_INV_G11
XG14325 XI11_1/XI0/XI0_12/d_14_ XI11_1/XI0/XI0_12/d__14_ DECAP_INV_G11
XG14326 XI11_1/XI0/XI0_12/d_13_ XI11_1/XI0/XI0_12/d__13_ DECAP_INV_G11
XG14327 XI11_1/XI0/XI0_12/d_12_ XI11_1/XI0/XI0_12/d__12_ DECAP_INV_G11
XG14328 XI11_1/XI0/XI0_12/d_11_ XI11_1/XI0/XI0_12/d__11_ DECAP_INV_G11
XG14329 XI11_1/XI0/XI0_12/d_10_ XI11_1/XI0/XI0_12/d__10_ DECAP_INV_G11
XG14330 XI11_1/XI0/XI0_12/d_9_ XI11_1/XI0/XI0_12/d__9_ DECAP_INV_G11
XG14331 XI11_1/XI0/XI0_12/d_8_ XI11_1/XI0/XI0_12/d__8_ DECAP_INV_G11
XG14332 XI11_1/XI0/XI0_12/d_7_ XI11_1/XI0/XI0_12/d__7_ DECAP_INV_G11
XG14333 XI11_1/XI0/XI0_12/d_6_ XI11_1/XI0/XI0_12/d__6_ DECAP_INV_G11
XG14334 XI11_1/XI0/XI0_12/d_5_ XI11_1/XI0/XI0_12/d__5_ DECAP_INV_G11
XG14335 XI11_1/XI0/XI0_12/d_4_ XI11_1/XI0/XI0_12/d__4_ DECAP_INV_G11
XG14336 XI11_1/XI0/XI0_12/d_3_ XI11_1/XI0/XI0_12/d__3_ DECAP_INV_G11
XG14337 XI11_1/XI0/XI0_12/d_2_ XI11_1/XI0/XI0_12/d__2_ DECAP_INV_G11
XG14338 XI11_1/XI0/XI0_12/d_1_ XI11_1/XI0/XI0_12/d__1_ DECAP_INV_G11
XG14339 XI11_1/XI0/XI0_12/d_0_ XI11_1/XI0/XI0_12/d__0_ DECAP_INV_G11
XG14340 XI11_1/XI0/XI0_11/d__15_ XI11_1/XI0/XI0_11/d_15_ DECAP_INV_G11
XG14341 XI11_1/XI0/XI0_11/d__14_ XI11_1/XI0/XI0_11/d_14_ DECAP_INV_G11
XG14342 XI11_1/XI0/XI0_11/d__13_ XI11_1/XI0/XI0_11/d_13_ DECAP_INV_G11
XG14343 XI11_1/XI0/XI0_11/d__12_ XI11_1/XI0/XI0_11/d_12_ DECAP_INV_G11
XG14344 XI11_1/XI0/XI0_11/d__11_ XI11_1/XI0/XI0_11/d_11_ DECAP_INV_G11
XG14345 XI11_1/XI0/XI0_11/d__10_ XI11_1/XI0/XI0_11/d_10_ DECAP_INV_G11
XG14346 XI11_1/XI0/XI0_11/d__9_ XI11_1/XI0/XI0_11/d_9_ DECAP_INV_G11
XG14347 XI11_1/XI0/XI0_11/d__8_ XI11_1/XI0/XI0_11/d_8_ DECAP_INV_G11
XG14348 XI11_1/XI0/XI0_11/d__7_ XI11_1/XI0/XI0_11/d_7_ DECAP_INV_G11
XG14349 XI11_1/XI0/XI0_11/d__6_ XI11_1/XI0/XI0_11/d_6_ DECAP_INV_G11
XG14350 XI11_1/XI0/XI0_11/d__5_ XI11_1/XI0/XI0_11/d_5_ DECAP_INV_G11
XG14351 XI11_1/XI0/XI0_11/d__4_ XI11_1/XI0/XI0_11/d_4_ DECAP_INV_G11
XG14352 XI11_1/XI0/XI0_11/d__3_ XI11_1/XI0/XI0_11/d_3_ DECAP_INV_G11
XG14353 XI11_1/XI0/XI0_11/d__2_ XI11_1/XI0/XI0_11/d_2_ DECAP_INV_G11
XG14354 XI11_1/XI0/XI0_11/d__1_ XI11_1/XI0/XI0_11/d_1_ DECAP_INV_G11
XG14355 XI11_1/XI0/XI0_11/d__0_ XI11_1/XI0/XI0_11/d_0_ DECAP_INV_G11
XG14356 XI11_1/XI0/XI0_11/d_15_ XI11_1/XI0/XI0_11/d__15_ DECAP_INV_G11
XG14357 XI11_1/XI0/XI0_11/d_14_ XI11_1/XI0/XI0_11/d__14_ DECAP_INV_G11
XG14358 XI11_1/XI0/XI0_11/d_13_ XI11_1/XI0/XI0_11/d__13_ DECAP_INV_G11
XG14359 XI11_1/XI0/XI0_11/d_12_ XI11_1/XI0/XI0_11/d__12_ DECAP_INV_G11
XG14360 XI11_1/XI0/XI0_11/d_11_ XI11_1/XI0/XI0_11/d__11_ DECAP_INV_G11
XG14361 XI11_1/XI0/XI0_11/d_10_ XI11_1/XI0/XI0_11/d__10_ DECAP_INV_G11
XG14362 XI11_1/XI0/XI0_11/d_9_ XI11_1/XI0/XI0_11/d__9_ DECAP_INV_G11
XG14363 XI11_1/XI0/XI0_11/d_8_ XI11_1/XI0/XI0_11/d__8_ DECAP_INV_G11
XG14364 XI11_1/XI0/XI0_11/d_7_ XI11_1/XI0/XI0_11/d__7_ DECAP_INV_G11
XG14365 XI11_1/XI0/XI0_11/d_6_ XI11_1/XI0/XI0_11/d__6_ DECAP_INV_G11
XG14366 XI11_1/XI0/XI0_11/d_5_ XI11_1/XI0/XI0_11/d__5_ DECAP_INV_G11
XG14367 XI11_1/XI0/XI0_11/d_4_ XI11_1/XI0/XI0_11/d__4_ DECAP_INV_G11
XG14368 XI11_1/XI0/XI0_11/d_3_ XI11_1/XI0/XI0_11/d__3_ DECAP_INV_G11
XG14369 XI11_1/XI0/XI0_11/d_2_ XI11_1/XI0/XI0_11/d__2_ DECAP_INV_G11
XG14370 XI11_1/XI0/XI0_11/d_1_ XI11_1/XI0/XI0_11/d__1_ DECAP_INV_G11
XG14371 XI11_1/XI0/XI0_11/d_0_ XI11_1/XI0/XI0_11/d__0_ DECAP_INV_G11
XG14372 XI11_1/XI0/XI0_10/d__15_ XI11_1/XI0/XI0_10/d_15_ DECAP_INV_G11
XG14373 XI11_1/XI0/XI0_10/d__14_ XI11_1/XI0/XI0_10/d_14_ DECAP_INV_G11
XG14374 XI11_1/XI0/XI0_10/d__13_ XI11_1/XI0/XI0_10/d_13_ DECAP_INV_G11
XG14375 XI11_1/XI0/XI0_10/d__12_ XI11_1/XI0/XI0_10/d_12_ DECAP_INV_G11
XG14376 XI11_1/XI0/XI0_10/d__11_ XI11_1/XI0/XI0_10/d_11_ DECAP_INV_G11
XG14377 XI11_1/XI0/XI0_10/d__10_ XI11_1/XI0/XI0_10/d_10_ DECAP_INV_G11
XG14378 XI11_1/XI0/XI0_10/d__9_ XI11_1/XI0/XI0_10/d_9_ DECAP_INV_G11
XG14379 XI11_1/XI0/XI0_10/d__8_ XI11_1/XI0/XI0_10/d_8_ DECAP_INV_G11
XG14380 XI11_1/XI0/XI0_10/d__7_ XI11_1/XI0/XI0_10/d_7_ DECAP_INV_G11
XG14381 XI11_1/XI0/XI0_10/d__6_ XI11_1/XI0/XI0_10/d_6_ DECAP_INV_G11
XG14382 XI11_1/XI0/XI0_10/d__5_ XI11_1/XI0/XI0_10/d_5_ DECAP_INV_G11
XG14383 XI11_1/XI0/XI0_10/d__4_ XI11_1/XI0/XI0_10/d_4_ DECAP_INV_G11
XG14384 XI11_1/XI0/XI0_10/d__3_ XI11_1/XI0/XI0_10/d_3_ DECAP_INV_G11
XG14385 XI11_1/XI0/XI0_10/d__2_ XI11_1/XI0/XI0_10/d_2_ DECAP_INV_G11
XG14386 XI11_1/XI0/XI0_10/d__1_ XI11_1/XI0/XI0_10/d_1_ DECAP_INV_G11
XG14387 XI11_1/XI0/XI0_10/d__0_ XI11_1/XI0/XI0_10/d_0_ DECAP_INV_G11
XG14388 XI11_1/XI0/XI0_10/d_15_ XI11_1/XI0/XI0_10/d__15_ DECAP_INV_G11
XG14389 XI11_1/XI0/XI0_10/d_14_ XI11_1/XI0/XI0_10/d__14_ DECAP_INV_G11
XG14390 XI11_1/XI0/XI0_10/d_13_ XI11_1/XI0/XI0_10/d__13_ DECAP_INV_G11
XG14391 XI11_1/XI0/XI0_10/d_12_ XI11_1/XI0/XI0_10/d__12_ DECAP_INV_G11
XG14392 XI11_1/XI0/XI0_10/d_11_ XI11_1/XI0/XI0_10/d__11_ DECAP_INV_G11
XG14393 XI11_1/XI0/XI0_10/d_10_ XI11_1/XI0/XI0_10/d__10_ DECAP_INV_G11
XG14394 XI11_1/XI0/XI0_10/d_9_ XI11_1/XI0/XI0_10/d__9_ DECAP_INV_G11
XG14395 XI11_1/XI0/XI0_10/d_8_ XI11_1/XI0/XI0_10/d__8_ DECAP_INV_G11
XG14396 XI11_1/XI0/XI0_10/d_7_ XI11_1/XI0/XI0_10/d__7_ DECAP_INV_G11
XG14397 XI11_1/XI0/XI0_10/d_6_ XI11_1/XI0/XI0_10/d__6_ DECAP_INV_G11
XG14398 XI11_1/XI0/XI0_10/d_5_ XI11_1/XI0/XI0_10/d__5_ DECAP_INV_G11
XG14399 XI11_1/XI0/XI0_10/d_4_ XI11_1/XI0/XI0_10/d__4_ DECAP_INV_G11
XG14400 XI11_1/XI0/XI0_10/d_3_ XI11_1/XI0/XI0_10/d__3_ DECAP_INV_G11
XG14401 XI11_1/XI0/XI0_10/d_2_ XI11_1/XI0/XI0_10/d__2_ DECAP_INV_G11
XG14402 XI11_1/XI0/XI0_10/d_1_ XI11_1/XI0/XI0_10/d__1_ DECAP_INV_G11
XG14403 XI11_1/XI0/XI0_10/d_0_ XI11_1/XI0/XI0_10/d__0_ DECAP_INV_G11
XG14404 XI11_1/XI0/XI0_9/d__15_ XI11_1/XI0/XI0_9/d_15_ DECAP_INV_G11
XG14405 XI11_1/XI0/XI0_9/d__14_ XI11_1/XI0/XI0_9/d_14_ DECAP_INV_G11
XG14406 XI11_1/XI0/XI0_9/d__13_ XI11_1/XI0/XI0_9/d_13_ DECAP_INV_G11
XG14407 XI11_1/XI0/XI0_9/d__12_ XI11_1/XI0/XI0_9/d_12_ DECAP_INV_G11
XG14408 XI11_1/XI0/XI0_9/d__11_ XI11_1/XI0/XI0_9/d_11_ DECAP_INV_G11
XG14409 XI11_1/XI0/XI0_9/d__10_ XI11_1/XI0/XI0_9/d_10_ DECAP_INV_G11
XG14410 XI11_1/XI0/XI0_9/d__9_ XI11_1/XI0/XI0_9/d_9_ DECAP_INV_G11
XG14411 XI11_1/XI0/XI0_9/d__8_ XI11_1/XI0/XI0_9/d_8_ DECAP_INV_G11
XG14412 XI11_1/XI0/XI0_9/d__7_ XI11_1/XI0/XI0_9/d_7_ DECAP_INV_G11
XG14413 XI11_1/XI0/XI0_9/d__6_ XI11_1/XI0/XI0_9/d_6_ DECAP_INV_G11
XG14414 XI11_1/XI0/XI0_9/d__5_ XI11_1/XI0/XI0_9/d_5_ DECAP_INV_G11
XG14415 XI11_1/XI0/XI0_9/d__4_ XI11_1/XI0/XI0_9/d_4_ DECAP_INV_G11
XG14416 XI11_1/XI0/XI0_9/d__3_ XI11_1/XI0/XI0_9/d_3_ DECAP_INV_G11
XG14417 XI11_1/XI0/XI0_9/d__2_ XI11_1/XI0/XI0_9/d_2_ DECAP_INV_G11
XG14418 XI11_1/XI0/XI0_9/d__1_ XI11_1/XI0/XI0_9/d_1_ DECAP_INV_G11
XG14419 XI11_1/XI0/XI0_9/d__0_ XI11_1/XI0/XI0_9/d_0_ DECAP_INV_G11
XG14420 XI11_1/XI0/XI0_9/d_15_ XI11_1/XI0/XI0_9/d__15_ DECAP_INV_G11
XG14421 XI11_1/XI0/XI0_9/d_14_ XI11_1/XI0/XI0_9/d__14_ DECAP_INV_G11
XG14422 XI11_1/XI0/XI0_9/d_13_ XI11_1/XI0/XI0_9/d__13_ DECAP_INV_G11
XG14423 XI11_1/XI0/XI0_9/d_12_ XI11_1/XI0/XI0_9/d__12_ DECAP_INV_G11
XG14424 XI11_1/XI0/XI0_9/d_11_ XI11_1/XI0/XI0_9/d__11_ DECAP_INV_G11
XG14425 XI11_1/XI0/XI0_9/d_10_ XI11_1/XI0/XI0_9/d__10_ DECAP_INV_G11
XG14426 XI11_1/XI0/XI0_9/d_9_ XI11_1/XI0/XI0_9/d__9_ DECAP_INV_G11
XG14427 XI11_1/XI0/XI0_9/d_8_ XI11_1/XI0/XI0_9/d__8_ DECAP_INV_G11
XG14428 XI11_1/XI0/XI0_9/d_7_ XI11_1/XI0/XI0_9/d__7_ DECAP_INV_G11
XG14429 XI11_1/XI0/XI0_9/d_6_ XI11_1/XI0/XI0_9/d__6_ DECAP_INV_G11
XG14430 XI11_1/XI0/XI0_9/d_5_ XI11_1/XI0/XI0_9/d__5_ DECAP_INV_G11
XG14431 XI11_1/XI0/XI0_9/d_4_ XI11_1/XI0/XI0_9/d__4_ DECAP_INV_G11
XG14432 XI11_1/XI0/XI0_9/d_3_ XI11_1/XI0/XI0_9/d__3_ DECAP_INV_G11
XG14433 XI11_1/XI0/XI0_9/d_2_ XI11_1/XI0/XI0_9/d__2_ DECAP_INV_G11
XG14434 XI11_1/XI0/XI0_9/d_1_ XI11_1/XI0/XI0_9/d__1_ DECAP_INV_G11
XG14435 XI11_1/XI0/XI0_9/d_0_ XI11_1/XI0/XI0_9/d__0_ DECAP_INV_G11
XG14436 XI11_1/XI0/XI0_8/d__15_ XI11_1/XI0/XI0_8/d_15_ DECAP_INV_G11
XG14437 XI11_1/XI0/XI0_8/d__14_ XI11_1/XI0/XI0_8/d_14_ DECAP_INV_G11
XG14438 XI11_1/XI0/XI0_8/d__13_ XI11_1/XI0/XI0_8/d_13_ DECAP_INV_G11
XG14439 XI11_1/XI0/XI0_8/d__12_ XI11_1/XI0/XI0_8/d_12_ DECAP_INV_G11
XG14440 XI11_1/XI0/XI0_8/d__11_ XI11_1/XI0/XI0_8/d_11_ DECAP_INV_G11
XG14441 XI11_1/XI0/XI0_8/d__10_ XI11_1/XI0/XI0_8/d_10_ DECAP_INV_G11
XG14442 XI11_1/XI0/XI0_8/d__9_ XI11_1/XI0/XI0_8/d_9_ DECAP_INV_G11
XG14443 XI11_1/XI0/XI0_8/d__8_ XI11_1/XI0/XI0_8/d_8_ DECAP_INV_G11
XG14444 XI11_1/XI0/XI0_8/d__7_ XI11_1/XI0/XI0_8/d_7_ DECAP_INV_G11
XG14445 XI11_1/XI0/XI0_8/d__6_ XI11_1/XI0/XI0_8/d_6_ DECAP_INV_G11
XG14446 XI11_1/XI0/XI0_8/d__5_ XI11_1/XI0/XI0_8/d_5_ DECAP_INV_G11
XG14447 XI11_1/XI0/XI0_8/d__4_ XI11_1/XI0/XI0_8/d_4_ DECAP_INV_G11
XG14448 XI11_1/XI0/XI0_8/d__3_ XI11_1/XI0/XI0_8/d_3_ DECAP_INV_G11
XG14449 XI11_1/XI0/XI0_8/d__2_ XI11_1/XI0/XI0_8/d_2_ DECAP_INV_G11
XG14450 XI11_1/XI0/XI0_8/d__1_ XI11_1/XI0/XI0_8/d_1_ DECAP_INV_G11
XG14451 XI11_1/XI0/XI0_8/d__0_ XI11_1/XI0/XI0_8/d_0_ DECAP_INV_G11
XG14452 XI11_1/XI0/XI0_8/d_15_ XI11_1/XI0/XI0_8/d__15_ DECAP_INV_G11
XG14453 XI11_1/XI0/XI0_8/d_14_ XI11_1/XI0/XI0_8/d__14_ DECAP_INV_G11
XG14454 XI11_1/XI0/XI0_8/d_13_ XI11_1/XI0/XI0_8/d__13_ DECAP_INV_G11
XG14455 XI11_1/XI0/XI0_8/d_12_ XI11_1/XI0/XI0_8/d__12_ DECAP_INV_G11
XG14456 XI11_1/XI0/XI0_8/d_11_ XI11_1/XI0/XI0_8/d__11_ DECAP_INV_G11
XG14457 XI11_1/XI0/XI0_8/d_10_ XI11_1/XI0/XI0_8/d__10_ DECAP_INV_G11
XG14458 XI11_1/XI0/XI0_8/d_9_ XI11_1/XI0/XI0_8/d__9_ DECAP_INV_G11
XG14459 XI11_1/XI0/XI0_8/d_8_ XI11_1/XI0/XI0_8/d__8_ DECAP_INV_G11
XG14460 XI11_1/XI0/XI0_8/d_7_ XI11_1/XI0/XI0_8/d__7_ DECAP_INV_G11
XG14461 XI11_1/XI0/XI0_8/d_6_ XI11_1/XI0/XI0_8/d__6_ DECAP_INV_G11
XG14462 XI11_1/XI0/XI0_8/d_5_ XI11_1/XI0/XI0_8/d__5_ DECAP_INV_G11
XG14463 XI11_1/XI0/XI0_8/d_4_ XI11_1/XI0/XI0_8/d__4_ DECAP_INV_G11
XG14464 XI11_1/XI0/XI0_8/d_3_ XI11_1/XI0/XI0_8/d__3_ DECAP_INV_G11
XG14465 XI11_1/XI0/XI0_8/d_2_ XI11_1/XI0/XI0_8/d__2_ DECAP_INV_G11
XG14466 XI11_1/XI0/XI0_8/d_1_ XI11_1/XI0/XI0_8/d__1_ DECAP_INV_G11
XG14467 XI11_1/XI0/XI0_8/d_0_ XI11_1/XI0/XI0_8/d__0_ DECAP_INV_G11
XG14468 XI11_1/XI0/XI0_7/d__15_ XI11_1/XI0/XI0_7/d_15_ DECAP_INV_G11
XG14469 XI11_1/XI0/XI0_7/d__14_ XI11_1/XI0/XI0_7/d_14_ DECAP_INV_G11
XG14470 XI11_1/XI0/XI0_7/d__13_ XI11_1/XI0/XI0_7/d_13_ DECAP_INV_G11
XG14471 XI11_1/XI0/XI0_7/d__12_ XI11_1/XI0/XI0_7/d_12_ DECAP_INV_G11
XG14472 XI11_1/XI0/XI0_7/d__11_ XI11_1/XI0/XI0_7/d_11_ DECAP_INV_G11
XG14473 XI11_1/XI0/XI0_7/d__10_ XI11_1/XI0/XI0_7/d_10_ DECAP_INV_G11
XG14474 XI11_1/XI0/XI0_7/d__9_ XI11_1/XI0/XI0_7/d_9_ DECAP_INV_G11
XG14475 XI11_1/XI0/XI0_7/d__8_ XI11_1/XI0/XI0_7/d_8_ DECAP_INV_G11
XG14476 XI11_1/XI0/XI0_7/d__7_ XI11_1/XI0/XI0_7/d_7_ DECAP_INV_G11
XG14477 XI11_1/XI0/XI0_7/d__6_ XI11_1/XI0/XI0_7/d_6_ DECAP_INV_G11
XG14478 XI11_1/XI0/XI0_7/d__5_ XI11_1/XI0/XI0_7/d_5_ DECAP_INV_G11
XG14479 XI11_1/XI0/XI0_7/d__4_ XI11_1/XI0/XI0_7/d_4_ DECAP_INV_G11
XG14480 XI11_1/XI0/XI0_7/d__3_ XI11_1/XI0/XI0_7/d_3_ DECAP_INV_G11
XG14481 XI11_1/XI0/XI0_7/d__2_ XI11_1/XI0/XI0_7/d_2_ DECAP_INV_G11
XG14482 XI11_1/XI0/XI0_7/d__1_ XI11_1/XI0/XI0_7/d_1_ DECAP_INV_G11
XG14483 XI11_1/XI0/XI0_7/d__0_ XI11_1/XI0/XI0_7/d_0_ DECAP_INV_G11
XG14484 XI11_1/XI0/XI0_7/d_15_ XI11_1/XI0/XI0_7/d__15_ DECAP_INV_G11
XG14485 XI11_1/XI0/XI0_7/d_14_ XI11_1/XI0/XI0_7/d__14_ DECAP_INV_G11
XG14486 XI11_1/XI0/XI0_7/d_13_ XI11_1/XI0/XI0_7/d__13_ DECAP_INV_G11
XG14487 XI11_1/XI0/XI0_7/d_12_ XI11_1/XI0/XI0_7/d__12_ DECAP_INV_G11
XG14488 XI11_1/XI0/XI0_7/d_11_ XI11_1/XI0/XI0_7/d__11_ DECAP_INV_G11
XG14489 XI11_1/XI0/XI0_7/d_10_ XI11_1/XI0/XI0_7/d__10_ DECAP_INV_G11
XG14490 XI11_1/XI0/XI0_7/d_9_ XI11_1/XI0/XI0_7/d__9_ DECAP_INV_G11
XG14491 XI11_1/XI0/XI0_7/d_8_ XI11_1/XI0/XI0_7/d__8_ DECAP_INV_G11
XG14492 XI11_1/XI0/XI0_7/d_7_ XI11_1/XI0/XI0_7/d__7_ DECAP_INV_G11
XG14493 XI11_1/XI0/XI0_7/d_6_ XI11_1/XI0/XI0_7/d__6_ DECAP_INV_G11
XG14494 XI11_1/XI0/XI0_7/d_5_ XI11_1/XI0/XI0_7/d__5_ DECAP_INV_G11
XG14495 XI11_1/XI0/XI0_7/d_4_ XI11_1/XI0/XI0_7/d__4_ DECAP_INV_G11
XG14496 XI11_1/XI0/XI0_7/d_3_ XI11_1/XI0/XI0_7/d__3_ DECAP_INV_G11
XG14497 XI11_1/XI0/XI0_7/d_2_ XI11_1/XI0/XI0_7/d__2_ DECAP_INV_G11
XG14498 XI11_1/XI0/XI0_7/d_1_ XI11_1/XI0/XI0_7/d__1_ DECAP_INV_G11
XG14499 XI11_1/XI0/XI0_7/d_0_ XI11_1/XI0/XI0_7/d__0_ DECAP_INV_G11
XG14500 XI11_1/XI0/XI0_6/d__15_ XI11_1/XI0/XI0_6/d_15_ DECAP_INV_G11
XG14501 XI11_1/XI0/XI0_6/d__14_ XI11_1/XI0/XI0_6/d_14_ DECAP_INV_G11
XG14502 XI11_1/XI0/XI0_6/d__13_ XI11_1/XI0/XI0_6/d_13_ DECAP_INV_G11
XG14503 XI11_1/XI0/XI0_6/d__12_ XI11_1/XI0/XI0_6/d_12_ DECAP_INV_G11
XG14504 XI11_1/XI0/XI0_6/d__11_ XI11_1/XI0/XI0_6/d_11_ DECAP_INV_G11
XG14505 XI11_1/XI0/XI0_6/d__10_ XI11_1/XI0/XI0_6/d_10_ DECAP_INV_G11
XG14506 XI11_1/XI0/XI0_6/d__9_ XI11_1/XI0/XI0_6/d_9_ DECAP_INV_G11
XG14507 XI11_1/XI0/XI0_6/d__8_ XI11_1/XI0/XI0_6/d_8_ DECAP_INV_G11
XG14508 XI11_1/XI0/XI0_6/d__7_ XI11_1/XI0/XI0_6/d_7_ DECAP_INV_G11
XG14509 XI11_1/XI0/XI0_6/d__6_ XI11_1/XI0/XI0_6/d_6_ DECAP_INV_G11
XG14510 XI11_1/XI0/XI0_6/d__5_ XI11_1/XI0/XI0_6/d_5_ DECAP_INV_G11
XG14511 XI11_1/XI0/XI0_6/d__4_ XI11_1/XI0/XI0_6/d_4_ DECAP_INV_G11
XG14512 XI11_1/XI0/XI0_6/d__3_ XI11_1/XI0/XI0_6/d_3_ DECAP_INV_G11
XG14513 XI11_1/XI0/XI0_6/d__2_ XI11_1/XI0/XI0_6/d_2_ DECAP_INV_G11
XG14514 XI11_1/XI0/XI0_6/d__1_ XI11_1/XI0/XI0_6/d_1_ DECAP_INV_G11
XG14515 XI11_1/XI0/XI0_6/d__0_ XI11_1/XI0/XI0_6/d_0_ DECAP_INV_G11
XG14516 XI11_1/XI0/XI0_6/d_15_ XI11_1/XI0/XI0_6/d__15_ DECAP_INV_G11
XG14517 XI11_1/XI0/XI0_6/d_14_ XI11_1/XI0/XI0_6/d__14_ DECAP_INV_G11
XG14518 XI11_1/XI0/XI0_6/d_13_ XI11_1/XI0/XI0_6/d__13_ DECAP_INV_G11
XG14519 XI11_1/XI0/XI0_6/d_12_ XI11_1/XI0/XI0_6/d__12_ DECAP_INV_G11
XG14520 XI11_1/XI0/XI0_6/d_11_ XI11_1/XI0/XI0_6/d__11_ DECAP_INV_G11
XG14521 XI11_1/XI0/XI0_6/d_10_ XI11_1/XI0/XI0_6/d__10_ DECAP_INV_G11
XG14522 XI11_1/XI0/XI0_6/d_9_ XI11_1/XI0/XI0_6/d__9_ DECAP_INV_G11
XG14523 XI11_1/XI0/XI0_6/d_8_ XI11_1/XI0/XI0_6/d__8_ DECAP_INV_G11
XG14524 XI11_1/XI0/XI0_6/d_7_ XI11_1/XI0/XI0_6/d__7_ DECAP_INV_G11
XG14525 XI11_1/XI0/XI0_6/d_6_ XI11_1/XI0/XI0_6/d__6_ DECAP_INV_G11
XG14526 XI11_1/XI0/XI0_6/d_5_ XI11_1/XI0/XI0_6/d__5_ DECAP_INV_G11
XG14527 XI11_1/XI0/XI0_6/d_4_ XI11_1/XI0/XI0_6/d__4_ DECAP_INV_G11
XG14528 XI11_1/XI0/XI0_6/d_3_ XI11_1/XI0/XI0_6/d__3_ DECAP_INV_G11
XG14529 XI11_1/XI0/XI0_6/d_2_ XI11_1/XI0/XI0_6/d__2_ DECAP_INV_G11
XG14530 XI11_1/XI0/XI0_6/d_1_ XI11_1/XI0/XI0_6/d__1_ DECAP_INV_G11
XG14531 XI11_1/XI0/XI0_6/d_0_ XI11_1/XI0/XI0_6/d__0_ DECAP_INV_G11
XG14532 XI11_1/XI0/XI0_5/d__15_ XI11_1/XI0/XI0_5/d_15_ DECAP_INV_G11
XG14533 XI11_1/XI0/XI0_5/d__14_ XI11_1/XI0/XI0_5/d_14_ DECAP_INV_G11
XG14534 XI11_1/XI0/XI0_5/d__13_ XI11_1/XI0/XI0_5/d_13_ DECAP_INV_G11
XG14535 XI11_1/XI0/XI0_5/d__12_ XI11_1/XI0/XI0_5/d_12_ DECAP_INV_G11
XG14536 XI11_1/XI0/XI0_5/d__11_ XI11_1/XI0/XI0_5/d_11_ DECAP_INV_G11
XG14537 XI11_1/XI0/XI0_5/d__10_ XI11_1/XI0/XI0_5/d_10_ DECAP_INV_G11
XG14538 XI11_1/XI0/XI0_5/d__9_ XI11_1/XI0/XI0_5/d_9_ DECAP_INV_G11
XG14539 XI11_1/XI0/XI0_5/d__8_ XI11_1/XI0/XI0_5/d_8_ DECAP_INV_G11
XG14540 XI11_1/XI0/XI0_5/d__7_ XI11_1/XI0/XI0_5/d_7_ DECAP_INV_G11
XG14541 XI11_1/XI0/XI0_5/d__6_ XI11_1/XI0/XI0_5/d_6_ DECAP_INV_G11
XG14542 XI11_1/XI0/XI0_5/d__5_ XI11_1/XI0/XI0_5/d_5_ DECAP_INV_G11
XG14543 XI11_1/XI0/XI0_5/d__4_ XI11_1/XI0/XI0_5/d_4_ DECAP_INV_G11
XG14544 XI11_1/XI0/XI0_5/d__3_ XI11_1/XI0/XI0_5/d_3_ DECAP_INV_G11
XG14545 XI11_1/XI0/XI0_5/d__2_ XI11_1/XI0/XI0_5/d_2_ DECAP_INV_G11
XG14546 XI11_1/XI0/XI0_5/d__1_ XI11_1/XI0/XI0_5/d_1_ DECAP_INV_G11
XG14547 XI11_1/XI0/XI0_5/d__0_ XI11_1/XI0/XI0_5/d_0_ DECAP_INV_G11
XG14548 XI11_1/XI0/XI0_5/d_15_ XI11_1/XI0/XI0_5/d__15_ DECAP_INV_G11
XG14549 XI11_1/XI0/XI0_5/d_14_ XI11_1/XI0/XI0_5/d__14_ DECAP_INV_G11
XG14550 XI11_1/XI0/XI0_5/d_13_ XI11_1/XI0/XI0_5/d__13_ DECAP_INV_G11
XG14551 XI11_1/XI0/XI0_5/d_12_ XI11_1/XI0/XI0_5/d__12_ DECAP_INV_G11
XG14552 XI11_1/XI0/XI0_5/d_11_ XI11_1/XI0/XI0_5/d__11_ DECAP_INV_G11
XG14553 XI11_1/XI0/XI0_5/d_10_ XI11_1/XI0/XI0_5/d__10_ DECAP_INV_G11
XG14554 XI11_1/XI0/XI0_5/d_9_ XI11_1/XI0/XI0_5/d__9_ DECAP_INV_G11
XG14555 XI11_1/XI0/XI0_5/d_8_ XI11_1/XI0/XI0_5/d__8_ DECAP_INV_G11
XG14556 XI11_1/XI0/XI0_5/d_7_ XI11_1/XI0/XI0_5/d__7_ DECAP_INV_G11
XG14557 XI11_1/XI0/XI0_5/d_6_ XI11_1/XI0/XI0_5/d__6_ DECAP_INV_G11
XG14558 XI11_1/XI0/XI0_5/d_5_ XI11_1/XI0/XI0_5/d__5_ DECAP_INV_G11
XG14559 XI11_1/XI0/XI0_5/d_4_ XI11_1/XI0/XI0_5/d__4_ DECAP_INV_G11
XG14560 XI11_1/XI0/XI0_5/d_3_ XI11_1/XI0/XI0_5/d__3_ DECAP_INV_G11
XG14561 XI11_1/XI0/XI0_5/d_2_ XI11_1/XI0/XI0_5/d__2_ DECAP_INV_G11
XG14562 XI11_1/XI0/XI0_5/d_1_ XI11_1/XI0/XI0_5/d__1_ DECAP_INV_G11
XG14563 XI11_1/XI0/XI0_5/d_0_ XI11_1/XI0/XI0_5/d__0_ DECAP_INV_G11
XG14564 XI11_1/XI0/XI0_4/d__15_ XI11_1/XI0/XI0_4/d_15_ DECAP_INV_G11
XG14565 XI11_1/XI0/XI0_4/d__14_ XI11_1/XI0/XI0_4/d_14_ DECAP_INV_G11
XG14566 XI11_1/XI0/XI0_4/d__13_ XI11_1/XI0/XI0_4/d_13_ DECAP_INV_G11
XG14567 XI11_1/XI0/XI0_4/d__12_ XI11_1/XI0/XI0_4/d_12_ DECAP_INV_G11
XG14568 XI11_1/XI0/XI0_4/d__11_ XI11_1/XI0/XI0_4/d_11_ DECAP_INV_G11
XG14569 XI11_1/XI0/XI0_4/d__10_ XI11_1/XI0/XI0_4/d_10_ DECAP_INV_G11
XG14570 XI11_1/XI0/XI0_4/d__9_ XI11_1/XI0/XI0_4/d_9_ DECAP_INV_G11
XG14571 XI11_1/XI0/XI0_4/d__8_ XI11_1/XI0/XI0_4/d_8_ DECAP_INV_G11
XG14572 XI11_1/XI0/XI0_4/d__7_ XI11_1/XI0/XI0_4/d_7_ DECAP_INV_G11
XG14573 XI11_1/XI0/XI0_4/d__6_ XI11_1/XI0/XI0_4/d_6_ DECAP_INV_G11
XG14574 XI11_1/XI0/XI0_4/d__5_ XI11_1/XI0/XI0_4/d_5_ DECAP_INV_G11
XG14575 XI11_1/XI0/XI0_4/d__4_ XI11_1/XI0/XI0_4/d_4_ DECAP_INV_G11
XG14576 XI11_1/XI0/XI0_4/d__3_ XI11_1/XI0/XI0_4/d_3_ DECAP_INV_G11
XG14577 XI11_1/XI0/XI0_4/d__2_ XI11_1/XI0/XI0_4/d_2_ DECAP_INV_G11
XG14578 XI11_1/XI0/XI0_4/d__1_ XI11_1/XI0/XI0_4/d_1_ DECAP_INV_G11
XG14579 XI11_1/XI0/XI0_4/d__0_ XI11_1/XI0/XI0_4/d_0_ DECAP_INV_G11
XG14580 XI11_1/XI0/XI0_4/d_15_ XI11_1/XI0/XI0_4/d__15_ DECAP_INV_G11
XG14581 XI11_1/XI0/XI0_4/d_14_ XI11_1/XI0/XI0_4/d__14_ DECAP_INV_G11
XG14582 XI11_1/XI0/XI0_4/d_13_ XI11_1/XI0/XI0_4/d__13_ DECAP_INV_G11
XG14583 XI11_1/XI0/XI0_4/d_12_ XI11_1/XI0/XI0_4/d__12_ DECAP_INV_G11
XG14584 XI11_1/XI0/XI0_4/d_11_ XI11_1/XI0/XI0_4/d__11_ DECAP_INV_G11
XG14585 XI11_1/XI0/XI0_4/d_10_ XI11_1/XI0/XI0_4/d__10_ DECAP_INV_G11
XG14586 XI11_1/XI0/XI0_4/d_9_ XI11_1/XI0/XI0_4/d__9_ DECAP_INV_G11
XG14587 XI11_1/XI0/XI0_4/d_8_ XI11_1/XI0/XI0_4/d__8_ DECAP_INV_G11
XG14588 XI11_1/XI0/XI0_4/d_7_ XI11_1/XI0/XI0_4/d__7_ DECAP_INV_G11
XG14589 XI11_1/XI0/XI0_4/d_6_ XI11_1/XI0/XI0_4/d__6_ DECAP_INV_G11
XG14590 XI11_1/XI0/XI0_4/d_5_ XI11_1/XI0/XI0_4/d__5_ DECAP_INV_G11
XG14591 XI11_1/XI0/XI0_4/d_4_ XI11_1/XI0/XI0_4/d__4_ DECAP_INV_G11
XG14592 XI11_1/XI0/XI0_4/d_3_ XI11_1/XI0/XI0_4/d__3_ DECAP_INV_G11
XG14593 XI11_1/XI0/XI0_4/d_2_ XI11_1/XI0/XI0_4/d__2_ DECAP_INV_G11
XG14594 XI11_1/XI0/XI0_4/d_1_ XI11_1/XI0/XI0_4/d__1_ DECAP_INV_G11
XG14595 XI11_1/XI0/XI0_4/d_0_ XI11_1/XI0/XI0_4/d__0_ DECAP_INV_G11
XG14596 XI11_1/XI0/XI0_3/d__15_ XI11_1/XI0/XI0_3/d_15_ DECAP_INV_G11
XG14597 XI11_1/XI0/XI0_3/d__14_ XI11_1/XI0/XI0_3/d_14_ DECAP_INV_G11
XG14598 XI11_1/XI0/XI0_3/d__13_ XI11_1/XI0/XI0_3/d_13_ DECAP_INV_G11
XG14599 XI11_1/XI0/XI0_3/d__12_ XI11_1/XI0/XI0_3/d_12_ DECAP_INV_G11
XG14600 XI11_1/XI0/XI0_3/d__11_ XI11_1/XI0/XI0_3/d_11_ DECAP_INV_G11
XG14601 XI11_1/XI0/XI0_3/d__10_ XI11_1/XI0/XI0_3/d_10_ DECAP_INV_G11
XG14602 XI11_1/XI0/XI0_3/d__9_ XI11_1/XI0/XI0_3/d_9_ DECAP_INV_G11
XG14603 XI11_1/XI0/XI0_3/d__8_ XI11_1/XI0/XI0_3/d_8_ DECAP_INV_G11
XG14604 XI11_1/XI0/XI0_3/d__7_ XI11_1/XI0/XI0_3/d_7_ DECAP_INV_G11
XG14605 XI11_1/XI0/XI0_3/d__6_ XI11_1/XI0/XI0_3/d_6_ DECAP_INV_G11
XG14606 XI11_1/XI0/XI0_3/d__5_ XI11_1/XI0/XI0_3/d_5_ DECAP_INV_G11
XG14607 XI11_1/XI0/XI0_3/d__4_ XI11_1/XI0/XI0_3/d_4_ DECAP_INV_G11
XG14608 XI11_1/XI0/XI0_3/d__3_ XI11_1/XI0/XI0_3/d_3_ DECAP_INV_G11
XG14609 XI11_1/XI0/XI0_3/d__2_ XI11_1/XI0/XI0_3/d_2_ DECAP_INV_G11
XG14610 XI11_1/XI0/XI0_3/d__1_ XI11_1/XI0/XI0_3/d_1_ DECAP_INV_G11
XG14611 XI11_1/XI0/XI0_3/d__0_ XI11_1/XI0/XI0_3/d_0_ DECAP_INV_G11
XG14612 XI11_1/XI0/XI0_3/d_15_ XI11_1/XI0/XI0_3/d__15_ DECAP_INV_G11
XG14613 XI11_1/XI0/XI0_3/d_14_ XI11_1/XI0/XI0_3/d__14_ DECAP_INV_G11
XG14614 XI11_1/XI0/XI0_3/d_13_ XI11_1/XI0/XI0_3/d__13_ DECAP_INV_G11
XG14615 XI11_1/XI0/XI0_3/d_12_ XI11_1/XI0/XI0_3/d__12_ DECAP_INV_G11
XG14616 XI11_1/XI0/XI0_3/d_11_ XI11_1/XI0/XI0_3/d__11_ DECAP_INV_G11
XG14617 XI11_1/XI0/XI0_3/d_10_ XI11_1/XI0/XI0_3/d__10_ DECAP_INV_G11
XG14618 XI11_1/XI0/XI0_3/d_9_ XI11_1/XI0/XI0_3/d__9_ DECAP_INV_G11
XG14619 XI11_1/XI0/XI0_3/d_8_ XI11_1/XI0/XI0_3/d__8_ DECAP_INV_G11
XG14620 XI11_1/XI0/XI0_3/d_7_ XI11_1/XI0/XI0_3/d__7_ DECAP_INV_G11
XG14621 XI11_1/XI0/XI0_3/d_6_ XI11_1/XI0/XI0_3/d__6_ DECAP_INV_G11
XG14622 XI11_1/XI0/XI0_3/d_5_ XI11_1/XI0/XI0_3/d__5_ DECAP_INV_G11
XG14623 XI11_1/XI0/XI0_3/d_4_ XI11_1/XI0/XI0_3/d__4_ DECAP_INV_G11
XG14624 XI11_1/XI0/XI0_3/d_3_ XI11_1/XI0/XI0_3/d__3_ DECAP_INV_G11
XG14625 XI11_1/XI0/XI0_3/d_2_ XI11_1/XI0/XI0_3/d__2_ DECAP_INV_G11
XG14626 XI11_1/XI0/XI0_3/d_1_ XI11_1/XI0/XI0_3/d__1_ DECAP_INV_G11
XG14627 XI11_1/XI0/XI0_3/d_0_ XI11_1/XI0/XI0_3/d__0_ DECAP_INV_G11
XG14628 XI11_1/XI0/XI0_2/d__15_ XI11_1/XI0/XI0_2/d_15_ DECAP_INV_G11
XG14629 XI11_1/XI0/XI0_2/d__14_ XI11_1/XI0/XI0_2/d_14_ DECAP_INV_G11
XG14630 XI11_1/XI0/XI0_2/d__13_ XI11_1/XI0/XI0_2/d_13_ DECAP_INV_G11
XG14631 XI11_1/XI0/XI0_2/d__12_ XI11_1/XI0/XI0_2/d_12_ DECAP_INV_G11
XG14632 XI11_1/XI0/XI0_2/d__11_ XI11_1/XI0/XI0_2/d_11_ DECAP_INV_G11
XG14633 XI11_1/XI0/XI0_2/d__10_ XI11_1/XI0/XI0_2/d_10_ DECAP_INV_G11
XG14634 XI11_1/XI0/XI0_2/d__9_ XI11_1/XI0/XI0_2/d_9_ DECAP_INV_G11
XG14635 XI11_1/XI0/XI0_2/d__8_ XI11_1/XI0/XI0_2/d_8_ DECAP_INV_G11
XG14636 XI11_1/XI0/XI0_2/d__7_ XI11_1/XI0/XI0_2/d_7_ DECAP_INV_G11
XG14637 XI11_1/XI0/XI0_2/d__6_ XI11_1/XI0/XI0_2/d_6_ DECAP_INV_G11
XG14638 XI11_1/XI0/XI0_2/d__5_ XI11_1/XI0/XI0_2/d_5_ DECAP_INV_G11
XG14639 XI11_1/XI0/XI0_2/d__4_ XI11_1/XI0/XI0_2/d_4_ DECAP_INV_G11
XG14640 XI11_1/XI0/XI0_2/d__3_ XI11_1/XI0/XI0_2/d_3_ DECAP_INV_G11
XG14641 XI11_1/XI0/XI0_2/d__2_ XI11_1/XI0/XI0_2/d_2_ DECAP_INV_G11
XG14642 XI11_1/XI0/XI0_2/d__1_ XI11_1/XI0/XI0_2/d_1_ DECAP_INV_G11
XG14643 XI11_1/XI0/XI0_2/d__0_ XI11_1/XI0/XI0_2/d_0_ DECAP_INV_G11
XG14644 XI11_1/XI0/XI0_2/d_15_ XI11_1/XI0/XI0_2/d__15_ DECAP_INV_G11
XG14645 XI11_1/XI0/XI0_2/d_14_ XI11_1/XI0/XI0_2/d__14_ DECAP_INV_G11
XG14646 XI11_1/XI0/XI0_2/d_13_ XI11_1/XI0/XI0_2/d__13_ DECAP_INV_G11
XG14647 XI11_1/XI0/XI0_2/d_12_ XI11_1/XI0/XI0_2/d__12_ DECAP_INV_G11
XG14648 XI11_1/XI0/XI0_2/d_11_ XI11_1/XI0/XI0_2/d__11_ DECAP_INV_G11
XG14649 XI11_1/XI0/XI0_2/d_10_ XI11_1/XI0/XI0_2/d__10_ DECAP_INV_G11
XG14650 XI11_1/XI0/XI0_2/d_9_ XI11_1/XI0/XI0_2/d__9_ DECAP_INV_G11
XG14651 XI11_1/XI0/XI0_2/d_8_ XI11_1/XI0/XI0_2/d__8_ DECAP_INV_G11
XG14652 XI11_1/XI0/XI0_2/d_7_ XI11_1/XI0/XI0_2/d__7_ DECAP_INV_G11
XG14653 XI11_1/XI0/XI0_2/d_6_ XI11_1/XI0/XI0_2/d__6_ DECAP_INV_G11
XG14654 XI11_1/XI0/XI0_2/d_5_ XI11_1/XI0/XI0_2/d__5_ DECAP_INV_G11
XG14655 XI11_1/XI0/XI0_2/d_4_ XI11_1/XI0/XI0_2/d__4_ DECAP_INV_G11
XG14656 XI11_1/XI0/XI0_2/d_3_ XI11_1/XI0/XI0_2/d__3_ DECAP_INV_G11
XG14657 XI11_1/XI0/XI0_2/d_2_ XI11_1/XI0/XI0_2/d__2_ DECAP_INV_G11
XG14658 XI11_1/XI0/XI0_2/d_1_ XI11_1/XI0/XI0_2/d__1_ DECAP_INV_G11
XG14659 XI11_1/XI0/XI0_2/d_0_ XI11_1/XI0/XI0_2/d__0_ DECAP_INV_G11
XG14660 XI11_1/XI0/XI0_1/d__15_ XI11_1/XI0/XI0_1/d_15_ DECAP_INV_G11
XG14661 XI11_1/XI0/XI0_1/d__14_ XI11_1/XI0/XI0_1/d_14_ DECAP_INV_G11
XG14662 XI11_1/XI0/XI0_1/d__13_ XI11_1/XI0/XI0_1/d_13_ DECAP_INV_G11
XG14663 XI11_1/XI0/XI0_1/d__12_ XI11_1/XI0/XI0_1/d_12_ DECAP_INV_G11
XG14664 XI11_1/XI0/XI0_1/d__11_ XI11_1/XI0/XI0_1/d_11_ DECAP_INV_G11
XG14665 XI11_1/XI0/XI0_1/d__10_ XI11_1/XI0/XI0_1/d_10_ DECAP_INV_G11
XG14666 XI11_1/XI0/XI0_1/d__9_ XI11_1/XI0/XI0_1/d_9_ DECAP_INV_G11
XG14667 XI11_1/XI0/XI0_1/d__8_ XI11_1/XI0/XI0_1/d_8_ DECAP_INV_G11
XG14668 XI11_1/XI0/XI0_1/d__7_ XI11_1/XI0/XI0_1/d_7_ DECAP_INV_G11
XG14669 XI11_1/XI0/XI0_1/d__6_ XI11_1/XI0/XI0_1/d_6_ DECAP_INV_G11
XG14670 XI11_1/XI0/XI0_1/d__5_ XI11_1/XI0/XI0_1/d_5_ DECAP_INV_G11
XG14671 XI11_1/XI0/XI0_1/d__4_ XI11_1/XI0/XI0_1/d_4_ DECAP_INV_G11
XG14672 XI11_1/XI0/XI0_1/d__3_ XI11_1/XI0/XI0_1/d_3_ DECAP_INV_G11
XG14673 XI11_1/XI0/XI0_1/d__2_ XI11_1/XI0/XI0_1/d_2_ DECAP_INV_G11
XG14674 XI11_1/XI0/XI0_1/d__1_ XI11_1/XI0/XI0_1/d_1_ DECAP_INV_G11
XG14675 XI11_1/XI0/XI0_1/d__0_ XI11_1/XI0/XI0_1/d_0_ DECAP_INV_G11
XG14676 XI11_1/XI0/XI0_1/d_15_ XI11_1/XI0/XI0_1/d__15_ DECAP_INV_G11
XG14677 XI11_1/XI0/XI0_1/d_14_ XI11_1/XI0/XI0_1/d__14_ DECAP_INV_G11
XG14678 XI11_1/XI0/XI0_1/d_13_ XI11_1/XI0/XI0_1/d__13_ DECAP_INV_G11
XG14679 XI11_1/XI0/XI0_1/d_12_ XI11_1/XI0/XI0_1/d__12_ DECAP_INV_G11
XG14680 XI11_1/XI0/XI0_1/d_11_ XI11_1/XI0/XI0_1/d__11_ DECAP_INV_G11
XG14681 XI11_1/XI0/XI0_1/d_10_ XI11_1/XI0/XI0_1/d__10_ DECAP_INV_G11
XG14682 XI11_1/XI0/XI0_1/d_9_ XI11_1/XI0/XI0_1/d__9_ DECAP_INV_G11
XG14683 XI11_1/XI0/XI0_1/d_8_ XI11_1/XI0/XI0_1/d__8_ DECAP_INV_G11
XG14684 XI11_1/XI0/XI0_1/d_7_ XI11_1/XI0/XI0_1/d__7_ DECAP_INV_G11
XG14685 XI11_1/XI0/XI0_1/d_6_ XI11_1/XI0/XI0_1/d__6_ DECAP_INV_G11
XG14686 XI11_1/XI0/XI0_1/d_5_ XI11_1/XI0/XI0_1/d__5_ DECAP_INV_G11
XG14687 XI11_1/XI0/XI0_1/d_4_ XI11_1/XI0/XI0_1/d__4_ DECAP_INV_G11
XG14688 XI11_1/XI0/XI0_1/d_3_ XI11_1/XI0/XI0_1/d__3_ DECAP_INV_G11
XG14689 XI11_1/XI0/XI0_1/d_2_ XI11_1/XI0/XI0_1/d__2_ DECAP_INV_G11
XG14690 XI11_1/XI0/XI0_1/d_1_ XI11_1/XI0/XI0_1/d__1_ DECAP_INV_G11
XG14691 XI11_1/XI0/XI0_1/d_0_ XI11_1/XI0/XI0_1/d__0_ DECAP_INV_G11
XG14692 XI11_1/XI0/XI0_0/d__15_ XI11_1/XI0/XI0_0/d_15_ DECAP_INV_G11
XG14693 XI11_1/XI0/XI0_0/d__14_ XI11_1/XI0/XI0_0/d_14_ DECAP_INV_G11
XG14694 XI11_1/XI0/XI0_0/d__13_ XI11_1/XI0/XI0_0/d_13_ DECAP_INV_G11
XG14695 XI11_1/XI0/XI0_0/d__12_ XI11_1/XI0/XI0_0/d_12_ DECAP_INV_G11
XG14696 XI11_1/XI0/XI0_0/d__11_ XI11_1/XI0/XI0_0/d_11_ DECAP_INV_G11
XG14697 XI11_1/XI0/XI0_0/d__10_ XI11_1/XI0/XI0_0/d_10_ DECAP_INV_G11
XG14698 XI11_1/XI0/XI0_0/d__9_ XI11_1/XI0/XI0_0/d_9_ DECAP_INV_G11
XG14699 XI11_1/XI0/XI0_0/d__8_ XI11_1/XI0/XI0_0/d_8_ DECAP_INV_G11
XG14700 XI11_1/XI0/XI0_0/d__7_ XI11_1/XI0/XI0_0/d_7_ DECAP_INV_G11
XG14701 XI11_1/XI0/XI0_0/d__6_ XI11_1/XI0/XI0_0/d_6_ DECAP_INV_G11
XG14702 XI11_1/XI0/XI0_0/d__5_ XI11_1/XI0/XI0_0/d_5_ DECAP_INV_G11
XG14703 XI11_1/XI0/XI0_0/d__4_ XI11_1/XI0/XI0_0/d_4_ DECAP_INV_G11
XG14704 XI11_1/XI0/XI0_0/d__3_ XI11_1/XI0/XI0_0/d_3_ DECAP_INV_G11
XG14705 XI11_1/XI0/XI0_0/d__2_ XI11_1/XI0/XI0_0/d_2_ DECAP_INV_G11
XG14706 XI11_1/XI0/XI0_0/d__1_ XI11_1/XI0/XI0_0/d_1_ DECAP_INV_G11
XG14707 XI11_1/XI0/XI0_0/d__0_ XI11_1/XI0/XI0_0/d_0_ DECAP_INV_G11
XG14708 XI11_1/XI0/XI0_0/d_15_ XI11_1/XI0/XI0_0/d__15_ DECAP_INV_G11
XG14709 XI11_1/XI0/XI0_0/d_14_ XI11_1/XI0/XI0_0/d__14_ DECAP_INV_G11
XG14710 XI11_1/XI0/XI0_0/d_13_ XI11_1/XI0/XI0_0/d__13_ DECAP_INV_G11
XG14711 XI11_1/XI0/XI0_0/d_12_ XI11_1/XI0/XI0_0/d__12_ DECAP_INV_G11
XG14712 XI11_1/XI0/XI0_0/d_11_ XI11_1/XI0/XI0_0/d__11_ DECAP_INV_G11
XG14713 XI11_1/XI0/XI0_0/d_10_ XI11_1/XI0/XI0_0/d__10_ DECAP_INV_G11
XG14714 XI11_1/XI0/XI0_0/d_9_ XI11_1/XI0/XI0_0/d__9_ DECAP_INV_G11
XG14715 XI11_1/XI0/XI0_0/d_8_ XI11_1/XI0/XI0_0/d__8_ DECAP_INV_G11
XG14716 XI11_1/XI0/XI0_0/d_7_ XI11_1/XI0/XI0_0/d__7_ DECAP_INV_G11
XG14717 XI11_1/XI0/XI0_0/d_6_ XI11_1/XI0/XI0_0/d__6_ DECAP_INV_G11
XG14718 XI11_1/XI0/XI0_0/d_5_ XI11_1/XI0/XI0_0/d__5_ DECAP_INV_G11
XG14719 XI11_1/XI0/XI0_0/d_4_ XI11_1/XI0/XI0_0/d__4_ DECAP_INV_G11
XG14720 XI11_1/XI0/XI0_0/d_3_ XI11_1/XI0/XI0_0/d__3_ DECAP_INV_G11
XG14721 XI11_1/XI0/XI0_0/d_2_ XI11_1/XI0/XI0_0/d__2_ DECAP_INV_G11
XG14722 XI11_1/XI0/XI0_0/d_1_ XI11_1/XI0/XI0_0/d__1_ DECAP_INV_G11
XG14723 XI11_1/XI0/XI0_0/d_0_ XI11_1/XI0/XI0_0/d__0_ DECAP_INV_G11
XG14724 XI11_0/XI3/net17 XI11_0/XI3/net5 DECAP_INV_G7
XG14725 XI11_0/XI3/net5 XI11_0/preck DECAP_INV_G8
XG14726 sck_bar XI11_0/XI3/net018 DECAP_INV_G9
XG14727 XI11_0/XI3/net018 XI11_0/XI3/net012 DECAP_INV_G9
XG14728 XI11_0/XI3/net014 XI11_0/XI3/net7 DECAP_INV_G9
XG14729 XI11_0/XI3/net012 XI11_0/XI3/net014 DECAP_INV_G9
XG14730 XI11_0/XI4/net063 XI11_0/XI4/net0112 DECAP_INV_G10
XG14731 XI11_0/XI4/net26 XI11_0/XI4/net089 DECAP_INV_G10
XG14732 XI11_0/XI4/data_out XI11_0/XI4/data_out_ DECAP_INV_G10
XG14733 XI11_0/XI4/net20 XI11_0/XI4/net0103 DECAP_INV_G10
XG14734 XI11_0/net12 XI11_0/XI4/net32 DECAP_INV_G7
XG14735 XI11_0/net9 XI11_0/XI4/net52 DECAP_INV_G7
XG14736 XI11_0/XI4/data_out_ XI11_0/XI4/data_out DECAP_INV_G10
XG14737 XI11_0/XI0/XI0_63/d__15_ XI11_0/XI0/XI0_63/d_15_ DECAP_INV_G11
XG14738 XI11_0/XI0/XI0_63/d__14_ XI11_0/XI0/XI0_63/d_14_ DECAP_INV_G11
XG14739 XI11_0/XI0/XI0_63/d__13_ XI11_0/XI0/XI0_63/d_13_ DECAP_INV_G11
XG14740 XI11_0/XI0/XI0_63/d__12_ XI11_0/XI0/XI0_63/d_12_ DECAP_INV_G11
XG14741 XI11_0/XI0/XI0_63/d__11_ XI11_0/XI0/XI0_63/d_11_ DECAP_INV_G11
XG14742 XI11_0/XI0/XI0_63/d__10_ XI11_0/XI0/XI0_63/d_10_ DECAP_INV_G11
XG14743 XI11_0/XI0/XI0_63/d__9_ XI11_0/XI0/XI0_63/d_9_ DECAP_INV_G11
XG14744 XI11_0/XI0/XI0_63/d__8_ XI11_0/XI0/XI0_63/d_8_ DECAP_INV_G11
XG14745 XI11_0/XI0/XI0_63/d__7_ XI11_0/XI0/XI0_63/d_7_ DECAP_INV_G11
XG14746 XI11_0/XI0/XI0_63/d__6_ XI11_0/XI0/XI0_63/d_6_ DECAP_INV_G11
XG14747 XI11_0/XI0/XI0_63/d__5_ XI11_0/XI0/XI0_63/d_5_ DECAP_INV_G11
XG14748 XI11_0/XI0/XI0_63/d__4_ XI11_0/XI0/XI0_63/d_4_ DECAP_INV_G11
XG14749 XI11_0/XI0/XI0_63/d__3_ XI11_0/XI0/XI0_63/d_3_ DECAP_INV_G11
XG14750 XI11_0/XI0/XI0_63/d__2_ XI11_0/XI0/XI0_63/d_2_ DECAP_INV_G11
XG14751 XI11_0/XI0/XI0_63/d__1_ XI11_0/XI0/XI0_63/d_1_ DECAP_INV_G11
XG14752 XI11_0/XI0/XI0_63/d__0_ XI11_0/XI0/XI0_63/d_0_ DECAP_INV_G11
XG14753 XI11_0/XI0/XI0_63/d_15_ XI11_0/XI0/XI0_63/d__15_ DECAP_INV_G11
XG14754 XI11_0/XI0/XI0_63/d_14_ XI11_0/XI0/XI0_63/d__14_ DECAP_INV_G11
XG14755 XI11_0/XI0/XI0_63/d_13_ XI11_0/XI0/XI0_63/d__13_ DECAP_INV_G11
XG14756 XI11_0/XI0/XI0_63/d_12_ XI11_0/XI0/XI0_63/d__12_ DECAP_INV_G11
XG14757 XI11_0/XI0/XI0_63/d_11_ XI11_0/XI0/XI0_63/d__11_ DECAP_INV_G11
XG14758 XI11_0/XI0/XI0_63/d_10_ XI11_0/XI0/XI0_63/d__10_ DECAP_INV_G11
XG14759 XI11_0/XI0/XI0_63/d_9_ XI11_0/XI0/XI0_63/d__9_ DECAP_INV_G11
XG14760 XI11_0/XI0/XI0_63/d_8_ XI11_0/XI0/XI0_63/d__8_ DECAP_INV_G11
XG14761 XI11_0/XI0/XI0_63/d_7_ XI11_0/XI0/XI0_63/d__7_ DECAP_INV_G11
XG14762 XI11_0/XI0/XI0_63/d_6_ XI11_0/XI0/XI0_63/d__6_ DECAP_INV_G11
XG14763 XI11_0/XI0/XI0_63/d_5_ XI11_0/XI0/XI0_63/d__5_ DECAP_INV_G11
XG14764 XI11_0/XI0/XI0_63/d_4_ XI11_0/XI0/XI0_63/d__4_ DECAP_INV_G11
XG14765 XI11_0/XI0/XI0_63/d_3_ XI11_0/XI0/XI0_63/d__3_ DECAP_INV_G11
XG14766 XI11_0/XI0/XI0_63/d_2_ XI11_0/XI0/XI0_63/d__2_ DECAP_INV_G11
XG14767 XI11_0/XI0/XI0_63/d_1_ XI11_0/XI0/XI0_63/d__1_ DECAP_INV_G11
XG14768 XI11_0/XI0/XI0_63/d_0_ XI11_0/XI0/XI0_63/d__0_ DECAP_INV_G11
XG14769 XI11_0/XI0/XI0_62/d__15_ XI11_0/XI0/XI0_62/d_15_ DECAP_INV_G11
XG14770 XI11_0/XI0/XI0_62/d__14_ XI11_0/XI0/XI0_62/d_14_ DECAP_INV_G11
XG14771 XI11_0/XI0/XI0_62/d__13_ XI11_0/XI0/XI0_62/d_13_ DECAP_INV_G11
XG14772 XI11_0/XI0/XI0_62/d__12_ XI11_0/XI0/XI0_62/d_12_ DECAP_INV_G11
XG14773 XI11_0/XI0/XI0_62/d__11_ XI11_0/XI0/XI0_62/d_11_ DECAP_INV_G11
XG14774 XI11_0/XI0/XI0_62/d__10_ XI11_0/XI0/XI0_62/d_10_ DECAP_INV_G11
XG14775 XI11_0/XI0/XI0_62/d__9_ XI11_0/XI0/XI0_62/d_9_ DECAP_INV_G11
XG14776 XI11_0/XI0/XI0_62/d__8_ XI11_0/XI0/XI0_62/d_8_ DECAP_INV_G11
XG14777 XI11_0/XI0/XI0_62/d__7_ XI11_0/XI0/XI0_62/d_7_ DECAP_INV_G11
XG14778 XI11_0/XI0/XI0_62/d__6_ XI11_0/XI0/XI0_62/d_6_ DECAP_INV_G11
XG14779 XI11_0/XI0/XI0_62/d__5_ XI11_0/XI0/XI0_62/d_5_ DECAP_INV_G11
XG14780 XI11_0/XI0/XI0_62/d__4_ XI11_0/XI0/XI0_62/d_4_ DECAP_INV_G11
XG14781 XI11_0/XI0/XI0_62/d__3_ XI11_0/XI0/XI0_62/d_3_ DECAP_INV_G11
XG14782 XI11_0/XI0/XI0_62/d__2_ XI11_0/XI0/XI0_62/d_2_ DECAP_INV_G11
XG14783 XI11_0/XI0/XI0_62/d__1_ XI11_0/XI0/XI0_62/d_1_ DECAP_INV_G11
XG14784 XI11_0/XI0/XI0_62/d__0_ XI11_0/XI0/XI0_62/d_0_ DECAP_INV_G11
XG14785 XI11_0/XI0/XI0_62/d_15_ XI11_0/XI0/XI0_62/d__15_ DECAP_INV_G11
XG14786 XI11_0/XI0/XI0_62/d_14_ XI11_0/XI0/XI0_62/d__14_ DECAP_INV_G11
XG14787 XI11_0/XI0/XI0_62/d_13_ XI11_0/XI0/XI0_62/d__13_ DECAP_INV_G11
XG14788 XI11_0/XI0/XI0_62/d_12_ XI11_0/XI0/XI0_62/d__12_ DECAP_INV_G11
XG14789 XI11_0/XI0/XI0_62/d_11_ XI11_0/XI0/XI0_62/d__11_ DECAP_INV_G11
XG14790 XI11_0/XI0/XI0_62/d_10_ XI11_0/XI0/XI0_62/d__10_ DECAP_INV_G11
XG14791 XI11_0/XI0/XI0_62/d_9_ XI11_0/XI0/XI0_62/d__9_ DECAP_INV_G11
XG14792 XI11_0/XI0/XI0_62/d_8_ XI11_0/XI0/XI0_62/d__8_ DECAP_INV_G11
XG14793 XI11_0/XI0/XI0_62/d_7_ XI11_0/XI0/XI0_62/d__7_ DECAP_INV_G11
XG14794 XI11_0/XI0/XI0_62/d_6_ XI11_0/XI0/XI0_62/d__6_ DECAP_INV_G11
XG14795 XI11_0/XI0/XI0_62/d_5_ XI11_0/XI0/XI0_62/d__5_ DECAP_INV_G11
XG14796 XI11_0/XI0/XI0_62/d_4_ XI11_0/XI0/XI0_62/d__4_ DECAP_INV_G11
XG14797 XI11_0/XI0/XI0_62/d_3_ XI11_0/XI0/XI0_62/d__3_ DECAP_INV_G11
XG14798 XI11_0/XI0/XI0_62/d_2_ XI11_0/XI0/XI0_62/d__2_ DECAP_INV_G11
XG14799 XI11_0/XI0/XI0_62/d_1_ XI11_0/XI0/XI0_62/d__1_ DECAP_INV_G11
XG14800 XI11_0/XI0/XI0_62/d_0_ XI11_0/XI0/XI0_62/d__0_ DECAP_INV_G11
XG14801 XI11_0/XI0/XI0_61/d__15_ XI11_0/XI0/XI0_61/d_15_ DECAP_INV_G11
XG14802 XI11_0/XI0/XI0_61/d__14_ XI11_0/XI0/XI0_61/d_14_ DECAP_INV_G11
XG14803 XI11_0/XI0/XI0_61/d__13_ XI11_0/XI0/XI0_61/d_13_ DECAP_INV_G11
XG14804 XI11_0/XI0/XI0_61/d__12_ XI11_0/XI0/XI0_61/d_12_ DECAP_INV_G11
XG14805 XI11_0/XI0/XI0_61/d__11_ XI11_0/XI0/XI0_61/d_11_ DECAP_INV_G11
XG14806 XI11_0/XI0/XI0_61/d__10_ XI11_0/XI0/XI0_61/d_10_ DECAP_INV_G11
XG14807 XI11_0/XI0/XI0_61/d__9_ XI11_0/XI0/XI0_61/d_9_ DECAP_INV_G11
XG14808 XI11_0/XI0/XI0_61/d__8_ XI11_0/XI0/XI0_61/d_8_ DECAP_INV_G11
XG14809 XI11_0/XI0/XI0_61/d__7_ XI11_0/XI0/XI0_61/d_7_ DECAP_INV_G11
XG14810 XI11_0/XI0/XI0_61/d__6_ XI11_0/XI0/XI0_61/d_6_ DECAP_INV_G11
XG14811 XI11_0/XI0/XI0_61/d__5_ XI11_0/XI0/XI0_61/d_5_ DECAP_INV_G11
XG14812 XI11_0/XI0/XI0_61/d__4_ XI11_0/XI0/XI0_61/d_4_ DECAP_INV_G11
XG14813 XI11_0/XI0/XI0_61/d__3_ XI11_0/XI0/XI0_61/d_3_ DECAP_INV_G11
XG14814 XI11_0/XI0/XI0_61/d__2_ XI11_0/XI0/XI0_61/d_2_ DECAP_INV_G11
XG14815 XI11_0/XI0/XI0_61/d__1_ XI11_0/XI0/XI0_61/d_1_ DECAP_INV_G11
XG14816 XI11_0/XI0/XI0_61/d__0_ XI11_0/XI0/XI0_61/d_0_ DECAP_INV_G11
XG14817 XI11_0/XI0/XI0_61/d_15_ XI11_0/XI0/XI0_61/d__15_ DECAP_INV_G11
XG14818 XI11_0/XI0/XI0_61/d_14_ XI11_0/XI0/XI0_61/d__14_ DECAP_INV_G11
XG14819 XI11_0/XI0/XI0_61/d_13_ XI11_0/XI0/XI0_61/d__13_ DECAP_INV_G11
XG14820 XI11_0/XI0/XI0_61/d_12_ XI11_0/XI0/XI0_61/d__12_ DECAP_INV_G11
XG14821 XI11_0/XI0/XI0_61/d_11_ XI11_0/XI0/XI0_61/d__11_ DECAP_INV_G11
XG14822 XI11_0/XI0/XI0_61/d_10_ XI11_0/XI0/XI0_61/d__10_ DECAP_INV_G11
XG14823 XI11_0/XI0/XI0_61/d_9_ XI11_0/XI0/XI0_61/d__9_ DECAP_INV_G11
XG14824 XI11_0/XI0/XI0_61/d_8_ XI11_0/XI0/XI0_61/d__8_ DECAP_INV_G11
XG14825 XI11_0/XI0/XI0_61/d_7_ XI11_0/XI0/XI0_61/d__7_ DECAP_INV_G11
XG14826 XI11_0/XI0/XI0_61/d_6_ XI11_0/XI0/XI0_61/d__6_ DECAP_INV_G11
XG14827 XI11_0/XI0/XI0_61/d_5_ XI11_0/XI0/XI0_61/d__5_ DECAP_INV_G11
XG14828 XI11_0/XI0/XI0_61/d_4_ XI11_0/XI0/XI0_61/d__4_ DECAP_INV_G11
XG14829 XI11_0/XI0/XI0_61/d_3_ XI11_0/XI0/XI0_61/d__3_ DECAP_INV_G11
XG14830 XI11_0/XI0/XI0_61/d_2_ XI11_0/XI0/XI0_61/d__2_ DECAP_INV_G11
XG14831 XI11_0/XI0/XI0_61/d_1_ XI11_0/XI0/XI0_61/d__1_ DECAP_INV_G11
XG14832 XI11_0/XI0/XI0_61/d_0_ XI11_0/XI0/XI0_61/d__0_ DECAP_INV_G11
XG14833 XI11_0/XI0/XI0_60/d__15_ XI11_0/XI0/XI0_60/d_15_ DECAP_INV_G11
XG14834 XI11_0/XI0/XI0_60/d__14_ XI11_0/XI0/XI0_60/d_14_ DECAP_INV_G11
XG14835 XI11_0/XI0/XI0_60/d__13_ XI11_0/XI0/XI0_60/d_13_ DECAP_INV_G11
XG14836 XI11_0/XI0/XI0_60/d__12_ XI11_0/XI0/XI0_60/d_12_ DECAP_INV_G11
XG14837 XI11_0/XI0/XI0_60/d__11_ XI11_0/XI0/XI0_60/d_11_ DECAP_INV_G11
XG14838 XI11_0/XI0/XI0_60/d__10_ XI11_0/XI0/XI0_60/d_10_ DECAP_INV_G11
XG14839 XI11_0/XI0/XI0_60/d__9_ XI11_0/XI0/XI0_60/d_9_ DECAP_INV_G11
XG14840 XI11_0/XI0/XI0_60/d__8_ XI11_0/XI0/XI0_60/d_8_ DECAP_INV_G11
XG14841 XI11_0/XI0/XI0_60/d__7_ XI11_0/XI0/XI0_60/d_7_ DECAP_INV_G11
XG14842 XI11_0/XI0/XI0_60/d__6_ XI11_0/XI0/XI0_60/d_6_ DECAP_INV_G11
XG14843 XI11_0/XI0/XI0_60/d__5_ XI11_0/XI0/XI0_60/d_5_ DECAP_INV_G11
XG14844 XI11_0/XI0/XI0_60/d__4_ XI11_0/XI0/XI0_60/d_4_ DECAP_INV_G11
XG14845 XI11_0/XI0/XI0_60/d__3_ XI11_0/XI0/XI0_60/d_3_ DECAP_INV_G11
XG14846 XI11_0/XI0/XI0_60/d__2_ XI11_0/XI0/XI0_60/d_2_ DECAP_INV_G11
XG14847 XI11_0/XI0/XI0_60/d__1_ XI11_0/XI0/XI0_60/d_1_ DECAP_INV_G11
XG14848 XI11_0/XI0/XI0_60/d__0_ XI11_0/XI0/XI0_60/d_0_ DECAP_INV_G11
XG14849 XI11_0/XI0/XI0_60/d_15_ XI11_0/XI0/XI0_60/d__15_ DECAP_INV_G11
XG14850 XI11_0/XI0/XI0_60/d_14_ XI11_0/XI0/XI0_60/d__14_ DECAP_INV_G11
XG14851 XI11_0/XI0/XI0_60/d_13_ XI11_0/XI0/XI0_60/d__13_ DECAP_INV_G11
XG14852 XI11_0/XI0/XI0_60/d_12_ XI11_0/XI0/XI0_60/d__12_ DECAP_INV_G11
XG14853 XI11_0/XI0/XI0_60/d_11_ XI11_0/XI0/XI0_60/d__11_ DECAP_INV_G11
XG14854 XI11_0/XI0/XI0_60/d_10_ XI11_0/XI0/XI0_60/d__10_ DECAP_INV_G11
XG14855 XI11_0/XI0/XI0_60/d_9_ XI11_0/XI0/XI0_60/d__9_ DECAP_INV_G11
XG14856 XI11_0/XI0/XI0_60/d_8_ XI11_0/XI0/XI0_60/d__8_ DECAP_INV_G11
XG14857 XI11_0/XI0/XI0_60/d_7_ XI11_0/XI0/XI0_60/d__7_ DECAP_INV_G11
XG14858 XI11_0/XI0/XI0_60/d_6_ XI11_0/XI0/XI0_60/d__6_ DECAP_INV_G11
XG14859 XI11_0/XI0/XI0_60/d_5_ XI11_0/XI0/XI0_60/d__5_ DECAP_INV_G11
XG14860 XI11_0/XI0/XI0_60/d_4_ XI11_0/XI0/XI0_60/d__4_ DECAP_INV_G11
XG14861 XI11_0/XI0/XI0_60/d_3_ XI11_0/XI0/XI0_60/d__3_ DECAP_INV_G11
XG14862 XI11_0/XI0/XI0_60/d_2_ XI11_0/XI0/XI0_60/d__2_ DECAP_INV_G11
XG14863 XI11_0/XI0/XI0_60/d_1_ XI11_0/XI0/XI0_60/d__1_ DECAP_INV_G11
XG14864 XI11_0/XI0/XI0_60/d_0_ XI11_0/XI0/XI0_60/d__0_ DECAP_INV_G11
XG14865 XI11_0/XI0/XI0_59/d__15_ XI11_0/XI0/XI0_59/d_15_ DECAP_INV_G11
XG14866 XI11_0/XI0/XI0_59/d__14_ XI11_0/XI0/XI0_59/d_14_ DECAP_INV_G11
XG14867 XI11_0/XI0/XI0_59/d__13_ XI11_0/XI0/XI0_59/d_13_ DECAP_INV_G11
XG14868 XI11_0/XI0/XI0_59/d__12_ XI11_0/XI0/XI0_59/d_12_ DECAP_INV_G11
XG14869 XI11_0/XI0/XI0_59/d__11_ XI11_0/XI0/XI0_59/d_11_ DECAP_INV_G11
XG14870 XI11_0/XI0/XI0_59/d__10_ XI11_0/XI0/XI0_59/d_10_ DECAP_INV_G11
XG14871 XI11_0/XI0/XI0_59/d__9_ XI11_0/XI0/XI0_59/d_9_ DECAP_INV_G11
XG14872 XI11_0/XI0/XI0_59/d__8_ XI11_0/XI0/XI0_59/d_8_ DECAP_INV_G11
XG14873 XI11_0/XI0/XI0_59/d__7_ XI11_0/XI0/XI0_59/d_7_ DECAP_INV_G11
XG14874 XI11_0/XI0/XI0_59/d__6_ XI11_0/XI0/XI0_59/d_6_ DECAP_INV_G11
XG14875 XI11_0/XI0/XI0_59/d__5_ XI11_0/XI0/XI0_59/d_5_ DECAP_INV_G11
XG14876 XI11_0/XI0/XI0_59/d__4_ XI11_0/XI0/XI0_59/d_4_ DECAP_INV_G11
XG14877 XI11_0/XI0/XI0_59/d__3_ XI11_0/XI0/XI0_59/d_3_ DECAP_INV_G11
XG14878 XI11_0/XI0/XI0_59/d__2_ XI11_0/XI0/XI0_59/d_2_ DECAP_INV_G11
XG14879 XI11_0/XI0/XI0_59/d__1_ XI11_0/XI0/XI0_59/d_1_ DECAP_INV_G11
XG14880 XI11_0/XI0/XI0_59/d__0_ XI11_0/XI0/XI0_59/d_0_ DECAP_INV_G11
XG14881 XI11_0/XI0/XI0_59/d_15_ XI11_0/XI0/XI0_59/d__15_ DECAP_INV_G11
XG14882 XI11_0/XI0/XI0_59/d_14_ XI11_0/XI0/XI0_59/d__14_ DECAP_INV_G11
XG14883 XI11_0/XI0/XI0_59/d_13_ XI11_0/XI0/XI0_59/d__13_ DECAP_INV_G11
XG14884 XI11_0/XI0/XI0_59/d_12_ XI11_0/XI0/XI0_59/d__12_ DECAP_INV_G11
XG14885 XI11_0/XI0/XI0_59/d_11_ XI11_0/XI0/XI0_59/d__11_ DECAP_INV_G11
XG14886 XI11_0/XI0/XI0_59/d_10_ XI11_0/XI0/XI0_59/d__10_ DECAP_INV_G11
XG14887 XI11_0/XI0/XI0_59/d_9_ XI11_0/XI0/XI0_59/d__9_ DECAP_INV_G11
XG14888 XI11_0/XI0/XI0_59/d_8_ XI11_0/XI0/XI0_59/d__8_ DECAP_INV_G11
XG14889 XI11_0/XI0/XI0_59/d_7_ XI11_0/XI0/XI0_59/d__7_ DECAP_INV_G11
XG14890 XI11_0/XI0/XI0_59/d_6_ XI11_0/XI0/XI0_59/d__6_ DECAP_INV_G11
XG14891 XI11_0/XI0/XI0_59/d_5_ XI11_0/XI0/XI0_59/d__5_ DECAP_INV_G11
XG14892 XI11_0/XI0/XI0_59/d_4_ XI11_0/XI0/XI0_59/d__4_ DECAP_INV_G11
XG14893 XI11_0/XI0/XI0_59/d_3_ XI11_0/XI0/XI0_59/d__3_ DECAP_INV_G11
XG14894 XI11_0/XI0/XI0_59/d_2_ XI11_0/XI0/XI0_59/d__2_ DECAP_INV_G11
XG14895 XI11_0/XI0/XI0_59/d_1_ XI11_0/XI0/XI0_59/d__1_ DECAP_INV_G11
XG14896 XI11_0/XI0/XI0_59/d_0_ XI11_0/XI0/XI0_59/d__0_ DECAP_INV_G11
XG14897 XI11_0/XI0/XI0_58/d__15_ XI11_0/XI0/XI0_58/d_15_ DECAP_INV_G11
XG14898 XI11_0/XI0/XI0_58/d__14_ XI11_0/XI0/XI0_58/d_14_ DECAP_INV_G11
XG14899 XI11_0/XI0/XI0_58/d__13_ XI11_0/XI0/XI0_58/d_13_ DECAP_INV_G11
XG14900 XI11_0/XI0/XI0_58/d__12_ XI11_0/XI0/XI0_58/d_12_ DECAP_INV_G11
XG14901 XI11_0/XI0/XI0_58/d__11_ XI11_0/XI0/XI0_58/d_11_ DECAP_INV_G11
XG14902 XI11_0/XI0/XI0_58/d__10_ XI11_0/XI0/XI0_58/d_10_ DECAP_INV_G11
XG14903 XI11_0/XI0/XI0_58/d__9_ XI11_0/XI0/XI0_58/d_9_ DECAP_INV_G11
XG14904 XI11_0/XI0/XI0_58/d__8_ XI11_0/XI0/XI0_58/d_8_ DECAP_INV_G11
XG14905 XI11_0/XI0/XI0_58/d__7_ XI11_0/XI0/XI0_58/d_7_ DECAP_INV_G11
XG14906 XI11_0/XI0/XI0_58/d__6_ XI11_0/XI0/XI0_58/d_6_ DECAP_INV_G11
XG14907 XI11_0/XI0/XI0_58/d__5_ XI11_0/XI0/XI0_58/d_5_ DECAP_INV_G11
XG14908 XI11_0/XI0/XI0_58/d__4_ XI11_0/XI0/XI0_58/d_4_ DECAP_INV_G11
XG14909 XI11_0/XI0/XI0_58/d__3_ XI11_0/XI0/XI0_58/d_3_ DECAP_INV_G11
XG14910 XI11_0/XI0/XI0_58/d__2_ XI11_0/XI0/XI0_58/d_2_ DECAP_INV_G11
XG14911 XI11_0/XI0/XI0_58/d__1_ XI11_0/XI0/XI0_58/d_1_ DECAP_INV_G11
XG14912 XI11_0/XI0/XI0_58/d__0_ XI11_0/XI0/XI0_58/d_0_ DECAP_INV_G11
XG14913 XI11_0/XI0/XI0_58/d_15_ XI11_0/XI0/XI0_58/d__15_ DECAP_INV_G11
XG14914 XI11_0/XI0/XI0_58/d_14_ XI11_0/XI0/XI0_58/d__14_ DECAP_INV_G11
XG14915 XI11_0/XI0/XI0_58/d_13_ XI11_0/XI0/XI0_58/d__13_ DECAP_INV_G11
XG14916 XI11_0/XI0/XI0_58/d_12_ XI11_0/XI0/XI0_58/d__12_ DECAP_INV_G11
XG14917 XI11_0/XI0/XI0_58/d_11_ XI11_0/XI0/XI0_58/d__11_ DECAP_INV_G11
XG14918 XI11_0/XI0/XI0_58/d_10_ XI11_0/XI0/XI0_58/d__10_ DECAP_INV_G11
XG14919 XI11_0/XI0/XI0_58/d_9_ XI11_0/XI0/XI0_58/d__9_ DECAP_INV_G11
XG14920 XI11_0/XI0/XI0_58/d_8_ XI11_0/XI0/XI0_58/d__8_ DECAP_INV_G11
XG14921 XI11_0/XI0/XI0_58/d_7_ XI11_0/XI0/XI0_58/d__7_ DECAP_INV_G11
XG14922 XI11_0/XI0/XI0_58/d_6_ XI11_0/XI0/XI0_58/d__6_ DECAP_INV_G11
XG14923 XI11_0/XI0/XI0_58/d_5_ XI11_0/XI0/XI0_58/d__5_ DECAP_INV_G11
XG14924 XI11_0/XI0/XI0_58/d_4_ XI11_0/XI0/XI0_58/d__4_ DECAP_INV_G11
XG14925 XI11_0/XI0/XI0_58/d_3_ XI11_0/XI0/XI0_58/d__3_ DECAP_INV_G11
XG14926 XI11_0/XI0/XI0_58/d_2_ XI11_0/XI0/XI0_58/d__2_ DECAP_INV_G11
XG14927 XI11_0/XI0/XI0_58/d_1_ XI11_0/XI0/XI0_58/d__1_ DECAP_INV_G11
XG14928 XI11_0/XI0/XI0_58/d_0_ XI11_0/XI0/XI0_58/d__0_ DECAP_INV_G11
XG14929 XI11_0/XI0/XI0_57/d__15_ XI11_0/XI0/XI0_57/d_15_ DECAP_INV_G11
XG14930 XI11_0/XI0/XI0_57/d__14_ XI11_0/XI0/XI0_57/d_14_ DECAP_INV_G11
XG14931 XI11_0/XI0/XI0_57/d__13_ XI11_0/XI0/XI0_57/d_13_ DECAP_INV_G11
XG14932 XI11_0/XI0/XI0_57/d__12_ XI11_0/XI0/XI0_57/d_12_ DECAP_INV_G11
XG14933 XI11_0/XI0/XI0_57/d__11_ XI11_0/XI0/XI0_57/d_11_ DECAP_INV_G11
XG14934 XI11_0/XI0/XI0_57/d__10_ XI11_0/XI0/XI0_57/d_10_ DECAP_INV_G11
XG14935 XI11_0/XI0/XI0_57/d__9_ XI11_0/XI0/XI0_57/d_9_ DECAP_INV_G11
XG14936 XI11_0/XI0/XI0_57/d__8_ XI11_0/XI0/XI0_57/d_8_ DECAP_INV_G11
XG14937 XI11_0/XI0/XI0_57/d__7_ XI11_0/XI0/XI0_57/d_7_ DECAP_INV_G11
XG14938 XI11_0/XI0/XI0_57/d__6_ XI11_0/XI0/XI0_57/d_6_ DECAP_INV_G11
XG14939 XI11_0/XI0/XI0_57/d__5_ XI11_0/XI0/XI0_57/d_5_ DECAP_INV_G11
XG14940 XI11_0/XI0/XI0_57/d__4_ XI11_0/XI0/XI0_57/d_4_ DECAP_INV_G11
XG14941 XI11_0/XI0/XI0_57/d__3_ XI11_0/XI0/XI0_57/d_3_ DECAP_INV_G11
XG14942 XI11_0/XI0/XI0_57/d__2_ XI11_0/XI0/XI0_57/d_2_ DECAP_INV_G11
XG14943 XI11_0/XI0/XI0_57/d__1_ XI11_0/XI0/XI0_57/d_1_ DECAP_INV_G11
XG14944 XI11_0/XI0/XI0_57/d__0_ XI11_0/XI0/XI0_57/d_0_ DECAP_INV_G11
XG14945 XI11_0/XI0/XI0_57/d_15_ XI11_0/XI0/XI0_57/d__15_ DECAP_INV_G11
XG14946 XI11_0/XI0/XI0_57/d_14_ XI11_0/XI0/XI0_57/d__14_ DECAP_INV_G11
XG14947 XI11_0/XI0/XI0_57/d_13_ XI11_0/XI0/XI0_57/d__13_ DECAP_INV_G11
XG14948 XI11_0/XI0/XI0_57/d_12_ XI11_0/XI0/XI0_57/d__12_ DECAP_INV_G11
XG14949 XI11_0/XI0/XI0_57/d_11_ XI11_0/XI0/XI0_57/d__11_ DECAP_INV_G11
XG14950 XI11_0/XI0/XI0_57/d_10_ XI11_0/XI0/XI0_57/d__10_ DECAP_INV_G11
XG14951 XI11_0/XI0/XI0_57/d_9_ XI11_0/XI0/XI0_57/d__9_ DECAP_INV_G11
XG14952 XI11_0/XI0/XI0_57/d_8_ XI11_0/XI0/XI0_57/d__8_ DECAP_INV_G11
XG14953 XI11_0/XI0/XI0_57/d_7_ XI11_0/XI0/XI0_57/d__7_ DECAP_INV_G11
XG14954 XI11_0/XI0/XI0_57/d_6_ XI11_0/XI0/XI0_57/d__6_ DECAP_INV_G11
XG14955 XI11_0/XI0/XI0_57/d_5_ XI11_0/XI0/XI0_57/d__5_ DECAP_INV_G11
XG14956 XI11_0/XI0/XI0_57/d_4_ XI11_0/XI0/XI0_57/d__4_ DECAP_INV_G11
XG14957 XI11_0/XI0/XI0_57/d_3_ XI11_0/XI0/XI0_57/d__3_ DECAP_INV_G11
XG14958 XI11_0/XI0/XI0_57/d_2_ XI11_0/XI0/XI0_57/d__2_ DECAP_INV_G11
XG14959 XI11_0/XI0/XI0_57/d_1_ XI11_0/XI0/XI0_57/d__1_ DECAP_INV_G11
XG14960 XI11_0/XI0/XI0_57/d_0_ XI11_0/XI0/XI0_57/d__0_ DECAP_INV_G11
XG14961 XI11_0/XI0/XI0_56/d__15_ XI11_0/XI0/XI0_56/d_15_ DECAP_INV_G11
XG14962 XI11_0/XI0/XI0_56/d__14_ XI11_0/XI0/XI0_56/d_14_ DECAP_INV_G11
XG14963 XI11_0/XI0/XI0_56/d__13_ XI11_0/XI0/XI0_56/d_13_ DECAP_INV_G11
XG14964 XI11_0/XI0/XI0_56/d__12_ XI11_0/XI0/XI0_56/d_12_ DECAP_INV_G11
XG14965 XI11_0/XI0/XI0_56/d__11_ XI11_0/XI0/XI0_56/d_11_ DECAP_INV_G11
XG14966 XI11_0/XI0/XI0_56/d__10_ XI11_0/XI0/XI0_56/d_10_ DECAP_INV_G11
XG14967 XI11_0/XI0/XI0_56/d__9_ XI11_0/XI0/XI0_56/d_9_ DECAP_INV_G11
XG14968 XI11_0/XI0/XI0_56/d__8_ XI11_0/XI0/XI0_56/d_8_ DECAP_INV_G11
XG14969 XI11_0/XI0/XI0_56/d__7_ XI11_0/XI0/XI0_56/d_7_ DECAP_INV_G11
XG14970 XI11_0/XI0/XI0_56/d__6_ XI11_0/XI0/XI0_56/d_6_ DECAP_INV_G11
XG14971 XI11_0/XI0/XI0_56/d__5_ XI11_0/XI0/XI0_56/d_5_ DECAP_INV_G11
XG14972 XI11_0/XI0/XI0_56/d__4_ XI11_0/XI0/XI0_56/d_4_ DECAP_INV_G11
XG14973 XI11_0/XI0/XI0_56/d__3_ XI11_0/XI0/XI0_56/d_3_ DECAP_INV_G11
XG14974 XI11_0/XI0/XI0_56/d__2_ XI11_0/XI0/XI0_56/d_2_ DECAP_INV_G11
XG14975 XI11_0/XI0/XI0_56/d__1_ XI11_0/XI0/XI0_56/d_1_ DECAP_INV_G11
XG14976 XI11_0/XI0/XI0_56/d__0_ XI11_0/XI0/XI0_56/d_0_ DECAP_INV_G11
XG14977 XI11_0/XI0/XI0_56/d_15_ XI11_0/XI0/XI0_56/d__15_ DECAP_INV_G11
XG14978 XI11_0/XI0/XI0_56/d_14_ XI11_0/XI0/XI0_56/d__14_ DECAP_INV_G11
XG14979 XI11_0/XI0/XI0_56/d_13_ XI11_0/XI0/XI0_56/d__13_ DECAP_INV_G11
XG14980 XI11_0/XI0/XI0_56/d_12_ XI11_0/XI0/XI0_56/d__12_ DECAP_INV_G11
XG14981 XI11_0/XI0/XI0_56/d_11_ XI11_0/XI0/XI0_56/d__11_ DECAP_INV_G11
XG14982 XI11_0/XI0/XI0_56/d_10_ XI11_0/XI0/XI0_56/d__10_ DECAP_INV_G11
XG14983 XI11_0/XI0/XI0_56/d_9_ XI11_0/XI0/XI0_56/d__9_ DECAP_INV_G11
XG14984 XI11_0/XI0/XI0_56/d_8_ XI11_0/XI0/XI0_56/d__8_ DECAP_INV_G11
XG14985 XI11_0/XI0/XI0_56/d_7_ XI11_0/XI0/XI0_56/d__7_ DECAP_INV_G11
XG14986 XI11_0/XI0/XI0_56/d_6_ XI11_0/XI0/XI0_56/d__6_ DECAP_INV_G11
XG14987 XI11_0/XI0/XI0_56/d_5_ XI11_0/XI0/XI0_56/d__5_ DECAP_INV_G11
XG14988 XI11_0/XI0/XI0_56/d_4_ XI11_0/XI0/XI0_56/d__4_ DECAP_INV_G11
XG14989 XI11_0/XI0/XI0_56/d_3_ XI11_0/XI0/XI0_56/d__3_ DECAP_INV_G11
XG14990 XI11_0/XI0/XI0_56/d_2_ XI11_0/XI0/XI0_56/d__2_ DECAP_INV_G11
XG14991 XI11_0/XI0/XI0_56/d_1_ XI11_0/XI0/XI0_56/d__1_ DECAP_INV_G11
XG14992 XI11_0/XI0/XI0_56/d_0_ XI11_0/XI0/XI0_56/d__0_ DECAP_INV_G11
XG14993 XI11_0/XI0/XI0_55/d__15_ XI11_0/XI0/XI0_55/d_15_ DECAP_INV_G11
XG14994 XI11_0/XI0/XI0_55/d__14_ XI11_0/XI0/XI0_55/d_14_ DECAP_INV_G11
XG14995 XI11_0/XI0/XI0_55/d__13_ XI11_0/XI0/XI0_55/d_13_ DECAP_INV_G11
XG14996 XI11_0/XI0/XI0_55/d__12_ XI11_0/XI0/XI0_55/d_12_ DECAP_INV_G11
XG14997 XI11_0/XI0/XI0_55/d__11_ XI11_0/XI0/XI0_55/d_11_ DECAP_INV_G11
XG14998 XI11_0/XI0/XI0_55/d__10_ XI11_0/XI0/XI0_55/d_10_ DECAP_INV_G11
XG14999 XI11_0/XI0/XI0_55/d__9_ XI11_0/XI0/XI0_55/d_9_ DECAP_INV_G11
XG15000 XI11_0/XI0/XI0_55/d__8_ XI11_0/XI0/XI0_55/d_8_ DECAP_INV_G11
XG15001 XI11_0/XI0/XI0_55/d__7_ XI11_0/XI0/XI0_55/d_7_ DECAP_INV_G11
XG15002 XI11_0/XI0/XI0_55/d__6_ XI11_0/XI0/XI0_55/d_6_ DECAP_INV_G11
XG15003 XI11_0/XI0/XI0_55/d__5_ XI11_0/XI0/XI0_55/d_5_ DECAP_INV_G11
XG15004 XI11_0/XI0/XI0_55/d__4_ XI11_0/XI0/XI0_55/d_4_ DECAP_INV_G11
XG15005 XI11_0/XI0/XI0_55/d__3_ XI11_0/XI0/XI0_55/d_3_ DECAP_INV_G11
XG15006 XI11_0/XI0/XI0_55/d__2_ XI11_0/XI0/XI0_55/d_2_ DECAP_INV_G11
XG15007 XI11_0/XI0/XI0_55/d__1_ XI11_0/XI0/XI0_55/d_1_ DECAP_INV_G11
XG15008 XI11_0/XI0/XI0_55/d__0_ XI11_0/XI0/XI0_55/d_0_ DECAP_INV_G11
XG15009 XI11_0/XI0/XI0_55/d_15_ XI11_0/XI0/XI0_55/d__15_ DECAP_INV_G11
XG15010 XI11_0/XI0/XI0_55/d_14_ XI11_0/XI0/XI0_55/d__14_ DECAP_INV_G11
XG15011 XI11_0/XI0/XI0_55/d_13_ XI11_0/XI0/XI0_55/d__13_ DECAP_INV_G11
XG15012 XI11_0/XI0/XI0_55/d_12_ XI11_0/XI0/XI0_55/d__12_ DECAP_INV_G11
XG15013 XI11_0/XI0/XI0_55/d_11_ XI11_0/XI0/XI0_55/d__11_ DECAP_INV_G11
XG15014 XI11_0/XI0/XI0_55/d_10_ XI11_0/XI0/XI0_55/d__10_ DECAP_INV_G11
XG15015 XI11_0/XI0/XI0_55/d_9_ XI11_0/XI0/XI0_55/d__9_ DECAP_INV_G11
XG15016 XI11_0/XI0/XI0_55/d_8_ XI11_0/XI0/XI0_55/d__8_ DECAP_INV_G11
XG15017 XI11_0/XI0/XI0_55/d_7_ XI11_0/XI0/XI0_55/d__7_ DECAP_INV_G11
XG15018 XI11_0/XI0/XI0_55/d_6_ XI11_0/XI0/XI0_55/d__6_ DECAP_INV_G11
XG15019 XI11_0/XI0/XI0_55/d_5_ XI11_0/XI0/XI0_55/d__5_ DECAP_INV_G11
XG15020 XI11_0/XI0/XI0_55/d_4_ XI11_0/XI0/XI0_55/d__4_ DECAP_INV_G11
XG15021 XI11_0/XI0/XI0_55/d_3_ XI11_0/XI0/XI0_55/d__3_ DECAP_INV_G11
XG15022 XI11_0/XI0/XI0_55/d_2_ XI11_0/XI0/XI0_55/d__2_ DECAP_INV_G11
XG15023 XI11_0/XI0/XI0_55/d_1_ XI11_0/XI0/XI0_55/d__1_ DECAP_INV_G11
XG15024 XI11_0/XI0/XI0_55/d_0_ XI11_0/XI0/XI0_55/d__0_ DECAP_INV_G11
XG15025 XI11_0/XI0/XI0_54/d__15_ XI11_0/XI0/XI0_54/d_15_ DECAP_INV_G11
XG15026 XI11_0/XI0/XI0_54/d__14_ XI11_0/XI0/XI0_54/d_14_ DECAP_INV_G11
XG15027 XI11_0/XI0/XI0_54/d__13_ XI11_0/XI0/XI0_54/d_13_ DECAP_INV_G11
XG15028 XI11_0/XI0/XI0_54/d__12_ XI11_0/XI0/XI0_54/d_12_ DECAP_INV_G11
XG15029 XI11_0/XI0/XI0_54/d__11_ XI11_0/XI0/XI0_54/d_11_ DECAP_INV_G11
XG15030 XI11_0/XI0/XI0_54/d__10_ XI11_0/XI0/XI0_54/d_10_ DECAP_INV_G11
XG15031 XI11_0/XI0/XI0_54/d__9_ XI11_0/XI0/XI0_54/d_9_ DECAP_INV_G11
XG15032 XI11_0/XI0/XI0_54/d__8_ XI11_0/XI0/XI0_54/d_8_ DECAP_INV_G11
XG15033 XI11_0/XI0/XI0_54/d__7_ XI11_0/XI0/XI0_54/d_7_ DECAP_INV_G11
XG15034 XI11_0/XI0/XI0_54/d__6_ XI11_0/XI0/XI0_54/d_6_ DECAP_INV_G11
XG15035 XI11_0/XI0/XI0_54/d__5_ XI11_0/XI0/XI0_54/d_5_ DECAP_INV_G11
XG15036 XI11_0/XI0/XI0_54/d__4_ XI11_0/XI0/XI0_54/d_4_ DECAP_INV_G11
XG15037 XI11_0/XI0/XI0_54/d__3_ XI11_0/XI0/XI0_54/d_3_ DECAP_INV_G11
XG15038 XI11_0/XI0/XI0_54/d__2_ XI11_0/XI0/XI0_54/d_2_ DECAP_INV_G11
XG15039 XI11_0/XI0/XI0_54/d__1_ XI11_0/XI0/XI0_54/d_1_ DECAP_INV_G11
XG15040 XI11_0/XI0/XI0_54/d__0_ XI11_0/XI0/XI0_54/d_0_ DECAP_INV_G11
XG15041 XI11_0/XI0/XI0_54/d_15_ XI11_0/XI0/XI0_54/d__15_ DECAP_INV_G11
XG15042 XI11_0/XI0/XI0_54/d_14_ XI11_0/XI0/XI0_54/d__14_ DECAP_INV_G11
XG15043 XI11_0/XI0/XI0_54/d_13_ XI11_0/XI0/XI0_54/d__13_ DECAP_INV_G11
XG15044 XI11_0/XI0/XI0_54/d_12_ XI11_0/XI0/XI0_54/d__12_ DECAP_INV_G11
XG15045 XI11_0/XI0/XI0_54/d_11_ XI11_0/XI0/XI0_54/d__11_ DECAP_INV_G11
XG15046 XI11_0/XI0/XI0_54/d_10_ XI11_0/XI0/XI0_54/d__10_ DECAP_INV_G11
XG15047 XI11_0/XI0/XI0_54/d_9_ XI11_0/XI0/XI0_54/d__9_ DECAP_INV_G11
XG15048 XI11_0/XI0/XI0_54/d_8_ XI11_0/XI0/XI0_54/d__8_ DECAP_INV_G11
XG15049 XI11_0/XI0/XI0_54/d_7_ XI11_0/XI0/XI0_54/d__7_ DECAP_INV_G11
XG15050 XI11_0/XI0/XI0_54/d_6_ XI11_0/XI0/XI0_54/d__6_ DECAP_INV_G11
XG15051 XI11_0/XI0/XI0_54/d_5_ XI11_0/XI0/XI0_54/d__5_ DECAP_INV_G11
XG15052 XI11_0/XI0/XI0_54/d_4_ XI11_0/XI0/XI0_54/d__4_ DECAP_INV_G11
XG15053 XI11_0/XI0/XI0_54/d_3_ XI11_0/XI0/XI0_54/d__3_ DECAP_INV_G11
XG15054 XI11_0/XI0/XI0_54/d_2_ XI11_0/XI0/XI0_54/d__2_ DECAP_INV_G11
XG15055 XI11_0/XI0/XI0_54/d_1_ XI11_0/XI0/XI0_54/d__1_ DECAP_INV_G11
XG15056 XI11_0/XI0/XI0_54/d_0_ XI11_0/XI0/XI0_54/d__0_ DECAP_INV_G11
XG15057 XI11_0/XI0/XI0_53/d__15_ XI11_0/XI0/XI0_53/d_15_ DECAP_INV_G11
XG15058 XI11_0/XI0/XI0_53/d__14_ XI11_0/XI0/XI0_53/d_14_ DECAP_INV_G11
XG15059 XI11_0/XI0/XI0_53/d__13_ XI11_0/XI0/XI0_53/d_13_ DECAP_INV_G11
XG15060 XI11_0/XI0/XI0_53/d__12_ XI11_0/XI0/XI0_53/d_12_ DECAP_INV_G11
XG15061 XI11_0/XI0/XI0_53/d__11_ XI11_0/XI0/XI0_53/d_11_ DECAP_INV_G11
XG15062 XI11_0/XI0/XI0_53/d__10_ XI11_0/XI0/XI0_53/d_10_ DECAP_INV_G11
XG15063 XI11_0/XI0/XI0_53/d__9_ XI11_0/XI0/XI0_53/d_9_ DECAP_INV_G11
XG15064 XI11_0/XI0/XI0_53/d__8_ XI11_0/XI0/XI0_53/d_8_ DECAP_INV_G11
XG15065 XI11_0/XI0/XI0_53/d__7_ XI11_0/XI0/XI0_53/d_7_ DECAP_INV_G11
XG15066 XI11_0/XI0/XI0_53/d__6_ XI11_0/XI0/XI0_53/d_6_ DECAP_INV_G11
XG15067 XI11_0/XI0/XI0_53/d__5_ XI11_0/XI0/XI0_53/d_5_ DECAP_INV_G11
XG15068 XI11_0/XI0/XI0_53/d__4_ XI11_0/XI0/XI0_53/d_4_ DECAP_INV_G11
XG15069 XI11_0/XI0/XI0_53/d__3_ XI11_0/XI0/XI0_53/d_3_ DECAP_INV_G11
XG15070 XI11_0/XI0/XI0_53/d__2_ XI11_0/XI0/XI0_53/d_2_ DECAP_INV_G11
XG15071 XI11_0/XI0/XI0_53/d__1_ XI11_0/XI0/XI0_53/d_1_ DECAP_INV_G11
XG15072 XI11_0/XI0/XI0_53/d__0_ XI11_0/XI0/XI0_53/d_0_ DECAP_INV_G11
XG15073 XI11_0/XI0/XI0_53/d_15_ XI11_0/XI0/XI0_53/d__15_ DECAP_INV_G11
XG15074 XI11_0/XI0/XI0_53/d_14_ XI11_0/XI0/XI0_53/d__14_ DECAP_INV_G11
XG15075 XI11_0/XI0/XI0_53/d_13_ XI11_0/XI0/XI0_53/d__13_ DECAP_INV_G11
XG15076 XI11_0/XI0/XI0_53/d_12_ XI11_0/XI0/XI0_53/d__12_ DECAP_INV_G11
XG15077 XI11_0/XI0/XI0_53/d_11_ XI11_0/XI0/XI0_53/d__11_ DECAP_INV_G11
XG15078 XI11_0/XI0/XI0_53/d_10_ XI11_0/XI0/XI0_53/d__10_ DECAP_INV_G11
XG15079 XI11_0/XI0/XI0_53/d_9_ XI11_0/XI0/XI0_53/d__9_ DECAP_INV_G11
XG15080 XI11_0/XI0/XI0_53/d_8_ XI11_0/XI0/XI0_53/d__8_ DECAP_INV_G11
XG15081 XI11_0/XI0/XI0_53/d_7_ XI11_0/XI0/XI0_53/d__7_ DECAP_INV_G11
XG15082 XI11_0/XI0/XI0_53/d_6_ XI11_0/XI0/XI0_53/d__6_ DECAP_INV_G11
XG15083 XI11_0/XI0/XI0_53/d_5_ XI11_0/XI0/XI0_53/d__5_ DECAP_INV_G11
XG15084 XI11_0/XI0/XI0_53/d_4_ XI11_0/XI0/XI0_53/d__4_ DECAP_INV_G11
XG15085 XI11_0/XI0/XI0_53/d_3_ XI11_0/XI0/XI0_53/d__3_ DECAP_INV_G11
XG15086 XI11_0/XI0/XI0_53/d_2_ XI11_0/XI0/XI0_53/d__2_ DECAP_INV_G11
XG15087 XI11_0/XI0/XI0_53/d_1_ XI11_0/XI0/XI0_53/d__1_ DECAP_INV_G11
XG15088 XI11_0/XI0/XI0_53/d_0_ XI11_0/XI0/XI0_53/d__0_ DECAP_INV_G11
XG15089 XI11_0/XI0/XI0_52/d__15_ XI11_0/XI0/XI0_52/d_15_ DECAP_INV_G11
XG15090 XI11_0/XI0/XI0_52/d__14_ XI11_0/XI0/XI0_52/d_14_ DECAP_INV_G11
XG15091 XI11_0/XI0/XI0_52/d__13_ XI11_0/XI0/XI0_52/d_13_ DECAP_INV_G11
XG15092 XI11_0/XI0/XI0_52/d__12_ XI11_0/XI0/XI0_52/d_12_ DECAP_INV_G11
XG15093 XI11_0/XI0/XI0_52/d__11_ XI11_0/XI0/XI0_52/d_11_ DECAP_INV_G11
XG15094 XI11_0/XI0/XI0_52/d__10_ XI11_0/XI0/XI0_52/d_10_ DECAP_INV_G11
XG15095 XI11_0/XI0/XI0_52/d__9_ XI11_0/XI0/XI0_52/d_9_ DECAP_INV_G11
XG15096 XI11_0/XI0/XI0_52/d__8_ XI11_0/XI0/XI0_52/d_8_ DECAP_INV_G11
XG15097 XI11_0/XI0/XI0_52/d__7_ XI11_0/XI0/XI0_52/d_7_ DECAP_INV_G11
XG15098 XI11_0/XI0/XI0_52/d__6_ XI11_0/XI0/XI0_52/d_6_ DECAP_INV_G11
XG15099 XI11_0/XI0/XI0_52/d__5_ XI11_0/XI0/XI0_52/d_5_ DECAP_INV_G11
XG15100 XI11_0/XI0/XI0_52/d__4_ XI11_0/XI0/XI0_52/d_4_ DECAP_INV_G11
XG15101 XI11_0/XI0/XI0_52/d__3_ XI11_0/XI0/XI0_52/d_3_ DECAP_INV_G11
XG15102 XI11_0/XI0/XI0_52/d__2_ XI11_0/XI0/XI0_52/d_2_ DECAP_INV_G11
XG15103 XI11_0/XI0/XI0_52/d__1_ XI11_0/XI0/XI0_52/d_1_ DECAP_INV_G11
XG15104 XI11_0/XI0/XI0_52/d__0_ XI11_0/XI0/XI0_52/d_0_ DECAP_INV_G11
XG15105 XI11_0/XI0/XI0_52/d_15_ XI11_0/XI0/XI0_52/d__15_ DECAP_INV_G11
XG15106 XI11_0/XI0/XI0_52/d_14_ XI11_0/XI0/XI0_52/d__14_ DECAP_INV_G11
XG15107 XI11_0/XI0/XI0_52/d_13_ XI11_0/XI0/XI0_52/d__13_ DECAP_INV_G11
XG15108 XI11_0/XI0/XI0_52/d_12_ XI11_0/XI0/XI0_52/d__12_ DECAP_INV_G11
XG15109 XI11_0/XI0/XI0_52/d_11_ XI11_0/XI0/XI0_52/d__11_ DECAP_INV_G11
XG15110 XI11_0/XI0/XI0_52/d_10_ XI11_0/XI0/XI0_52/d__10_ DECAP_INV_G11
XG15111 XI11_0/XI0/XI0_52/d_9_ XI11_0/XI0/XI0_52/d__9_ DECAP_INV_G11
XG15112 XI11_0/XI0/XI0_52/d_8_ XI11_0/XI0/XI0_52/d__8_ DECAP_INV_G11
XG15113 XI11_0/XI0/XI0_52/d_7_ XI11_0/XI0/XI0_52/d__7_ DECAP_INV_G11
XG15114 XI11_0/XI0/XI0_52/d_6_ XI11_0/XI0/XI0_52/d__6_ DECAP_INV_G11
XG15115 XI11_0/XI0/XI0_52/d_5_ XI11_0/XI0/XI0_52/d__5_ DECAP_INV_G11
XG15116 XI11_0/XI0/XI0_52/d_4_ XI11_0/XI0/XI0_52/d__4_ DECAP_INV_G11
XG15117 XI11_0/XI0/XI0_52/d_3_ XI11_0/XI0/XI0_52/d__3_ DECAP_INV_G11
XG15118 XI11_0/XI0/XI0_52/d_2_ XI11_0/XI0/XI0_52/d__2_ DECAP_INV_G11
XG15119 XI11_0/XI0/XI0_52/d_1_ XI11_0/XI0/XI0_52/d__1_ DECAP_INV_G11
XG15120 XI11_0/XI0/XI0_52/d_0_ XI11_0/XI0/XI0_52/d__0_ DECAP_INV_G11
XG15121 XI11_0/XI0/XI0_51/d__15_ XI11_0/XI0/XI0_51/d_15_ DECAP_INV_G11
XG15122 XI11_0/XI0/XI0_51/d__14_ XI11_0/XI0/XI0_51/d_14_ DECAP_INV_G11
XG15123 XI11_0/XI0/XI0_51/d__13_ XI11_0/XI0/XI0_51/d_13_ DECAP_INV_G11
XG15124 XI11_0/XI0/XI0_51/d__12_ XI11_0/XI0/XI0_51/d_12_ DECAP_INV_G11
XG15125 XI11_0/XI0/XI0_51/d__11_ XI11_0/XI0/XI0_51/d_11_ DECAP_INV_G11
XG15126 XI11_0/XI0/XI0_51/d__10_ XI11_0/XI0/XI0_51/d_10_ DECAP_INV_G11
XG15127 XI11_0/XI0/XI0_51/d__9_ XI11_0/XI0/XI0_51/d_9_ DECAP_INV_G11
XG15128 XI11_0/XI0/XI0_51/d__8_ XI11_0/XI0/XI0_51/d_8_ DECAP_INV_G11
XG15129 XI11_0/XI0/XI0_51/d__7_ XI11_0/XI0/XI0_51/d_7_ DECAP_INV_G11
XG15130 XI11_0/XI0/XI0_51/d__6_ XI11_0/XI0/XI0_51/d_6_ DECAP_INV_G11
XG15131 XI11_0/XI0/XI0_51/d__5_ XI11_0/XI0/XI0_51/d_5_ DECAP_INV_G11
XG15132 XI11_0/XI0/XI0_51/d__4_ XI11_0/XI0/XI0_51/d_4_ DECAP_INV_G11
XG15133 XI11_0/XI0/XI0_51/d__3_ XI11_0/XI0/XI0_51/d_3_ DECAP_INV_G11
XG15134 XI11_0/XI0/XI0_51/d__2_ XI11_0/XI0/XI0_51/d_2_ DECAP_INV_G11
XG15135 XI11_0/XI0/XI0_51/d__1_ XI11_0/XI0/XI0_51/d_1_ DECAP_INV_G11
XG15136 XI11_0/XI0/XI0_51/d__0_ XI11_0/XI0/XI0_51/d_0_ DECAP_INV_G11
XG15137 XI11_0/XI0/XI0_51/d_15_ XI11_0/XI0/XI0_51/d__15_ DECAP_INV_G11
XG15138 XI11_0/XI0/XI0_51/d_14_ XI11_0/XI0/XI0_51/d__14_ DECAP_INV_G11
XG15139 XI11_0/XI0/XI0_51/d_13_ XI11_0/XI0/XI0_51/d__13_ DECAP_INV_G11
XG15140 XI11_0/XI0/XI0_51/d_12_ XI11_0/XI0/XI0_51/d__12_ DECAP_INV_G11
XG15141 XI11_0/XI0/XI0_51/d_11_ XI11_0/XI0/XI0_51/d__11_ DECAP_INV_G11
XG15142 XI11_0/XI0/XI0_51/d_10_ XI11_0/XI0/XI0_51/d__10_ DECAP_INV_G11
XG15143 XI11_0/XI0/XI0_51/d_9_ XI11_0/XI0/XI0_51/d__9_ DECAP_INV_G11
XG15144 XI11_0/XI0/XI0_51/d_8_ XI11_0/XI0/XI0_51/d__8_ DECAP_INV_G11
XG15145 XI11_0/XI0/XI0_51/d_7_ XI11_0/XI0/XI0_51/d__7_ DECAP_INV_G11
XG15146 XI11_0/XI0/XI0_51/d_6_ XI11_0/XI0/XI0_51/d__6_ DECAP_INV_G11
XG15147 XI11_0/XI0/XI0_51/d_5_ XI11_0/XI0/XI0_51/d__5_ DECAP_INV_G11
XG15148 XI11_0/XI0/XI0_51/d_4_ XI11_0/XI0/XI0_51/d__4_ DECAP_INV_G11
XG15149 XI11_0/XI0/XI0_51/d_3_ XI11_0/XI0/XI0_51/d__3_ DECAP_INV_G11
XG15150 XI11_0/XI0/XI0_51/d_2_ XI11_0/XI0/XI0_51/d__2_ DECAP_INV_G11
XG15151 XI11_0/XI0/XI0_51/d_1_ XI11_0/XI0/XI0_51/d__1_ DECAP_INV_G11
XG15152 XI11_0/XI0/XI0_51/d_0_ XI11_0/XI0/XI0_51/d__0_ DECAP_INV_G11
XG15153 XI11_0/XI0/XI0_50/d__15_ XI11_0/XI0/XI0_50/d_15_ DECAP_INV_G11
XG15154 XI11_0/XI0/XI0_50/d__14_ XI11_0/XI0/XI0_50/d_14_ DECAP_INV_G11
XG15155 XI11_0/XI0/XI0_50/d__13_ XI11_0/XI0/XI0_50/d_13_ DECAP_INV_G11
XG15156 XI11_0/XI0/XI0_50/d__12_ XI11_0/XI0/XI0_50/d_12_ DECAP_INV_G11
XG15157 XI11_0/XI0/XI0_50/d__11_ XI11_0/XI0/XI0_50/d_11_ DECAP_INV_G11
XG15158 XI11_0/XI0/XI0_50/d__10_ XI11_0/XI0/XI0_50/d_10_ DECAP_INV_G11
XG15159 XI11_0/XI0/XI0_50/d__9_ XI11_0/XI0/XI0_50/d_9_ DECAP_INV_G11
XG15160 XI11_0/XI0/XI0_50/d__8_ XI11_0/XI0/XI0_50/d_8_ DECAP_INV_G11
XG15161 XI11_0/XI0/XI0_50/d__7_ XI11_0/XI0/XI0_50/d_7_ DECAP_INV_G11
XG15162 XI11_0/XI0/XI0_50/d__6_ XI11_0/XI0/XI0_50/d_6_ DECAP_INV_G11
XG15163 XI11_0/XI0/XI0_50/d__5_ XI11_0/XI0/XI0_50/d_5_ DECAP_INV_G11
XG15164 XI11_0/XI0/XI0_50/d__4_ XI11_0/XI0/XI0_50/d_4_ DECAP_INV_G11
XG15165 XI11_0/XI0/XI0_50/d__3_ XI11_0/XI0/XI0_50/d_3_ DECAP_INV_G11
XG15166 XI11_0/XI0/XI0_50/d__2_ XI11_0/XI0/XI0_50/d_2_ DECAP_INV_G11
XG15167 XI11_0/XI0/XI0_50/d__1_ XI11_0/XI0/XI0_50/d_1_ DECAP_INV_G11
XG15168 XI11_0/XI0/XI0_50/d__0_ XI11_0/XI0/XI0_50/d_0_ DECAP_INV_G11
XG15169 XI11_0/XI0/XI0_50/d_15_ XI11_0/XI0/XI0_50/d__15_ DECAP_INV_G11
XG15170 XI11_0/XI0/XI0_50/d_14_ XI11_0/XI0/XI0_50/d__14_ DECAP_INV_G11
XG15171 XI11_0/XI0/XI0_50/d_13_ XI11_0/XI0/XI0_50/d__13_ DECAP_INV_G11
XG15172 XI11_0/XI0/XI0_50/d_12_ XI11_0/XI0/XI0_50/d__12_ DECAP_INV_G11
XG15173 XI11_0/XI0/XI0_50/d_11_ XI11_0/XI0/XI0_50/d__11_ DECAP_INV_G11
XG15174 XI11_0/XI0/XI0_50/d_10_ XI11_0/XI0/XI0_50/d__10_ DECAP_INV_G11
XG15175 XI11_0/XI0/XI0_50/d_9_ XI11_0/XI0/XI0_50/d__9_ DECAP_INV_G11
XG15176 XI11_0/XI0/XI0_50/d_8_ XI11_0/XI0/XI0_50/d__8_ DECAP_INV_G11
XG15177 XI11_0/XI0/XI0_50/d_7_ XI11_0/XI0/XI0_50/d__7_ DECAP_INV_G11
XG15178 XI11_0/XI0/XI0_50/d_6_ XI11_0/XI0/XI0_50/d__6_ DECAP_INV_G11
XG15179 XI11_0/XI0/XI0_50/d_5_ XI11_0/XI0/XI0_50/d__5_ DECAP_INV_G11
XG15180 XI11_0/XI0/XI0_50/d_4_ XI11_0/XI0/XI0_50/d__4_ DECAP_INV_G11
XG15181 XI11_0/XI0/XI0_50/d_3_ XI11_0/XI0/XI0_50/d__3_ DECAP_INV_G11
XG15182 XI11_0/XI0/XI0_50/d_2_ XI11_0/XI0/XI0_50/d__2_ DECAP_INV_G11
XG15183 XI11_0/XI0/XI0_50/d_1_ XI11_0/XI0/XI0_50/d__1_ DECAP_INV_G11
XG15184 XI11_0/XI0/XI0_50/d_0_ XI11_0/XI0/XI0_50/d__0_ DECAP_INV_G11
XG15185 XI11_0/XI0/XI0_49/d__15_ XI11_0/XI0/XI0_49/d_15_ DECAP_INV_G11
XG15186 XI11_0/XI0/XI0_49/d__14_ XI11_0/XI0/XI0_49/d_14_ DECAP_INV_G11
XG15187 XI11_0/XI0/XI0_49/d__13_ XI11_0/XI0/XI0_49/d_13_ DECAP_INV_G11
XG15188 XI11_0/XI0/XI0_49/d__12_ XI11_0/XI0/XI0_49/d_12_ DECAP_INV_G11
XG15189 XI11_0/XI0/XI0_49/d__11_ XI11_0/XI0/XI0_49/d_11_ DECAP_INV_G11
XG15190 XI11_0/XI0/XI0_49/d__10_ XI11_0/XI0/XI0_49/d_10_ DECAP_INV_G11
XG15191 XI11_0/XI0/XI0_49/d__9_ XI11_0/XI0/XI0_49/d_9_ DECAP_INV_G11
XG15192 XI11_0/XI0/XI0_49/d__8_ XI11_0/XI0/XI0_49/d_8_ DECAP_INV_G11
XG15193 XI11_0/XI0/XI0_49/d__7_ XI11_0/XI0/XI0_49/d_7_ DECAP_INV_G11
XG15194 XI11_0/XI0/XI0_49/d__6_ XI11_0/XI0/XI0_49/d_6_ DECAP_INV_G11
XG15195 XI11_0/XI0/XI0_49/d__5_ XI11_0/XI0/XI0_49/d_5_ DECAP_INV_G11
XG15196 XI11_0/XI0/XI0_49/d__4_ XI11_0/XI0/XI0_49/d_4_ DECAP_INV_G11
XG15197 XI11_0/XI0/XI0_49/d__3_ XI11_0/XI0/XI0_49/d_3_ DECAP_INV_G11
XG15198 XI11_0/XI0/XI0_49/d__2_ XI11_0/XI0/XI0_49/d_2_ DECAP_INV_G11
XG15199 XI11_0/XI0/XI0_49/d__1_ XI11_0/XI0/XI0_49/d_1_ DECAP_INV_G11
XG15200 XI11_0/XI0/XI0_49/d__0_ XI11_0/XI0/XI0_49/d_0_ DECAP_INV_G11
XG15201 XI11_0/XI0/XI0_49/d_15_ XI11_0/XI0/XI0_49/d__15_ DECAP_INV_G11
XG15202 XI11_0/XI0/XI0_49/d_14_ XI11_0/XI0/XI0_49/d__14_ DECAP_INV_G11
XG15203 XI11_0/XI0/XI0_49/d_13_ XI11_0/XI0/XI0_49/d__13_ DECAP_INV_G11
XG15204 XI11_0/XI0/XI0_49/d_12_ XI11_0/XI0/XI0_49/d__12_ DECAP_INV_G11
XG15205 XI11_0/XI0/XI0_49/d_11_ XI11_0/XI0/XI0_49/d__11_ DECAP_INV_G11
XG15206 XI11_0/XI0/XI0_49/d_10_ XI11_0/XI0/XI0_49/d__10_ DECAP_INV_G11
XG15207 XI11_0/XI0/XI0_49/d_9_ XI11_0/XI0/XI0_49/d__9_ DECAP_INV_G11
XG15208 XI11_0/XI0/XI0_49/d_8_ XI11_0/XI0/XI0_49/d__8_ DECAP_INV_G11
XG15209 XI11_0/XI0/XI0_49/d_7_ XI11_0/XI0/XI0_49/d__7_ DECAP_INV_G11
XG15210 XI11_0/XI0/XI0_49/d_6_ XI11_0/XI0/XI0_49/d__6_ DECAP_INV_G11
XG15211 XI11_0/XI0/XI0_49/d_5_ XI11_0/XI0/XI0_49/d__5_ DECAP_INV_G11
XG15212 XI11_0/XI0/XI0_49/d_4_ XI11_0/XI0/XI0_49/d__4_ DECAP_INV_G11
XG15213 XI11_0/XI0/XI0_49/d_3_ XI11_0/XI0/XI0_49/d__3_ DECAP_INV_G11
XG15214 XI11_0/XI0/XI0_49/d_2_ XI11_0/XI0/XI0_49/d__2_ DECAP_INV_G11
XG15215 XI11_0/XI0/XI0_49/d_1_ XI11_0/XI0/XI0_49/d__1_ DECAP_INV_G11
XG15216 XI11_0/XI0/XI0_49/d_0_ XI11_0/XI0/XI0_49/d__0_ DECAP_INV_G11
XG15217 XI11_0/XI0/XI0_48/d__15_ XI11_0/XI0/XI0_48/d_15_ DECAP_INV_G11
XG15218 XI11_0/XI0/XI0_48/d__14_ XI11_0/XI0/XI0_48/d_14_ DECAP_INV_G11
XG15219 XI11_0/XI0/XI0_48/d__13_ XI11_0/XI0/XI0_48/d_13_ DECAP_INV_G11
XG15220 XI11_0/XI0/XI0_48/d__12_ XI11_0/XI0/XI0_48/d_12_ DECAP_INV_G11
XG15221 XI11_0/XI0/XI0_48/d__11_ XI11_0/XI0/XI0_48/d_11_ DECAP_INV_G11
XG15222 XI11_0/XI0/XI0_48/d__10_ XI11_0/XI0/XI0_48/d_10_ DECAP_INV_G11
XG15223 XI11_0/XI0/XI0_48/d__9_ XI11_0/XI0/XI0_48/d_9_ DECAP_INV_G11
XG15224 XI11_0/XI0/XI0_48/d__8_ XI11_0/XI0/XI0_48/d_8_ DECAP_INV_G11
XG15225 XI11_0/XI0/XI0_48/d__7_ XI11_0/XI0/XI0_48/d_7_ DECAP_INV_G11
XG15226 XI11_0/XI0/XI0_48/d__6_ XI11_0/XI0/XI0_48/d_6_ DECAP_INV_G11
XG15227 XI11_0/XI0/XI0_48/d__5_ XI11_0/XI0/XI0_48/d_5_ DECAP_INV_G11
XG15228 XI11_0/XI0/XI0_48/d__4_ XI11_0/XI0/XI0_48/d_4_ DECAP_INV_G11
XG15229 XI11_0/XI0/XI0_48/d__3_ XI11_0/XI0/XI0_48/d_3_ DECAP_INV_G11
XG15230 XI11_0/XI0/XI0_48/d__2_ XI11_0/XI0/XI0_48/d_2_ DECAP_INV_G11
XG15231 XI11_0/XI0/XI0_48/d__1_ XI11_0/XI0/XI0_48/d_1_ DECAP_INV_G11
XG15232 XI11_0/XI0/XI0_48/d__0_ XI11_0/XI0/XI0_48/d_0_ DECAP_INV_G11
XG15233 XI11_0/XI0/XI0_48/d_15_ XI11_0/XI0/XI0_48/d__15_ DECAP_INV_G11
XG15234 XI11_0/XI0/XI0_48/d_14_ XI11_0/XI0/XI0_48/d__14_ DECAP_INV_G11
XG15235 XI11_0/XI0/XI0_48/d_13_ XI11_0/XI0/XI0_48/d__13_ DECAP_INV_G11
XG15236 XI11_0/XI0/XI0_48/d_12_ XI11_0/XI0/XI0_48/d__12_ DECAP_INV_G11
XG15237 XI11_0/XI0/XI0_48/d_11_ XI11_0/XI0/XI0_48/d__11_ DECAP_INV_G11
XG15238 XI11_0/XI0/XI0_48/d_10_ XI11_0/XI0/XI0_48/d__10_ DECAP_INV_G11
XG15239 XI11_0/XI0/XI0_48/d_9_ XI11_0/XI0/XI0_48/d__9_ DECAP_INV_G11
XG15240 XI11_0/XI0/XI0_48/d_8_ XI11_0/XI0/XI0_48/d__8_ DECAP_INV_G11
XG15241 XI11_0/XI0/XI0_48/d_7_ XI11_0/XI0/XI0_48/d__7_ DECAP_INV_G11
XG15242 XI11_0/XI0/XI0_48/d_6_ XI11_0/XI0/XI0_48/d__6_ DECAP_INV_G11
XG15243 XI11_0/XI0/XI0_48/d_5_ XI11_0/XI0/XI0_48/d__5_ DECAP_INV_G11
XG15244 XI11_0/XI0/XI0_48/d_4_ XI11_0/XI0/XI0_48/d__4_ DECAP_INV_G11
XG15245 XI11_0/XI0/XI0_48/d_3_ XI11_0/XI0/XI0_48/d__3_ DECAP_INV_G11
XG15246 XI11_0/XI0/XI0_48/d_2_ XI11_0/XI0/XI0_48/d__2_ DECAP_INV_G11
XG15247 XI11_0/XI0/XI0_48/d_1_ XI11_0/XI0/XI0_48/d__1_ DECAP_INV_G11
XG15248 XI11_0/XI0/XI0_48/d_0_ XI11_0/XI0/XI0_48/d__0_ DECAP_INV_G11
XG15249 XI11_0/XI0/XI0_47/d__15_ XI11_0/XI0/XI0_47/d_15_ DECAP_INV_G11
XG15250 XI11_0/XI0/XI0_47/d__14_ XI11_0/XI0/XI0_47/d_14_ DECAP_INV_G11
XG15251 XI11_0/XI0/XI0_47/d__13_ XI11_0/XI0/XI0_47/d_13_ DECAP_INV_G11
XG15252 XI11_0/XI0/XI0_47/d__12_ XI11_0/XI0/XI0_47/d_12_ DECAP_INV_G11
XG15253 XI11_0/XI0/XI0_47/d__11_ XI11_0/XI0/XI0_47/d_11_ DECAP_INV_G11
XG15254 XI11_0/XI0/XI0_47/d__10_ XI11_0/XI0/XI0_47/d_10_ DECAP_INV_G11
XG15255 XI11_0/XI0/XI0_47/d__9_ XI11_0/XI0/XI0_47/d_9_ DECAP_INV_G11
XG15256 XI11_0/XI0/XI0_47/d__8_ XI11_0/XI0/XI0_47/d_8_ DECAP_INV_G11
XG15257 XI11_0/XI0/XI0_47/d__7_ XI11_0/XI0/XI0_47/d_7_ DECAP_INV_G11
XG15258 XI11_0/XI0/XI0_47/d__6_ XI11_0/XI0/XI0_47/d_6_ DECAP_INV_G11
XG15259 XI11_0/XI0/XI0_47/d__5_ XI11_0/XI0/XI0_47/d_5_ DECAP_INV_G11
XG15260 XI11_0/XI0/XI0_47/d__4_ XI11_0/XI0/XI0_47/d_4_ DECAP_INV_G11
XG15261 XI11_0/XI0/XI0_47/d__3_ XI11_0/XI0/XI0_47/d_3_ DECAP_INV_G11
XG15262 XI11_0/XI0/XI0_47/d__2_ XI11_0/XI0/XI0_47/d_2_ DECAP_INV_G11
XG15263 XI11_0/XI0/XI0_47/d__1_ XI11_0/XI0/XI0_47/d_1_ DECAP_INV_G11
XG15264 XI11_0/XI0/XI0_47/d__0_ XI11_0/XI0/XI0_47/d_0_ DECAP_INV_G11
XG15265 XI11_0/XI0/XI0_47/d_15_ XI11_0/XI0/XI0_47/d__15_ DECAP_INV_G11
XG15266 XI11_0/XI0/XI0_47/d_14_ XI11_0/XI0/XI0_47/d__14_ DECAP_INV_G11
XG15267 XI11_0/XI0/XI0_47/d_13_ XI11_0/XI0/XI0_47/d__13_ DECAP_INV_G11
XG15268 XI11_0/XI0/XI0_47/d_12_ XI11_0/XI0/XI0_47/d__12_ DECAP_INV_G11
XG15269 XI11_0/XI0/XI0_47/d_11_ XI11_0/XI0/XI0_47/d__11_ DECAP_INV_G11
XG15270 XI11_0/XI0/XI0_47/d_10_ XI11_0/XI0/XI0_47/d__10_ DECAP_INV_G11
XG15271 XI11_0/XI0/XI0_47/d_9_ XI11_0/XI0/XI0_47/d__9_ DECAP_INV_G11
XG15272 XI11_0/XI0/XI0_47/d_8_ XI11_0/XI0/XI0_47/d__8_ DECAP_INV_G11
XG15273 XI11_0/XI0/XI0_47/d_7_ XI11_0/XI0/XI0_47/d__7_ DECAP_INV_G11
XG15274 XI11_0/XI0/XI0_47/d_6_ XI11_0/XI0/XI0_47/d__6_ DECAP_INV_G11
XG15275 XI11_0/XI0/XI0_47/d_5_ XI11_0/XI0/XI0_47/d__5_ DECAP_INV_G11
XG15276 XI11_0/XI0/XI0_47/d_4_ XI11_0/XI0/XI0_47/d__4_ DECAP_INV_G11
XG15277 XI11_0/XI0/XI0_47/d_3_ XI11_0/XI0/XI0_47/d__3_ DECAP_INV_G11
XG15278 XI11_0/XI0/XI0_47/d_2_ XI11_0/XI0/XI0_47/d__2_ DECAP_INV_G11
XG15279 XI11_0/XI0/XI0_47/d_1_ XI11_0/XI0/XI0_47/d__1_ DECAP_INV_G11
XG15280 XI11_0/XI0/XI0_47/d_0_ XI11_0/XI0/XI0_47/d__0_ DECAP_INV_G11
XG15281 XI11_0/XI0/XI0_46/d__15_ XI11_0/XI0/XI0_46/d_15_ DECAP_INV_G11
XG15282 XI11_0/XI0/XI0_46/d__14_ XI11_0/XI0/XI0_46/d_14_ DECAP_INV_G11
XG15283 XI11_0/XI0/XI0_46/d__13_ XI11_0/XI0/XI0_46/d_13_ DECAP_INV_G11
XG15284 XI11_0/XI0/XI0_46/d__12_ XI11_0/XI0/XI0_46/d_12_ DECAP_INV_G11
XG15285 XI11_0/XI0/XI0_46/d__11_ XI11_0/XI0/XI0_46/d_11_ DECAP_INV_G11
XG15286 XI11_0/XI0/XI0_46/d__10_ XI11_0/XI0/XI0_46/d_10_ DECAP_INV_G11
XG15287 XI11_0/XI0/XI0_46/d__9_ XI11_0/XI0/XI0_46/d_9_ DECAP_INV_G11
XG15288 XI11_0/XI0/XI0_46/d__8_ XI11_0/XI0/XI0_46/d_8_ DECAP_INV_G11
XG15289 XI11_0/XI0/XI0_46/d__7_ XI11_0/XI0/XI0_46/d_7_ DECAP_INV_G11
XG15290 XI11_0/XI0/XI0_46/d__6_ XI11_0/XI0/XI0_46/d_6_ DECAP_INV_G11
XG15291 XI11_0/XI0/XI0_46/d__5_ XI11_0/XI0/XI0_46/d_5_ DECAP_INV_G11
XG15292 XI11_0/XI0/XI0_46/d__4_ XI11_0/XI0/XI0_46/d_4_ DECAP_INV_G11
XG15293 XI11_0/XI0/XI0_46/d__3_ XI11_0/XI0/XI0_46/d_3_ DECAP_INV_G11
XG15294 XI11_0/XI0/XI0_46/d__2_ XI11_0/XI0/XI0_46/d_2_ DECAP_INV_G11
XG15295 XI11_0/XI0/XI0_46/d__1_ XI11_0/XI0/XI0_46/d_1_ DECAP_INV_G11
XG15296 XI11_0/XI0/XI0_46/d__0_ XI11_0/XI0/XI0_46/d_0_ DECAP_INV_G11
XG15297 XI11_0/XI0/XI0_46/d_15_ XI11_0/XI0/XI0_46/d__15_ DECAP_INV_G11
XG15298 XI11_0/XI0/XI0_46/d_14_ XI11_0/XI0/XI0_46/d__14_ DECAP_INV_G11
XG15299 XI11_0/XI0/XI0_46/d_13_ XI11_0/XI0/XI0_46/d__13_ DECAP_INV_G11
XG15300 XI11_0/XI0/XI0_46/d_12_ XI11_0/XI0/XI0_46/d__12_ DECAP_INV_G11
XG15301 XI11_0/XI0/XI0_46/d_11_ XI11_0/XI0/XI0_46/d__11_ DECAP_INV_G11
XG15302 XI11_0/XI0/XI0_46/d_10_ XI11_0/XI0/XI0_46/d__10_ DECAP_INV_G11
XG15303 XI11_0/XI0/XI0_46/d_9_ XI11_0/XI0/XI0_46/d__9_ DECAP_INV_G11
XG15304 XI11_0/XI0/XI0_46/d_8_ XI11_0/XI0/XI0_46/d__8_ DECAP_INV_G11
XG15305 XI11_0/XI0/XI0_46/d_7_ XI11_0/XI0/XI0_46/d__7_ DECAP_INV_G11
XG15306 XI11_0/XI0/XI0_46/d_6_ XI11_0/XI0/XI0_46/d__6_ DECAP_INV_G11
XG15307 XI11_0/XI0/XI0_46/d_5_ XI11_0/XI0/XI0_46/d__5_ DECAP_INV_G11
XG15308 XI11_0/XI0/XI0_46/d_4_ XI11_0/XI0/XI0_46/d__4_ DECAP_INV_G11
XG15309 XI11_0/XI0/XI0_46/d_3_ XI11_0/XI0/XI0_46/d__3_ DECAP_INV_G11
XG15310 XI11_0/XI0/XI0_46/d_2_ XI11_0/XI0/XI0_46/d__2_ DECAP_INV_G11
XG15311 XI11_0/XI0/XI0_46/d_1_ XI11_0/XI0/XI0_46/d__1_ DECAP_INV_G11
XG15312 XI11_0/XI0/XI0_46/d_0_ XI11_0/XI0/XI0_46/d__0_ DECAP_INV_G11
XG15313 XI11_0/XI0/XI0_45/d__15_ XI11_0/XI0/XI0_45/d_15_ DECAP_INV_G11
XG15314 XI11_0/XI0/XI0_45/d__14_ XI11_0/XI0/XI0_45/d_14_ DECAP_INV_G11
XG15315 XI11_0/XI0/XI0_45/d__13_ XI11_0/XI0/XI0_45/d_13_ DECAP_INV_G11
XG15316 XI11_0/XI0/XI0_45/d__12_ XI11_0/XI0/XI0_45/d_12_ DECAP_INV_G11
XG15317 XI11_0/XI0/XI0_45/d__11_ XI11_0/XI0/XI0_45/d_11_ DECAP_INV_G11
XG15318 XI11_0/XI0/XI0_45/d__10_ XI11_0/XI0/XI0_45/d_10_ DECAP_INV_G11
XG15319 XI11_0/XI0/XI0_45/d__9_ XI11_0/XI0/XI0_45/d_9_ DECAP_INV_G11
XG15320 XI11_0/XI0/XI0_45/d__8_ XI11_0/XI0/XI0_45/d_8_ DECAP_INV_G11
XG15321 XI11_0/XI0/XI0_45/d__7_ XI11_0/XI0/XI0_45/d_7_ DECAP_INV_G11
XG15322 XI11_0/XI0/XI0_45/d__6_ XI11_0/XI0/XI0_45/d_6_ DECAP_INV_G11
XG15323 XI11_0/XI0/XI0_45/d__5_ XI11_0/XI0/XI0_45/d_5_ DECAP_INV_G11
XG15324 XI11_0/XI0/XI0_45/d__4_ XI11_0/XI0/XI0_45/d_4_ DECAP_INV_G11
XG15325 XI11_0/XI0/XI0_45/d__3_ XI11_0/XI0/XI0_45/d_3_ DECAP_INV_G11
XG15326 XI11_0/XI0/XI0_45/d__2_ XI11_0/XI0/XI0_45/d_2_ DECAP_INV_G11
XG15327 XI11_0/XI0/XI0_45/d__1_ XI11_0/XI0/XI0_45/d_1_ DECAP_INV_G11
XG15328 XI11_0/XI0/XI0_45/d__0_ XI11_0/XI0/XI0_45/d_0_ DECAP_INV_G11
XG15329 XI11_0/XI0/XI0_45/d_15_ XI11_0/XI0/XI0_45/d__15_ DECAP_INV_G11
XG15330 XI11_0/XI0/XI0_45/d_14_ XI11_0/XI0/XI0_45/d__14_ DECAP_INV_G11
XG15331 XI11_0/XI0/XI0_45/d_13_ XI11_0/XI0/XI0_45/d__13_ DECAP_INV_G11
XG15332 XI11_0/XI0/XI0_45/d_12_ XI11_0/XI0/XI0_45/d__12_ DECAP_INV_G11
XG15333 XI11_0/XI0/XI0_45/d_11_ XI11_0/XI0/XI0_45/d__11_ DECAP_INV_G11
XG15334 XI11_0/XI0/XI0_45/d_10_ XI11_0/XI0/XI0_45/d__10_ DECAP_INV_G11
XG15335 XI11_0/XI0/XI0_45/d_9_ XI11_0/XI0/XI0_45/d__9_ DECAP_INV_G11
XG15336 XI11_0/XI0/XI0_45/d_8_ XI11_0/XI0/XI0_45/d__8_ DECAP_INV_G11
XG15337 XI11_0/XI0/XI0_45/d_7_ XI11_0/XI0/XI0_45/d__7_ DECAP_INV_G11
XG15338 XI11_0/XI0/XI0_45/d_6_ XI11_0/XI0/XI0_45/d__6_ DECAP_INV_G11
XG15339 XI11_0/XI0/XI0_45/d_5_ XI11_0/XI0/XI0_45/d__5_ DECAP_INV_G11
XG15340 XI11_0/XI0/XI0_45/d_4_ XI11_0/XI0/XI0_45/d__4_ DECAP_INV_G11
XG15341 XI11_0/XI0/XI0_45/d_3_ XI11_0/XI0/XI0_45/d__3_ DECAP_INV_G11
XG15342 XI11_0/XI0/XI0_45/d_2_ XI11_0/XI0/XI0_45/d__2_ DECAP_INV_G11
XG15343 XI11_0/XI0/XI0_45/d_1_ XI11_0/XI0/XI0_45/d__1_ DECAP_INV_G11
XG15344 XI11_0/XI0/XI0_45/d_0_ XI11_0/XI0/XI0_45/d__0_ DECAP_INV_G11
XG15345 XI11_0/XI0/XI0_44/d__15_ XI11_0/XI0/XI0_44/d_15_ DECAP_INV_G11
XG15346 XI11_0/XI0/XI0_44/d__14_ XI11_0/XI0/XI0_44/d_14_ DECAP_INV_G11
XG15347 XI11_0/XI0/XI0_44/d__13_ XI11_0/XI0/XI0_44/d_13_ DECAP_INV_G11
XG15348 XI11_0/XI0/XI0_44/d__12_ XI11_0/XI0/XI0_44/d_12_ DECAP_INV_G11
XG15349 XI11_0/XI0/XI0_44/d__11_ XI11_0/XI0/XI0_44/d_11_ DECAP_INV_G11
XG15350 XI11_0/XI0/XI0_44/d__10_ XI11_0/XI0/XI0_44/d_10_ DECAP_INV_G11
XG15351 XI11_0/XI0/XI0_44/d__9_ XI11_0/XI0/XI0_44/d_9_ DECAP_INV_G11
XG15352 XI11_0/XI0/XI0_44/d__8_ XI11_0/XI0/XI0_44/d_8_ DECAP_INV_G11
XG15353 XI11_0/XI0/XI0_44/d__7_ XI11_0/XI0/XI0_44/d_7_ DECAP_INV_G11
XG15354 XI11_0/XI0/XI0_44/d__6_ XI11_0/XI0/XI0_44/d_6_ DECAP_INV_G11
XG15355 XI11_0/XI0/XI0_44/d__5_ XI11_0/XI0/XI0_44/d_5_ DECAP_INV_G11
XG15356 XI11_0/XI0/XI0_44/d__4_ XI11_0/XI0/XI0_44/d_4_ DECAP_INV_G11
XG15357 XI11_0/XI0/XI0_44/d__3_ XI11_0/XI0/XI0_44/d_3_ DECAP_INV_G11
XG15358 XI11_0/XI0/XI0_44/d__2_ XI11_0/XI0/XI0_44/d_2_ DECAP_INV_G11
XG15359 XI11_0/XI0/XI0_44/d__1_ XI11_0/XI0/XI0_44/d_1_ DECAP_INV_G11
XG15360 XI11_0/XI0/XI0_44/d__0_ XI11_0/XI0/XI0_44/d_0_ DECAP_INV_G11
XG15361 XI11_0/XI0/XI0_44/d_15_ XI11_0/XI0/XI0_44/d__15_ DECAP_INV_G11
XG15362 XI11_0/XI0/XI0_44/d_14_ XI11_0/XI0/XI0_44/d__14_ DECAP_INV_G11
XG15363 XI11_0/XI0/XI0_44/d_13_ XI11_0/XI0/XI0_44/d__13_ DECAP_INV_G11
XG15364 XI11_0/XI0/XI0_44/d_12_ XI11_0/XI0/XI0_44/d__12_ DECAP_INV_G11
XG15365 XI11_0/XI0/XI0_44/d_11_ XI11_0/XI0/XI0_44/d__11_ DECAP_INV_G11
XG15366 XI11_0/XI0/XI0_44/d_10_ XI11_0/XI0/XI0_44/d__10_ DECAP_INV_G11
XG15367 XI11_0/XI0/XI0_44/d_9_ XI11_0/XI0/XI0_44/d__9_ DECAP_INV_G11
XG15368 XI11_0/XI0/XI0_44/d_8_ XI11_0/XI0/XI0_44/d__8_ DECAP_INV_G11
XG15369 XI11_0/XI0/XI0_44/d_7_ XI11_0/XI0/XI0_44/d__7_ DECAP_INV_G11
XG15370 XI11_0/XI0/XI0_44/d_6_ XI11_0/XI0/XI0_44/d__6_ DECAP_INV_G11
XG15371 XI11_0/XI0/XI0_44/d_5_ XI11_0/XI0/XI0_44/d__5_ DECAP_INV_G11
XG15372 XI11_0/XI0/XI0_44/d_4_ XI11_0/XI0/XI0_44/d__4_ DECAP_INV_G11
XG15373 XI11_0/XI0/XI0_44/d_3_ XI11_0/XI0/XI0_44/d__3_ DECAP_INV_G11
XG15374 XI11_0/XI0/XI0_44/d_2_ XI11_0/XI0/XI0_44/d__2_ DECAP_INV_G11
XG15375 XI11_0/XI0/XI0_44/d_1_ XI11_0/XI0/XI0_44/d__1_ DECAP_INV_G11
XG15376 XI11_0/XI0/XI0_44/d_0_ XI11_0/XI0/XI0_44/d__0_ DECAP_INV_G11
XG15377 XI11_0/XI0/XI0_43/d__15_ XI11_0/XI0/XI0_43/d_15_ DECAP_INV_G11
XG15378 XI11_0/XI0/XI0_43/d__14_ XI11_0/XI0/XI0_43/d_14_ DECAP_INV_G11
XG15379 XI11_0/XI0/XI0_43/d__13_ XI11_0/XI0/XI0_43/d_13_ DECAP_INV_G11
XG15380 XI11_0/XI0/XI0_43/d__12_ XI11_0/XI0/XI0_43/d_12_ DECAP_INV_G11
XG15381 XI11_0/XI0/XI0_43/d__11_ XI11_0/XI0/XI0_43/d_11_ DECAP_INV_G11
XG15382 XI11_0/XI0/XI0_43/d__10_ XI11_0/XI0/XI0_43/d_10_ DECAP_INV_G11
XG15383 XI11_0/XI0/XI0_43/d__9_ XI11_0/XI0/XI0_43/d_9_ DECAP_INV_G11
XG15384 XI11_0/XI0/XI0_43/d__8_ XI11_0/XI0/XI0_43/d_8_ DECAP_INV_G11
XG15385 XI11_0/XI0/XI0_43/d__7_ XI11_0/XI0/XI0_43/d_7_ DECAP_INV_G11
XG15386 XI11_0/XI0/XI0_43/d__6_ XI11_0/XI0/XI0_43/d_6_ DECAP_INV_G11
XG15387 XI11_0/XI0/XI0_43/d__5_ XI11_0/XI0/XI0_43/d_5_ DECAP_INV_G11
XG15388 XI11_0/XI0/XI0_43/d__4_ XI11_0/XI0/XI0_43/d_4_ DECAP_INV_G11
XG15389 XI11_0/XI0/XI0_43/d__3_ XI11_0/XI0/XI0_43/d_3_ DECAP_INV_G11
XG15390 XI11_0/XI0/XI0_43/d__2_ XI11_0/XI0/XI0_43/d_2_ DECAP_INV_G11
XG15391 XI11_0/XI0/XI0_43/d__1_ XI11_0/XI0/XI0_43/d_1_ DECAP_INV_G11
XG15392 XI11_0/XI0/XI0_43/d__0_ XI11_0/XI0/XI0_43/d_0_ DECAP_INV_G11
XG15393 XI11_0/XI0/XI0_43/d_15_ XI11_0/XI0/XI0_43/d__15_ DECAP_INV_G11
XG15394 XI11_0/XI0/XI0_43/d_14_ XI11_0/XI0/XI0_43/d__14_ DECAP_INV_G11
XG15395 XI11_0/XI0/XI0_43/d_13_ XI11_0/XI0/XI0_43/d__13_ DECAP_INV_G11
XG15396 XI11_0/XI0/XI0_43/d_12_ XI11_0/XI0/XI0_43/d__12_ DECAP_INV_G11
XG15397 XI11_0/XI0/XI0_43/d_11_ XI11_0/XI0/XI0_43/d__11_ DECAP_INV_G11
XG15398 XI11_0/XI0/XI0_43/d_10_ XI11_0/XI0/XI0_43/d__10_ DECAP_INV_G11
XG15399 XI11_0/XI0/XI0_43/d_9_ XI11_0/XI0/XI0_43/d__9_ DECAP_INV_G11
XG15400 XI11_0/XI0/XI0_43/d_8_ XI11_0/XI0/XI0_43/d__8_ DECAP_INV_G11
XG15401 XI11_0/XI0/XI0_43/d_7_ XI11_0/XI0/XI0_43/d__7_ DECAP_INV_G11
XG15402 XI11_0/XI0/XI0_43/d_6_ XI11_0/XI0/XI0_43/d__6_ DECAP_INV_G11
XG15403 XI11_0/XI0/XI0_43/d_5_ XI11_0/XI0/XI0_43/d__5_ DECAP_INV_G11
XG15404 XI11_0/XI0/XI0_43/d_4_ XI11_0/XI0/XI0_43/d__4_ DECAP_INV_G11
XG15405 XI11_0/XI0/XI0_43/d_3_ XI11_0/XI0/XI0_43/d__3_ DECAP_INV_G11
XG15406 XI11_0/XI0/XI0_43/d_2_ XI11_0/XI0/XI0_43/d__2_ DECAP_INV_G11
XG15407 XI11_0/XI0/XI0_43/d_1_ XI11_0/XI0/XI0_43/d__1_ DECAP_INV_G11
XG15408 XI11_0/XI0/XI0_43/d_0_ XI11_0/XI0/XI0_43/d__0_ DECAP_INV_G11
XG15409 XI11_0/XI0/XI0_42/d__15_ XI11_0/XI0/XI0_42/d_15_ DECAP_INV_G11
XG15410 XI11_0/XI0/XI0_42/d__14_ XI11_0/XI0/XI0_42/d_14_ DECAP_INV_G11
XG15411 XI11_0/XI0/XI0_42/d__13_ XI11_0/XI0/XI0_42/d_13_ DECAP_INV_G11
XG15412 XI11_0/XI0/XI0_42/d__12_ XI11_0/XI0/XI0_42/d_12_ DECAP_INV_G11
XG15413 XI11_0/XI0/XI0_42/d__11_ XI11_0/XI0/XI0_42/d_11_ DECAP_INV_G11
XG15414 XI11_0/XI0/XI0_42/d__10_ XI11_0/XI0/XI0_42/d_10_ DECAP_INV_G11
XG15415 XI11_0/XI0/XI0_42/d__9_ XI11_0/XI0/XI0_42/d_9_ DECAP_INV_G11
XG15416 XI11_0/XI0/XI0_42/d__8_ XI11_0/XI0/XI0_42/d_8_ DECAP_INV_G11
XG15417 XI11_0/XI0/XI0_42/d__7_ XI11_0/XI0/XI0_42/d_7_ DECAP_INV_G11
XG15418 XI11_0/XI0/XI0_42/d__6_ XI11_0/XI0/XI0_42/d_6_ DECAP_INV_G11
XG15419 XI11_0/XI0/XI0_42/d__5_ XI11_0/XI0/XI0_42/d_5_ DECAP_INV_G11
XG15420 XI11_0/XI0/XI0_42/d__4_ XI11_0/XI0/XI0_42/d_4_ DECAP_INV_G11
XG15421 XI11_0/XI0/XI0_42/d__3_ XI11_0/XI0/XI0_42/d_3_ DECAP_INV_G11
XG15422 XI11_0/XI0/XI0_42/d__2_ XI11_0/XI0/XI0_42/d_2_ DECAP_INV_G11
XG15423 XI11_0/XI0/XI0_42/d__1_ XI11_0/XI0/XI0_42/d_1_ DECAP_INV_G11
XG15424 XI11_0/XI0/XI0_42/d__0_ XI11_0/XI0/XI0_42/d_0_ DECAP_INV_G11
XG15425 XI11_0/XI0/XI0_42/d_15_ XI11_0/XI0/XI0_42/d__15_ DECAP_INV_G11
XG15426 XI11_0/XI0/XI0_42/d_14_ XI11_0/XI0/XI0_42/d__14_ DECAP_INV_G11
XG15427 XI11_0/XI0/XI0_42/d_13_ XI11_0/XI0/XI0_42/d__13_ DECAP_INV_G11
XG15428 XI11_0/XI0/XI0_42/d_12_ XI11_0/XI0/XI0_42/d__12_ DECAP_INV_G11
XG15429 XI11_0/XI0/XI0_42/d_11_ XI11_0/XI0/XI0_42/d__11_ DECAP_INV_G11
XG15430 XI11_0/XI0/XI0_42/d_10_ XI11_0/XI0/XI0_42/d__10_ DECAP_INV_G11
XG15431 XI11_0/XI0/XI0_42/d_9_ XI11_0/XI0/XI0_42/d__9_ DECAP_INV_G11
XG15432 XI11_0/XI0/XI0_42/d_8_ XI11_0/XI0/XI0_42/d__8_ DECAP_INV_G11
XG15433 XI11_0/XI0/XI0_42/d_7_ XI11_0/XI0/XI0_42/d__7_ DECAP_INV_G11
XG15434 XI11_0/XI0/XI0_42/d_6_ XI11_0/XI0/XI0_42/d__6_ DECAP_INV_G11
XG15435 XI11_0/XI0/XI0_42/d_5_ XI11_0/XI0/XI0_42/d__5_ DECAP_INV_G11
XG15436 XI11_0/XI0/XI0_42/d_4_ XI11_0/XI0/XI0_42/d__4_ DECAP_INV_G11
XG15437 XI11_0/XI0/XI0_42/d_3_ XI11_0/XI0/XI0_42/d__3_ DECAP_INV_G11
XG15438 XI11_0/XI0/XI0_42/d_2_ XI11_0/XI0/XI0_42/d__2_ DECAP_INV_G11
XG15439 XI11_0/XI0/XI0_42/d_1_ XI11_0/XI0/XI0_42/d__1_ DECAP_INV_G11
XG15440 XI11_0/XI0/XI0_42/d_0_ XI11_0/XI0/XI0_42/d__0_ DECAP_INV_G11
XG15441 XI11_0/XI0/XI0_41/d__15_ XI11_0/XI0/XI0_41/d_15_ DECAP_INV_G11
XG15442 XI11_0/XI0/XI0_41/d__14_ XI11_0/XI0/XI0_41/d_14_ DECAP_INV_G11
XG15443 XI11_0/XI0/XI0_41/d__13_ XI11_0/XI0/XI0_41/d_13_ DECAP_INV_G11
XG15444 XI11_0/XI0/XI0_41/d__12_ XI11_0/XI0/XI0_41/d_12_ DECAP_INV_G11
XG15445 XI11_0/XI0/XI0_41/d__11_ XI11_0/XI0/XI0_41/d_11_ DECAP_INV_G11
XG15446 XI11_0/XI0/XI0_41/d__10_ XI11_0/XI0/XI0_41/d_10_ DECAP_INV_G11
XG15447 XI11_0/XI0/XI0_41/d__9_ XI11_0/XI0/XI0_41/d_9_ DECAP_INV_G11
XG15448 XI11_0/XI0/XI0_41/d__8_ XI11_0/XI0/XI0_41/d_8_ DECAP_INV_G11
XG15449 XI11_0/XI0/XI0_41/d__7_ XI11_0/XI0/XI0_41/d_7_ DECAP_INV_G11
XG15450 XI11_0/XI0/XI0_41/d__6_ XI11_0/XI0/XI0_41/d_6_ DECAP_INV_G11
XG15451 XI11_0/XI0/XI0_41/d__5_ XI11_0/XI0/XI0_41/d_5_ DECAP_INV_G11
XG15452 XI11_0/XI0/XI0_41/d__4_ XI11_0/XI0/XI0_41/d_4_ DECAP_INV_G11
XG15453 XI11_0/XI0/XI0_41/d__3_ XI11_0/XI0/XI0_41/d_3_ DECAP_INV_G11
XG15454 XI11_0/XI0/XI0_41/d__2_ XI11_0/XI0/XI0_41/d_2_ DECAP_INV_G11
XG15455 XI11_0/XI0/XI0_41/d__1_ XI11_0/XI0/XI0_41/d_1_ DECAP_INV_G11
XG15456 XI11_0/XI0/XI0_41/d__0_ XI11_0/XI0/XI0_41/d_0_ DECAP_INV_G11
XG15457 XI11_0/XI0/XI0_41/d_15_ XI11_0/XI0/XI0_41/d__15_ DECAP_INV_G11
XG15458 XI11_0/XI0/XI0_41/d_14_ XI11_0/XI0/XI0_41/d__14_ DECAP_INV_G11
XG15459 XI11_0/XI0/XI0_41/d_13_ XI11_0/XI0/XI0_41/d__13_ DECAP_INV_G11
XG15460 XI11_0/XI0/XI0_41/d_12_ XI11_0/XI0/XI0_41/d__12_ DECAP_INV_G11
XG15461 XI11_0/XI0/XI0_41/d_11_ XI11_0/XI0/XI0_41/d__11_ DECAP_INV_G11
XG15462 XI11_0/XI0/XI0_41/d_10_ XI11_0/XI0/XI0_41/d__10_ DECAP_INV_G11
XG15463 XI11_0/XI0/XI0_41/d_9_ XI11_0/XI0/XI0_41/d__9_ DECAP_INV_G11
XG15464 XI11_0/XI0/XI0_41/d_8_ XI11_0/XI0/XI0_41/d__8_ DECAP_INV_G11
XG15465 XI11_0/XI0/XI0_41/d_7_ XI11_0/XI0/XI0_41/d__7_ DECAP_INV_G11
XG15466 XI11_0/XI0/XI0_41/d_6_ XI11_0/XI0/XI0_41/d__6_ DECAP_INV_G11
XG15467 XI11_0/XI0/XI0_41/d_5_ XI11_0/XI0/XI0_41/d__5_ DECAP_INV_G11
XG15468 XI11_0/XI0/XI0_41/d_4_ XI11_0/XI0/XI0_41/d__4_ DECAP_INV_G11
XG15469 XI11_0/XI0/XI0_41/d_3_ XI11_0/XI0/XI0_41/d__3_ DECAP_INV_G11
XG15470 XI11_0/XI0/XI0_41/d_2_ XI11_0/XI0/XI0_41/d__2_ DECAP_INV_G11
XG15471 XI11_0/XI0/XI0_41/d_1_ XI11_0/XI0/XI0_41/d__1_ DECAP_INV_G11
XG15472 XI11_0/XI0/XI0_41/d_0_ XI11_0/XI0/XI0_41/d__0_ DECAP_INV_G11
XG15473 XI11_0/XI0/XI0_40/d__15_ XI11_0/XI0/XI0_40/d_15_ DECAP_INV_G11
XG15474 XI11_0/XI0/XI0_40/d__14_ XI11_0/XI0/XI0_40/d_14_ DECAP_INV_G11
XG15475 XI11_0/XI0/XI0_40/d__13_ XI11_0/XI0/XI0_40/d_13_ DECAP_INV_G11
XG15476 XI11_0/XI0/XI0_40/d__12_ XI11_0/XI0/XI0_40/d_12_ DECAP_INV_G11
XG15477 XI11_0/XI0/XI0_40/d__11_ XI11_0/XI0/XI0_40/d_11_ DECAP_INV_G11
XG15478 XI11_0/XI0/XI0_40/d__10_ XI11_0/XI0/XI0_40/d_10_ DECAP_INV_G11
XG15479 XI11_0/XI0/XI0_40/d__9_ XI11_0/XI0/XI0_40/d_9_ DECAP_INV_G11
XG15480 XI11_0/XI0/XI0_40/d__8_ XI11_0/XI0/XI0_40/d_8_ DECAP_INV_G11
XG15481 XI11_0/XI0/XI0_40/d__7_ XI11_0/XI0/XI0_40/d_7_ DECAP_INV_G11
XG15482 XI11_0/XI0/XI0_40/d__6_ XI11_0/XI0/XI0_40/d_6_ DECAP_INV_G11
XG15483 XI11_0/XI0/XI0_40/d__5_ XI11_0/XI0/XI0_40/d_5_ DECAP_INV_G11
XG15484 XI11_0/XI0/XI0_40/d__4_ XI11_0/XI0/XI0_40/d_4_ DECAP_INV_G11
XG15485 XI11_0/XI0/XI0_40/d__3_ XI11_0/XI0/XI0_40/d_3_ DECAP_INV_G11
XG15486 XI11_0/XI0/XI0_40/d__2_ XI11_0/XI0/XI0_40/d_2_ DECAP_INV_G11
XG15487 XI11_0/XI0/XI0_40/d__1_ XI11_0/XI0/XI0_40/d_1_ DECAP_INV_G11
XG15488 XI11_0/XI0/XI0_40/d__0_ XI11_0/XI0/XI0_40/d_0_ DECAP_INV_G11
XG15489 XI11_0/XI0/XI0_40/d_15_ XI11_0/XI0/XI0_40/d__15_ DECAP_INV_G11
XG15490 XI11_0/XI0/XI0_40/d_14_ XI11_0/XI0/XI0_40/d__14_ DECAP_INV_G11
XG15491 XI11_0/XI0/XI0_40/d_13_ XI11_0/XI0/XI0_40/d__13_ DECAP_INV_G11
XG15492 XI11_0/XI0/XI0_40/d_12_ XI11_0/XI0/XI0_40/d__12_ DECAP_INV_G11
XG15493 XI11_0/XI0/XI0_40/d_11_ XI11_0/XI0/XI0_40/d__11_ DECAP_INV_G11
XG15494 XI11_0/XI0/XI0_40/d_10_ XI11_0/XI0/XI0_40/d__10_ DECAP_INV_G11
XG15495 XI11_0/XI0/XI0_40/d_9_ XI11_0/XI0/XI0_40/d__9_ DECAP_INV_G11
XG15496 XI11_0/XI0/XI0_40/d_8_ XI11_0/XI0/XI0_40/d__8_ DECAP_INV_G11
XG15497 XI11_0/XI0/XI0_40/d_7_ XI11_0/XI0/XI0_40/d__7_ DECAP_INV_G11
XG15498 XI11_0/XI0/XI0_40/d_6_ XI11_0/XI0/XI0_40/d__6_ DECAP_INV_G11
XG15499 XI11_0/XI0/XI0_40/d_5_ XI11_0/XI0/XI0_40/d__5_ DECAP_INV_G11
XG15500 XI11_0/XI0/XI0_40/d_4_ XI11_0/XI0/XI0_40/d__4_ DECAP_INV_G11
XG15501 XI11_0/XI0/XI0_40/d_3_ XI11_0/XI0/XI0_40/d__3_ DECAP_INV_G11
XG15502 XI11_0/XI0/XI0_40/d_2_ XI11_0/XI0/XI0_40/d__2_ DECAP_INV_G11
XG15503 XI11_0/XI0/XI0_40/d_1_ XI11_0/XI0/XI0_40/d__1_ DECAP_INV_G11
XG15504 XI11_0/XI0/XI0_40/d_0_ XI11_0/XI0/XI0_40/d__0_ DECAP_INV_G11
XG15505 XI11_0/XI0/XI0_39/d__15_ XI11_0/XI0/XI0_39/d_15_ DECAP_INV_G11
XG15506 XI11_0/XI0/XI0_39/d__14_ XI11_0/XI0/XI0_39/d_14_ DECAP_INV_G11
XG15507 XI11_0/XI0/XI0_39/d__13_ XI11_0/XI0/XI0_39/d_13_ DECAP_INV_G11
XG15508 XI11_0/XI0/XI0_39/d__12_ XI11_0/XI0/XI0_39/d_12_ DECAP_INV_G11
XG15509 XI11_0/XI0/XI0_39/d__11_ XI11_0/XI0/XI0_39/d_11_ DECAP_INV_G11
XG15510 XI11_0/XI0/XI0_39/d__10_ XI11_0/XI0/XI0_39/d_10_ DECAP_INV_G11
XG15511 XI11_0/XI0/XI0_39/d__9_ XI11_0/XI0/XI0_39/d_9_ DECAP_INV_G11
XG15512 XI11_0/XI0/XI0_39/d__8_ XI11_0/XI0/XI0_39/d_8_ DECAP_INV_G11
XG15513 XI11_0/XI0/XI0_39/d__7_ XI11_0/XI0/XI0_39/d_7_ DECAP_INV_G11
XG15514 XI11_0/XI0/XI0_39/d__6_ XI11_0/XI0/XI0_39/d_6_ DECAP_INV_G11
XG15515 XI11_0/XI0/XI0_39/d__5_ XI11_0/XI0/XI0_39/d_5_ DECAP_INV_G11
XG15516 XI11_0/XI0/XI0_39/d__4_ XI11_0/XI0/XI0_39/d_4_ DECAP_INV_G11
XG15517 XI11_0/XI0/XI0_39/d__3_ XI11_0/XI0/XI0_39/d_3_ DECAP_INV_G11
XG15518 XI11_0/XI0/XI0_39/d__2_ XI11_0/XI0/XI0_39/d_2_ DECAP_INV_G11
XG15519 XI11_0/XI0/XI0_39/d__1_ XI11_0/XI0/XI0_39/d_1_ DECAP_INV_G11
XG15520 XI11_0/XI0/XI0_39/d__0_ XI11_0/XI0/XI0_39/d_0_ DECAP_INV_G11
XG15521 XI11_0/XI0/XI0_39/d_15_ XI11_0/XI0/XI0_39/d__15_ DECAP_INV_G11
XG15522 XI11_0/XI0/XI0_39/d_14_ XI11_0/XI0/XI0_39/d__14_ DECAP_INV_G11
XG15523 XI11_0/XI0/XI0_39/d_13_ XI11_0/XI0/XI0_39/d__13_ DECAP_INV_G11
XG15524 XI11_0/XI0/XI0_39/d_12_ XI11_0/XI0/XI0_39/d__12_ DECAP_INV_G11
XG15525 XI11_0/XI0/XI0_39/d_11_ XI11_0/XI0/XI0_39/d__11_ DECAP_INV_G11
XG15526 XI11_0/XI0/XI0_39/d_10_ XI11_0/XI0/XI0_39/d__10_ DECAP_INV_G11
XG15527 XI11_0/XI0/XI0_39/d_9_ XI11_0/XI0/XI0_39/d__9_ DECAP_INV_G11
XG15528 XI11_0/XI0/XI0_39/d_8_ XI11_0/XI0/XI0_39/d__8_ DECAP_INV_G11
XG15529 XI11_0/XI0/XI0_39/d_7_ XI11_0/XI0/XI0_39/d__7_ DECAP_INV_G11
XG15530 XI11_0/XI0/XI0_39/d_6_ XI11_0/XI0/XI0_39/d__6_ DECAP_INV_G11
XG15531 XI11_0/XI0/XI0_39/d_5_ XI11_0/XI0/XI0_39/d__5_ DECAP_INV_G11
XG15532 XI11_0/XI0/XI0_39/d_4_ XI11_0/XI0/XI0_39/d__4_ DECAP_INV_G11
XG15533 XI11_0/XI0/XI0_39/d_3_ XI11_0/XI0/XI0_39/d__3_ DECAP_INV_G11
XG15534 XI11_0/XI0/XI0_39/d_2_ XI11_0/XI0/XI0_39/d__2_ DECAP_INV_G11
XG15535 XI11_0/XI0/XI0_39/d_1_ XI11_0/XI0/XI0_39/d__1_ DECAP_INV_G11
XG15536 XI11_0/XI0/XI0_39/d_0_ XI11_0/XI0/XI0_39/d__0_ DECAP_INV_G11
XG15537 XI11_0/XI0/XI0_38/d__15_ XI11_0/XI0/XI0_38/d_15_ DECAP_INV_G11
XG15538 XI11_0/XI0/XI0_38/d__14_ XI11_0/XI0/XI0_38/d_14_ DECAP_INV_G11
XG15539 XI11_0/XI0/XI0_38/d__13_ XI11_0/XI0/XI0_38/d_13_ DECAP_INV_G11
XG15540 XI11_0/XI0/XI0_38/d__12_ XI11_0/XI0/XI0_38/d_12_ DECAP_INV_G11
XG15541 XI11_0/XI0/XI0_38/d__11_ XI11_0/XI0/XI0_38/d_11_ DECAP_INV_G11
XG15542 XI11_0/XI0/XI0_38/d__10_ XI11_0/XI0/XI0_38/d_10_ DECAP_INV_G11
XG15543 XI11_0/XI0/XI0_38/d__9_ XI11_0/XI0/XI0_38/d_9_ DECAP_INV_G11
XG15544 XI11_0/XI0/XI0_38/d__8_ XI11_0/XI0/XI0_38/d_8_ DECAP_INV_G11
XG15545 XI11_0/XI0/XI0_38/d__7_ XI11_0/XI0/XI0_38/d_7_ DECAP_INV_G11
XG15546 XI11_0/XI0/XI0_38/d__6_ XI11_0/XI0/XI0_38/d_6_ DECAP_INV_G11
XG15547 XI11_0/XI0/XI0_38/d__5_ XI11_0/XI0/XI0_38/d_5_ DECAP_INV_G11
XG15548 XI11_0/XI0/XI0_38/d__4_ XI11_0/XI0/XI0_38/d_4_ DECAP_INV_G11
XG15549 XI11_0/XI0/XI0_38/d__3_ XI11_0/XI0/XI0_38/d_3_ DECAP_INV_G11
XG15550 XI11_0/XI0/XI0_38/d__2_ XI11_0/XI0/XI0_38/d_2_ DECAP_INV_G11
XG15551 XI11_0/XI0/XI0_38/d__1_ XI11_0/XI0/XI0_38/d_1_ DECAP_INV_G11
XG15552 XI11_0/XI0/XI0_38/d__0_ XI11_0/XI0/XI0_38/d_0_ DECAP_INV_G11
XG15553 XI11_0/XI0/XI0_38/d_15_ XI11_0/XI0/XI0_38/d__15_ DECAP_INV_G11
XG15554 XI11_0/XI0/XI0_38/d_14_ XI11_0/XI0/XI0_38/d__14_ DECAP_INV_G11
XG15555 XI11_0/XI0/XI0_38/d_13_ XI11_0/XI0/XI0_38/d__13_ DECAP_INV_G11
XG15556 XI11_0/XI0/XI0_38/d_12_ XI11_0/XI0/XI0_38/d__12_ DECAP_INV_G11
XG15557 XI11_0/XI0/XI0_38/d_11_ XI11_0/XI0/XI0_38/d__11_ DECAP_INV_G11
XG15558 XI11_0/XI0/XI0_38/d_10_ XI11_0/XI0/XI0_38/d__10_ DECAP_INV_G11
XG15559 XI11_0/XI0/XI0_38/d_9_ XI11_0/XI0/XI0_38/d__9_ DECAP_INV_G11
XG15560 XI11_0/XI0/XI0_38/d_8_ XI11_0/XI0/XI0_38/d__8_ DECAP_INV_G11
XG15561 XI11_0/XI0/XI0_38/d_7_ XI11_0/XI0/XI0_38/d__7_ DECAP_INV_G11
XG15562 XI11_0/XI0/XI0_38/d_6_ XI11_0/XI0/XI0_38/d__6_ DECAP_INV_G11
XG15563 XI11_0/XI0/XI0_38/d_5_ XI11_0/XI0/XI0_38/d__5_ DECAP_INV_G11
XG15564 XI11_0/XI0/XI0_38/d_4_ XI11_0/XI0/XI0_38/d__4_ DECAP_INV_G11
XG15565 XI11_0/XI0/XI0_38/d_3_ XI11_0/XI0/XI0_38/d__3_ DECAP_INV_G11
XG15566 XI11_0/XI0/XI0_38/d_2_ XI11_0/XI0/XI0_38/d__2_ DECAP_INV_G11
XG15567 XI11_0/XI0/XI0_38/d_1_ XI11_0/XI0/XI0_38/d__1_ DECAP_INV_G11
XG15568 XI11_0/XI0/XI0_38/d_0_ XI11_0/XI0/XI0_38/d__0_ DECAP_INV_G11
XG15569 XI11_0/XI0/XI0_37/d__15_ XI11_0/XI0/XI0_37/d_15_ DECAP_INV_G11
XG15570 XI11_0/XI0/XI0_37/d__14_ XI11_0/XI0/XI0_37/d_14_ DECAP_INV_G11
XG15571 XI11_0/XI0/XI0_37/d__13_ XI11_0/XI0/XI0_37/d_13_ DECAP_INV_G11
XG15572 XI11_0/XI0/XI0_37/d__12_ XI11_0/XI0/XI0_37/d_12_ DECAP_INV_G11
XG15573 XI11_0/XI0/XI0_37/d__11_ XI11_0/XI0/XI0_37/d_11_ DECAP_INV_G11
XG15574 XI11_0/XI0/XI0_37/d__10_ XI11_0/XI0/XI0_37/d_10_ DECAP_INV_G11
XG15575 XI11_0/XI0/XI0_37/d__9_ XI11_0/XI0/XI0_37/d_9_ DECAP_INV_G11
XG15576 XI11_0/XI0/XI0_37/d__8_ XI11_0/XI0/XI0_37/d_8_ DECAP_INV_G11
XG15577 XI11_0/XI0/XI0_37/d__7_ XI11_0/XI0/XI0_37/d_7_ DECAP_INV_G11
XG15578 XI11_0/XI0/XI0_37/d__6_ XI11_0/XI0/XI0_37/d_6_ DECAP_INV_G11
XG15579 XI11_0/XI0/XI0_37/d__5_ XI11_0/XI0/XI0_37/d_5_ DECAP_INV_G11
XG15580 XI11_0/XI0/XI0_37/d__4_ XI11_0/XI0/XI0_37/d_4_ DECAP_INV_G11
XG15581 XI11_0/XI0/XI0_37/d__3_ XI11_0/XI0/XI0_37/d_3_ DECAP_INV_G11
XG15582 XI11_0/XI0/XI0_37/d__2_ XI11_0/XI0/XI0_37/d_2_ DECAP_INV_G11
XG15583 XI11_0/XI0/XI0_37/d__1_ XI11_0/XI0/XI0_37/d_1_ DECAP_INV_G11
XG15584 XI11_0/XI0/XI0_37/d__0_ XI11_0/XI0/XI0_37/d_0_ DECAP_INV_G11
XG15585 XI11_0/XI0/XI0_37/d_15_ XI11_0/XI0/XI0_37/d__15_ DECAP_INV_G11
XG15586 XI11_0/XI0/XI0_37/d_14_ XI11_0/XI0/XI0_37/d__14_ DECAP_INV_G11
XG15587 XI11_0/XI0/XI0_37/d_13_ XI11_0/XI0/XI0_37/d__13_ DECAP_INV_G11
XG15588 XI11_0/XI0/XI0_37/d_12_ XI11_0/XI0/XI0_37/d__12_ DECAP_INV_G11
XG15589 XI11_0/XI0/XI0_37/d_11_ XI11_0/XI0/XI0_37/d__11_ DECAP_INV_G11
XG15590 XI11_0/XI0/XI0_37/d_10_ XI11_0/XI0/XI0_37/d__10_ DECAP_INV_G11
XG15591 XI11_0/XI0/XI0_37/d_9_ XI11_0/XI0/XI0_37/d__9_ DECAP_INV_G11
XG15592 XI11_0/XI0/XI0_37/d_8_ XI11_0/XI0/XI0_37/d__8_ DECAP_INV_G11
XG15593 XI11_0/XI0/XI0_37/d_7_ XI11_0/XI0/XI0_37/d__7_ DECAP_INV_G11
XG15594 XI11_0/XI0/XI0_37/d_6_ XI11_0/XI0/XI0_37/d__6_ DECAP_INV_G11
XG15595 XI11_0/XI0/XI0_37/d_5_ XI11_0/XI0/XI0_37/d__5_ DECAP_INV_G11
XG15596 XI11_0/XI0/XI0_37/d_4_ XI11_0/XI0/XI0_37/d__4_ DECAP_INV_G11
XG15597 XI11_0/XI0/XI0_37/d_3_ XI11_0/XI0/XI0_37/d__3_ DECAP_INV_G11
XG15598 XI11_0/XI0/XI0_37/d_2_ XI11_0/XI0/XI0_37/d__2_ DECAP_INV_G11
XG15599 XI11_0/XI0/XI0_37/d_1_ XI11_0/XI0/XI0_37/d__1_ DECAP_INV_G11
XG15600 XI11_0/XI0/XI0_37/d_0_ XI11_0/XI0/XI0_37/d__0_ DECAP_INV_G11
XG15601 XI11_0/XI0/XI0_36/d__15_ XI11_0/XI0/XI0_36/d_15_ DECAP_INV_G11
XG15602 XI11_0/XI0/XI0_36/d__14_ XI11_0/XI0/XI0_36/d_14_ DECAP_INV_G11
XG15603 XI11_0/XI0/XI0_36/d__13_ XI11_0/XI0/XI0_36/d_13_ DECAP_INV_G11
XG15604 XI11_0/XI0/XI0_36/d__12_ XI11_0/XI0/XI0_36/d_12_ DECAP_INV_G11
XG15605 XI11_0/XI0/XI0_36/d__11_ XI11_0/XI0/XI0_36/d_11_ DECAP_INV_G11
XG15606 XI11_0/XI0/XI0_36/d__10_ XI11_0/XI0/XI0_36/d_10_ DECAP_INV_G11
XG15607 XI11_0/XI0/XI0_36/d__9_ XI11_0/XI0/XI0_36/d_9_ DECAP_INV_G11
XG15608 XI11_0/XI0/XI0_36/d__8_ XI11_0/XI0/XI0_36/d_8_ DECAP_INV_G11
XG15609 XI11_0/XI0/XI0_36/d__7_ XI11_0/XI0/XI0_36/d_7_ DECAP_INV_G11
XG15610 XI11_0/XI0/XI0_36/d__6_ XI11_0/XI0/XI0_36/d_6_ DECAP_INV_G11
XG15611 XI11_0/XI0/XI0_36/d__5_ XI11_0/XI0/XI0_36/d_5_ DECAP_INV_G11
XG15612 XI11_0/XI0/XI0_36/d__4_ XI11_0/XI0/XI0_36/d_4_ DECAP_INV_G11
XG15613 XI11_0/XI0/XI0_36/d__3_ XI11_0/XI0/XI0_36/d_3_ DECAP_INV_G11
XG15614 XI11_0/XI0/XI0_36/d__2_ XI11_0/XI0/XI0_36/d_2_ DECAP_INV_G11
XG15615 XI11_0/XI0/XI0_36/d__1_ XI11_0/XI0/XI0_36/d_1_ DECAP_INV_G11
XG15616 XI11_0/XI0/XI0_36/d__0_ XI11_0/XI0/XI0_36/d_0_ DECAP_INV_G11
XG15617 XI11_0/XI0/XI0_36/d_15_ XI11_0/XI0/XI0_36/d__15_ DECAP_INV_G11
XG15618 XI11_0/XI0/XI0_36/d_14_ XI11_0/XI0/XI0_36/d__14_ DECAP_INV_G11
XG15619 XI11_0/XI0/XI0_36/d_13_ XI11_0/XI0/XI0_36/d__13_ DECAP_INV_G11
XG15620 XI11_0/XI0/XI0_36/d_12_ XI11_0/XI0/XI0_36/d__12_ DECAP_INV_G11
XG15621 XI11_0/XI0/XI0_36/d_11_ XI11_0/XI0/XI0_36/d__11_ DECAP_INV_G11
XG15622 XI11_0/XI0/XI0_36/d_10_ XI11_0/XI0/XI0_36/d__10_ DECAP_INV_G11
XG15623 XI11_0/XI0/XI0_36/d_9_ XI11_0/XI0/XI0_36/d__9_ DECAP_INV_G11
XG15624 XI11_0/XI0/XI0_36/d_8_ XI11_0/XI0/XI0_36/d__8_ DECAP_INV_G11
XG15625 XI11_0/XI0/XI0_36/d_7_ XI11_0/XI0/XI0_36/d__7_ DECAP_INV_G11
XG15626 XI11_0/XI0/XI0_36/d_6_ XI11_0/XI0/XI0_36/d__6_ DECAP_INV_G11
XG15627 XI11_0/XI0/XI0_36/d_5_ XI11_0/XI0/XI0_36/d__5_ DECAP_INV_G11
XG15628 XI11_0/XI0/XI0_36/d_4_ XI11_0/XI0/XI0_36/d__4_ DECAP_INV_G11
XG15629 XI11_0/XI0/XI0_36/d_3_ XI11_0/XI0/XI0_36/d__3_ DECAP_INV_G11
XG15630 XI11_0/XI0/XI0_36/d_2_ XI11_0/XI0/XI0_36/d__2_ DECAP_INV_G11
XG15631 XI11_0/XI0/XI0_36/d_1_ XI11_0/XI0/XI0_36/d__1_ DECAP_INV_G11
XG15632 XI11_0/XI0/XI0_36/d_0_ XI11_0/XI0/XI0_36/d__0_ DECAP_INV_G11
XG15633 XI11_0/XI0/XI0_35/d__15_ XI11_0/XI0/XI0_35/d_15_ DECAP_INV_G11
XG15634 XI11_0/XI0/XI0_35/d__14_ XI11_0/XI0/XI0_35/d_14_ DECAP_INV_G11
XG15635 XI11_0/XI0/XI0_35/d__13_ XI11_0/XI0/XI0_35/d_13_ DECAP_INV_G11
XG15636 XI11_0/XI0/XI0_35/d__12_ XI11_0/XI0/XI0_35/d_12_ DECAP_INV_G11
XG15637 XI11_0/XI0/XI0_35/d__11_ XI11_0/XI0/XI0_35/d_11_ DECAP_INV_G11
XG15638 XI11_0/XI0/XI0_35/d__10_ XI11_0/XI0/XI0_35/d_10_ DECAP_INV_G11
XG15639 XI11_0/XI0/XI0_35/d__9_ XI11_0/XI0/XI0_35/d_9_ DECAP_INV_G11
XG15640 XI11_0/XI0/XI0_35/d__8_ XI11_0/XI0/XI0_35/d_8_ DECAP_INV_G11
XG15641 XI11_0/XI0/XI0_35/d__7_ XI11_0/XI0/XI0_35/d_7_ DECAP_INV_G11
XG15642 XI11_0/XI0/XI0_35/d__6_ XI11_0/XI0/XI0_35/d_6_ DECAP_INV_G11
XG15643 XI11_0/XI0/XI0_35/d__5_ XI11_0/XI0/XI0_35/d_5_ DECAP_INV_G11
XG15644 XI11_0/XI0/XI0_35/d__4_ XI11_0/XI0/XI0_35/d_4_ DECAP_INV_G11
XG15645 XI11_0/XI0/XI0_35/d__3_ XI11_0/XI0/XI0_35/d_3_ DECAP_INV_G11
XG15646 XI11_0/XI0/XI0_35/d__2_ XI11_0/XI0/XI0_35/d_2_ DECAP_INV_G11
XG15647 XI11_0/XI0/XI0_35/d__1_ XI11_0/XI0/XI0_35/d_1_ DECAP_INV_G11
XG15648 XI11_0/XI0/XI0_35/d__0_ XI11_0/XI0/XI0_35/d_0_ DECAP_INV_G11
XG15649 XI11_0/XI0/XI0_35/d_15_ XI11_0/XI0/XI0_35/d__15_ DECAP_INV_G11
XG15650 XI11_0/XI0/XI0_35/d_14_ XI11_0/XI0/XI0_35/d__14_ DECAP_INV_G11
XG15651 XI11_0/XI0/XI0_35/d_13_ XI11_0/XI0/XI0_35/d__13_ DECAP_INV_G11
XG15652 XI11_0/XI0/XI0_35/d_12_ XI11_0/XI0/XI0_35/d__12_ DECAP_INV_G11
XG15653 XI11_0/XI0/XI0_35/d_11_ XI11_0/XI0/XI0_35/d__11_ DECAP_INV_G11
XG15654 XI11_0/XI0/XI0_35/d_10_ XI11_0/XI0/XI0_35/d__10_ DECAP_INV_G11
XG15655 XI11_0/XI0/XI0_35/d_9_ XI11_0/XI0/XI0_35/d__9_ DECAP_INV_G11
XG15656 XI11_0/XI0/XI0_35/d_8_ XI11_0/XI0/XI0_35/d__8_ DECAP_INV_G11
XG15657 XI11_0/XI0/XI0_35/d_7_ XI11_0/XI0/XI0_35/d__7_ DECAP_INV_G11
XG15658 XI11_0/XI0/XI0_35/d_6_ XI11_0/XI0/XI0_35/d__6_ DECAP_INV_G11
XG15659 XI11_0/XI0/XI0_35/d_5_ XI11_0/XI0/XI0_35/d__5_ DECAP_INV_G11
XG15660 XI11_0/XI0/XI0_35/d_4_ XI11_0/XI0/XI0_35/d__4_ DECAP_INV_G11
XG15661 XI11_0/XI0/XI0_35/d_3_ XI11_0/XI0/XI0_35/d__3_ DECAP_INV_G11
XG15662 XI11_0/XI0/XI0_35/d_2_ XI11_0/XI0/XI0_35/d__2_ DECAP_INV_G11
XG15663 XI11_0/XI0/XI0_35/d_1_ XI11_0/XI0/XI0_35/d__1_ DECAP_INV_G11
XG15664 XI11_0/XI0/XI0_35/d_0_ XI11_0/XI0/XI0_35/d__0_ DECAP_INV_G11
XG15665 XI11_0/XI0/XI0_34/d__15_ XI11_0/XI0/XI0_34/d_15_ DECAP_INV_G11
XG15666 XI11_0/XI0/XI0_34/d__14_ XI11_0/XI0/XI0_34/d_14_ DECAP_INV_G11
XG15667 XI11_0/XI0/XI0_34/d__13_ XI11_0/XI0/XI0_34/d_13_ DECAP_INV_G11
XG15668 XI11_0/XI0/XI0_34/d__12_ XI11_0/XI0/XI0_34/d_12_ DECAP_INV_G11
XG15669 XI11_0/XI0/XI0_34/d__11_ XI11_0/XI0/XI0_34/d_11_ DECAP_INV_G11
XG15670 XI11_0/XI0/XI0_34/d__10_ XI11_0/XI0/XI0_34/d_10_ DECAP_INV_G11
XG15671 XI11_0/XI0/XI0_34/d__9_ XI11_0/XI0/XI0_34/d_9_ DECAP_INV_G11
XG15672 XI11_0/XI0/XI0_34/d__8_ XI11_0/XI0/XI0_34/d_8_ DECAP_INV_G11
XG15673 XI11_0/XI0/XI0_34/d__7_ XI11_0/XI0/XI0_34/d_7_ DECAP_INV_G11
XG15674 XI11_0/XI0/XI0_34/d__6_ XI11_0/XI0/XI0_34/d_6_ DECAP_INV_G11
XG15675 XI11_0/XI0/XI0_34/d__5_ XI11_0/XI0/XI0_34/d_5_ DECAP_INV_G11
XG15676 XI11_0/XI0/XI0_34/d__4_ XI11_0/XI0/XI0_34/d_4_ DECAP_INV_G11
XG15677 XI11_0/XI0/XI0_34/d__3_ XI11_0/XI0/XI0_34/d_3_ DECAP_INV_G11
XG15678 XI11_0/XI0/XI0_34/d__2_ XI11_0/XI0/XI0_34/d_2_ DECAP_INV_G11
XG15679 XI11_0/XI0/XI0_34/d__1_ XI11_0/XI0/XI0_34/d_1_ DECAP_INV_G11
XG15680 XI11_0/XI0/XI0_34/d__0_ XI11_0/XI0/XI0_34/d_0_ DECAP_INV_G11
XG15681 XI11_0/XI0/XI0_34/d_15_ XI11_0/XI0/XI0_34/d__15_ DECAP_INV_G11
XG15682 XI11_0/XI0/XI0_34/d_14_ XI11_0/XI0/XI0_34/d__14_ DECAP_INV_G11
XG15683 XI11_0/XI0/XI0_34/d_13_ XI11_0/XI0/XI0_34/d__13_ DECAP_INV_G11
XG15684 XI11_0/XI0/XI0_34/d_12_ XI11_0/XI0/XI0_34/d__12_ DECAP_INV_G11
XG15685 XI11_0/XI0/XI0_34/d_11_ XI11_0/XI0/XI0_34/d__11_ DECAP_INV_G11
XG15686 XI11_0/XI0/XI0_34/d_10_ XI11_0/XI0/XI0_34/d__10_ DECAP_INV_G11
XG15687 XI11_0/XI0/XI0_34/d_9_ XI11_0/XI0/XI0_34/d__9_ DECAP_INV_G11
XG15688 XI11_0/XI0/XI0_34/d_8_ XI11_0/XI0/XI0_34/d__8_ DECAP_INV_G11
XG15689 XI11_0/XI0/XI0_34/d_7_ XI11_0/XI0/XI0_34/d__7_ DECAP_INV_G11
XG15690 XI11_0/XI0/XI0_34/d_6_ XI11_0/XI0/XI0_34/d__6_ DECAP_INV_G11
XG15691 XI11_0/XI0/XI0_34/d_5_ XI11_0/XI0/XI0_34/d__5_ DECAP_INV_G11
XG15692 XI11_0/XI0/XI0_34/d_4_ XI11_0/XI0/XI0_34/d__4_ DECAP_INV_G11
XG15693 XI11_0/XI0/XI0_34/d_3_ XI11_0/XI0/XI0_34/d__3_ DECAP_INV_G11
XG15694 XI11_0/XI0/XI0_34/d_2_ XI11_0/XI0/XI0_34/d__2_ DECAP_INV_G11
XG15695 XI11_0/XI0/XI0_34/d_1_ XI11_0/XI0/XI0_34/d__1_ DECAP_INV_G11
XG15696 XI11_0/XI0/XI0_34/d_0_ XI11_0/XI0/XI0_34/d__0_ DECAP_INV_G11
XG15697 XI11_0/XI0/XI0_33/d__15_ XI11_0/XI0/XI0_33/d_15_ DECAP_INV_G11
XG15698 XI11_0/XI0/XI0_33/d__14_ XI11_0/XI0/XI0_33/d_14_ DECAP_INV_G11
XG15699 XI11_0/XI0/XI0_33/d__13_ XI11_0/XI0/XI0_33/d_13_ DECAP_INV_G11
XG15700 XI11_0/XI0/XI0_33/d__12_ XI11_0/XI0/XI0_33/d_12_ DECAP_INV_G11
XG15701 XI11_0/XI0/XI0_33/d__11_ XI11_0/XI0/XI0_33/d_11_ DECAP_INV_G11
XG15702 XI11_0/XI0/XI0_33/d__10_ XI11_0/XI0/XI0_33/d_10_ DECAP_INV_G11
XG15703 XI11_0/XI0/XI0_33/d__9_ XI11_0/XI0/XI0_33/d_9_ DECAP_INV_G11
XG15704 XI11_0/XI0/XI0_33/d__8_ XI11_0/XI0/XI0_33/d_8_ DECAP_INV_G11
XG15705 XI11_0/XI0/XI0_33/d__7_ XI11_0/XI0/XI0_33/d_7_ DECAP_INV_G11
XG15706 XI11_0/XI0/XI0_33/d__6_ XI11_0/XI0/XI0_33/d_6_ DECAP_INV_G11
XG15707 XI11_0/XI0/XI0_33/d__5_ XI11_0/XI0/XI0_33/d_5_ DECAP_INV_G11
XG15708 XI11_0/XI0/XI0_33/d__4_ XI11_0/XI0/XI0_33/d_4_ DECAP_INV_G11
XG15709 XI11_0/XI0/XI0_33/d__3_ XI11_0/XI0/XI0_33/d_3_ DECAP_INV_G11
XG15710 XI11_0/XI0/XI0_33/d__2_ XI11_0/XI0/XI0_33/d_2_ DECAP_INV_G11
XG15711 XI11_0/XI0/XI0_33/d__1_ XI11_0/XI0/XI0_33/d_1_ DECAP_INV_G11
XG15712 XI11_0/XI0/XI0_33/d__0_ XI11_0/XI0/XI0_33/d_0_ DECAP_INV_G11
XG15713 XI11_0/XI0/XI0_33/d_15_ XI11_0/XI0/XI0_33/d__15_ DECAP_INV_G11
XG15714 XI11_0/XI0/XI0_33/d_14_ XI11_0/XI0/XI0_33/d__14_ DECAP_INV_G11
XG15715 XI11_0/XI0/XI0_33/d_13_ XI11_0/XI0/XI0_33/d__13_ DECAP_INV_G11
XG15716 XI11_0/XI0/XI0_33/d_12_ XI11_0/XI0/XI0_33/d__12_ DECAP_INV_G11
XG15717 XI11_0/XI0/XI0_33/d_11_ XI11_0/XI0/XI0_33/d__11_ DECAP_INV_G11
XG15718 XI11_0/XI0/XI0_33/d_10_ XI11_0/XI0/XI0_33/d__10_ DECAP_INV_G11
XG15719 XI11_0/XI0/XI0_33/d_9_ XI11_0/XI0/XI0_33/d__9_ DECAP_INV_G11
XG15720 XI11_0/XI0/XI0_33/d_8_ XI11_0/XI0/XI0_33/d__8_ DECAP_INV_G11
XG15721 XI11_0/XI0/XI0_33/d_7_ XI11_0/XI0/XI0_33/d__7_ DECAP_INV_G11
XG15722 XI11_0/XI0/XI0_33/d_6_ XI11_0/XI0/XI0_33/d__6_ DECAP_INV_G11
XG15723 XI11_0/XI0/XI0_33/d_5_ XI11_0/XI0/XI0_33/d__5_ DECAP_INV_G11
XG15724 XI11_0/XI0/XI0_33/d_4_ XI11_0/XI0/XI0_33/d__4_ DECAP_INV_G11
XG15725 XI11_0/XI0/XI0_33/d_3_ XI11_0/XI0/XI0_33/d__3_ DECAP_INV_G11
XG15726 XI11_0/XI0/XI0_33/d_2_ XI11_0/XI0/XI0_33/d__2_ DECAP_INV_G11
XG15727 XI11_0/XI0/XI0_33/d_1_ XI11_0/XI0/XI0_33/d__1_ DECAP_INV_G11
XG15728 XI11_0/XI0/XI0_33/d_0_ XI11_0/XI0/XI0_33/d__0_ DECAP_INV_G11
XG15729 XI11_0/XI0/XI0_32/d__15_ XI11_0/XI0/XI0_32/d_15_ DECAP_INV_G11
XG15730 XI11_0/XI0/XI0_32/d__14_ XI11_0/XI0/XI0_32/d_14_ DECAP_INV_G11
XG15731 XI11_0/XI0/XI0_32/d__13_ XI11_0/XI0/XI0_32/d_13_ DECAP_INV_G11
XG15732 XI11_0/XI0/XI0_32/d__12_ XI11_0/XI0/XI0_32/d_12_ DECAP_INV_G11
XG15733 XI11_0/XI0/XI0_32/d__11_ XI11_0/XI0/XI0_32/d_11_ DECAP_INV_G11
XG15734 XI11_0/XI0/XI0_32/d__10_ XI11_0/XI0/XI0_32/d_10_ DECAP_INV_G11
XG15735 XI11_0/XI0/XI0_32/d__9_ XI11_0/XI0/XI0_32/d_9_ DECAP_INV_G11
XG15736 XI11_0/XI0/XI0_32/d__8_ XI11_0/XI0/XI0_32/d_8_ DECAP_INV_G11
XG15737 XI11_0/XI0/XI0_32/d__7_ XI11_0/XI0/XI0_32/d_7_ DECAP_INV_G11
XG15738 XI11_0/XI0/XI0_32/d__6_ XI11_0/XI0/XI0_32/d_6_ DECAP_INV_G11
XG15739 XI11_0/XI0/XI0_32/d__5_ XI11_0/XI0/XI0_32/d_5_ DECAP_INV_G11
XG15740 XI11_0/XI0/XI0_32/d__4_ XI11_0/XI0/XI0_32/d_4_ DECAP_INV_G11
XG15741 XI11_0/XI0/XI0_32/d__3_ XI11_0/XI0/XI0_32/d_3_ DECAP_INV_G11
XG15742 XI11_0/XI0/XI0_32/d__2_ XI11_0/XI0/XI0_32/d_2_ DECAP_INV_G11
XG15743 XI11_0/XI0/XI0_32/d__1_ XI11_0/XI0/XI0_32/d_1_ DECAP_INV_G11
XG15744 XI11_0/XI0/XI0_32/d__0_ XI11_0/XI0/XI0_32/d_0_ DECAP_INV_G11
XG15745 XI11_0/XI0/XI0_32/d_15_ XI11_0/XI0/XI0_32/d__15_ DECAP_INV_G11
XG15746 XI11_0/XI0/XI0_32/d_14_ XI11_0/XI0/XI0_32/d__14_ DECAP_INV_G11
XG15747 XI11_0/XI0/XI0_32/d_13_ XI11_0/XI0/XI0_32/d__13_ DECAP_INV_G11
XG15748 XI11_0/XI0/XI0_32/d_12_ XI11_0/XI0/XI0_32/d__12_ DECAP_INV_G11
XG15749 XI11_0/XI0/XI0_32/d_11_ XI11_0/XI0/XI0_32/d__11_ DECAP_INV_G11
XG15750 XI11_0/XI0/XI0_32/d_10_ XI11_0/XI0/XI0_32/d__10_ DECAP_INV_G11
XG15751 XI11_0/XI0/XI0_32/d_9_ XI11_0/XI0/XI0_32/d__9_ DECAP_INV_G11
XG15752 XI11_0/XI0/XI0_32/d_8_ XI11_0/XI0/XI0_32/d__8_ DECAP_INV_G11
XG15753 XI11_0/XI0/XI0_32/d_7_ XI11_0/XI0/XI0_32/d__7_ DECAP_INV_G11
XG15754 XI11_0/XI0/XI0_32/d_6_ XI11_0/XI0/XI0_32/d__6_ DECAP_INV_G11
XG15755 XI11_0/XI0/XI0_32/d_5_ XI11_0/XI0/XI0_32/d__5_ DECAP_INV_G11
XG15756 XI11_0/XI0/XI0_32/d_4_ XI11_0/XI0/XI0_32/d__4_ DECAP_INV_G11
XG15757 XI11_0/XI0/XI0_32/d_3_ XI11_0/XI0/XI0_32/d__3_ DECAP_INV_G11
XG15758 XI11_0/XI0/XI0_32/d_2_ XI11_0/XI0/XI0_32/d__2_ DECAP_INV_G11
XG15759 XI11_0/XI0/XI0_32/d_1_ XI11_0/XI0/XI0_32/d__1_ DECAP_INV_G11
XG15760 XI11_0/XI0/XI0_32/d_0_ XI11_0/XI0/XI0_32/d__0_ DECAP_INV_G11
XG15761 XI11_0/XI0/XI0_31/d__15_ XI11_0/XI0/XI0_31/d_15_ DECAP_INV_G11
XG15762 XI11_0/XI0/XI0_31/d__14_ XI11_0/XI0/XI0_31/d_14_ DECAP_INV_G11
XG15763 XI11_0/XI0/XI0_31/d__13_ XI11_0/XI0/XI0_31/d_13_ DECAP_INV_G11
XG15764 XI11_0/XI0/XI0_31/d__12_ XI11_0/XI0/XI0_31/d_12_ DECAP_INV_G11
XG15765 XI11_0/XI0/XI0_31/d__11_ XI11_0/XI0/XI0_31/d_11_ DECAP_INV_G11
XG15766 XI11_0/XI0/XI0_31/d__10_ XI11_0/XI0/XI0_31/d_10_ DECAP_INV_G11
XG15767 XI11_0/XI0/XI0_31/d__9_ XI11_0/XI0/XI0_31/d_9_ DECAP_INV_G11
XG15768 XI11_0/XI0/XI0_31/d__8_ XI11_0/XI0/XI0_31/d_8_ DECAP_INV_G11
XG15769 XI11_0/XI0/XI0_31/d__7_ XI11_0/XI0/XI0_31/d_7_ DECAP_INV_G11
XG15770 XI11_0/XI0/XI0_31/d__6_ XI11_0/XI0/XI0_31/d_6_ DECAP_INV_G11
XG15771 XI11_0/XI0/XI0_31/d__5_ XI11_0/XI0/XI0_31/d_5_ DECAP_INV_G11
XG15772 XI11_0/XI0/XI0_31/d__4_ XI11_0/XI0/XI0_31/d_4_ DECAP_INV_G11
XG15773 XI11_0/XI0/XI0_31/d__3_ XI11_0/XI0/XI0_31/d_3_ DECAP_INV_G11
XG15774 XI11_0/XI0/XI0_31/d__2_ XI11_0/XI0/XI0_31/d_2_ DECAP_INV_G11
XG15775 XI11_0/XI0/XI0_31/d__1_ XI11_0/XI0/XI0_31/d_1_ DECAP_INV_G11
XG15776 XI11_0/XI0/XI0_31/d__0_ XI11_0/XI0/XI0_31/d_0_ DECAP_INV_G11
XG15777 XI11_0/XI0/XI0_31/d_15_ XI11_0/XI0/XI0_31/d__15_ DECAP_INV_G11
XG15778 XI11_0/XI0/XI0_31/d_14_ XI11_0/XI0/XI0_31/d__14_ DECAP_INV_G11
XG15779 XI11_0/XI0/XI0_31/d_13_ XI11_0/XI0/XI0_31/d__13_ DECAP_INV_G11
XG15780 XI11_0/XI0/XI0_31/d_12_ XI11_0/XI0/XI0_31/d__12_ DECAP_INV_G11
XG15781 XI11_0/XI0/XI0_31/d_11_ XI11_0/XI0/XI0_31/d__11_ DECAP_INV_G11
XG15782 XI11_0/XI0/XI0_31/d_10_ XI11_0/XI0/XI0_31/d__10_ DECAP_INV_G11
XG15783 XI11_0/XI0/XI0_31/d_9_ XI11_0/XI0/XI0_31/d__9_ DECAP_INV_G11
XG15784 XI11_0/XI0/XI0_31/d_8_ XI11_0/XI0/XI0_31/d__8_ DECAP_INV_G11
XG15785 XI11_0/XI0/XI0_31/d_7_ XI11_0/XI0/XI0_31/d__7_ DECAP_INV_G11
XG15786 XI11_0/XI0/XI0_31/d_6_ XI11_0/XI0/XI0_31/d__6_ DECAP_INV_G11
XG15787 XI11_0/XI0/XI0_31/d_5_ XI11_0/XI0/XI0_31/d__5_ DECAP_INV_G11
XG15788 XI11_0/XI0/XI0_31/d_4_ XI11_0/XI0/XI0_31/d__4_ DECAP_INV_G11
XG15789 XI11_0/XI0/XI0_31/d_3_ XI11_0/XI0/XI0_31/d__3_ DECAP_INV_G11
XG15790 XI11_0/XI0/XI0_31/d_2_ XI11_0/XI0/XI0_31/d__2_ DECAP_INV_G11
XG15791 XI11_0/XI0/XI0_31/d_1_ XI11_0/XI0/XI0_31/d__1_ DECAP_INV_G11
XG15792 XI11_0/XI0/XI0_31/d_0_ XI11_0/XI0/XI0_31/d__0_ DECAP_INV_G11
XG15793 XI11_0/XI0/XI0_30/d__15_ XI11_0/XI0/XI0_30/d_15_ DECAP_INV_G11
XG15794 XI11_0/XI0/XI0_30/d__14_ XI11_0/XI0/XI0_30/d_14_ DECAP_INV_G11
XG15795 XI11_0/XI0/XI0_30/d__13_ XI11_0/XI0/XI0_30/d_13_ DECAP_INV_G11
XG15796 XI11_0/XI0/XI0_30/d__12_ XI11_0/XI0/XI0_30/d_12_ DECAP_INV_G11
XG15797 XI11_0/XI0/XI0_30/d__11_ XI11_0/XI0/XI0_30/d_11_ DECAP_INV_G11
XG15798 XI11_0/XI0/XI0_30/d__10_ XI11_0/XI0/XI0_30/d_10_ DECAP_INV_G11
XG15799 XI11_0/XI0/XI0_30/d__9_ XI11_0/XI0/XI0_30/d_9_ DECAP_INV_G11
XG15800 XI11_0/XI0/XI0_30/d__8_ XI11_0/XI0/XI0_30/d_8_ DECAP_INV_G11
XG15801 XI11_0/XI0/XI0_30/d__7_ XI11_0/XI0/XI0_30/d_7_ DECAP_INV_G11
XG15802 XI11_0/XI0/XI0_30/d__6_ XI11_0/XI0/XI0_30/d_6_ DECAP_INV_G11
XG15803 XI11_0/XI0/XI0_30/d__5_ XI11_0/XI0/XI0_30/d_5_ DECAP_INV_G11
XG15804 XI11_0/XI0/XI0_30/d__4_ XI11_0/XI0/XI0_30/d_4_ DECAP_INV_G11
XG15805 XI11_0/XI0/XI0_30/d__3_ XI11_0/XI0/XI0_30/d_3_ DECAP_INV_G11
XG15806 XI11_0/XI0/XI0_30/d__2_ XI11_0/XI0/XI0_30/d_2_ DECAP_INV_G11
XG15807 XI11_0/XI0/XI0_30/d__1_ XI11_0/XI0/XI0_30/d_1_ DECAP_INV_G11
XG15808 XI11_0/XI0/XI0_30/d__0_ XI11_0/XI0/XI0_30/d_0_ DECAP_INV_G11
XG15809 XI11_0/XI0/XI0_30/d_15_ XI11_0/XI0/XI0_30/d__15_ DECAP_INV_G11
XG15810 XI11_0/XI0/XI0_30/d_14_ XI11_0/XI0/XI0_30/d__14_ DECAP_INV_G11
XG15811 XI11_0/XI0/XI0_30/d_13_ XI11_0/XI0/XI0_30/d__13_ DECAP_INV_G11
XG15812 XI11_0/XI0/XI0_30/d_12_ XI11_0/XI0/XI0_30/d__12_ DECAP_INV_G11
XG15813 XI11_0/XI0/XI0_30/d_11_ XI11_0/XI0/XI0_30/d__11_ DECAP_INV_G11
XG15814 XI11_0/XI0/XI0_30/d_10_ XI11_0/XI0/XI0_30/d__10_ DECAP_INV_G11
XG15815 XI11_0/XI0/XI0_30/d_9_ XI11_0/XI0/XI0_30/d__9_ DECAP_INV_G11
XG15816 XI11_0/XI0/XI0_30/d_8_ XI11_0/XI0/XI0_30/d__8_ DECAP_INV_G11
XG15817 XI11_0/XI0/XI0_30/d_7_ XI11_0/XI0/XI0_30/d__7_ DECAP_INV_G11
XG15818 XI11_0/XI0/XI0_30/d_6_ XI11_0/XI0/XI0_30/d__6_ DECAP_INV_G11
XG15819 XI11_0/XI0/XI0_30/d_5_ XI11_0/XI0/XI0_30/d__5_ DECAP_INV_G11
XG15820 XI11_0/XI0/XI0_30/d_4_ XI11_0/XI0/XI0_30/d__4_ DECAP_INV_G11
XG15821 XI11_0/XI0/XI0_30/d_3_ XI11_0/XI0/XI0_30/d__3_ DECAP_INV_G11
XG15822 XI11_0/XI0/XI0_30/d_2_ XI11_0/XI0/XI0_30/d__2_ DECAP_INV_G11
XG15823 XI11_0/XI0/XI0_30/d_1_ XI11_0/XI0/XI0_30/d__1_ DECAP_INV_G11
XG15824 XI11_0/XI0/XI0_30/d_0_ XI11_0/XI0/XI0_30/d__0_ DECAP_INV_G11
XG15825 XI11_0/XI0/XI0_29/d__15_ XI11_0/XI0/XI0_29/d_15_ DECAP_INV_G11
XG15826 XI11_0/XI0/XI0_29/d__14_ XI11_0/XI0/XI0_29/d_14_ DECAP_INV_G11
XG15827 XI11_0/XI0/XI0_29/d__13_ XI11_0/XI0/XI0_29/d_13_ DECAP_INV_G11
XG15828 XI11_0/XI0/XI0_29/d__12_ XI11_0/XI0/XI0_29/d_12_ DECAP_INV_G11
XG15829 XI11_0/XI0/XI0_29/d__11_ XI11_0/XI0/XI0_29/d_11_ DECAP_INV_G11
XG15830 XI11_0/XI0/XI0_29/d__10_ XI11_0/XI0/XI0_29/d_10_ DECAP_INV_G11
XG15831 XI11_0/XI0/XI0_29/d__9_ XI11_0/XI0/XI0_29/d_9_ DECAP_INV_G11
XG15832 XI11_0/XI0/XI0_29/d__8_ XI11_0/XI0/XI0_29/d_8_ DECAP_INV_G11
XG15833 XI11_0/XI0/XI0_29/d__7_ XI11_0/XI0/XI0_29/d_7_ DECAP_INV_G11
XG15834 XI11_0/XI0/XI0_29/d__6_ XI11_0/XI0/XI0_29/d_6_ DECAP_INV_G11
XG15835 XI11_0/XI0/XI0_29/d__5_ XI11_0/XI0/XI0_29/d_5_ DECAP_INV_G11
XG15836 XI11_0/XI0/XI0_29/d__4_ XI11_0/XI0/XI0_29/d_4_ DECAP_INV_G11
XG15837 XI11_0/XI0/XI0_29/d__3_ XI11_0/XI0/XI0_29/d_3_ DECAP_INV_G11
XG15838 XI11_0/XI0/XI0_29/d__2_ XI11_0/XI0/XI0_29/d_2_ DECAP_INV_G11
XG15839 XI11_0/XI0/XI0_29/d__1_ XI11_0/XI0/XI0_29/d_1_ DECAP_INV_G11
XG15840 XI11_0/XI0/XI0_29/d__0_ XI11_0/XI0/XI0_29/d_0_ DECAP_INV_G11
XG15841 XI11_0/XI0/XI0_29/d_15_ XI11_0/XI0/XI0_29/d__15_ DECAP_INV_G11
XG15842 XI11_0/XI0/XI0_29/d_14_ XI11_0/XI0/XI0_29/d__14_ DECAP_INV_G11
XG15843 XI11_0/XI0/XI0_29/d_13_ XI11_0/XI0/XI0_29/d__13_ DECAP_INV_G11
XG15844 XI11_0/XI0/XI0_29/d_12_ XI11_0/XI0/XI0_29/d__12_ DECAP_INV_G11
XG15845 XI11_0/XI0/XI0_29/d_11_ XI11_0/XI0/XI0_29/d__11_ DECAP_INV_G11
XG15846 XI11_0/XI0/XI0_29/d_10_ XI11_0/XI0/XI0_29/d__10_ DECAP_INV_G11
XG15847 XI11_0/XI0/XI0_29/d_9_ XI11_0/XI0/XI0_29/d__9_ DECAP_INV_G11
XG15848 XI11_0/XI0/XI0_29/d_8_ XI11_0/XI0/XI0_29/d__8_ DECAP_INV_G11
XG15849 XI11_0/XI0/XI0_29/d_7_ XI11_0/XI0/XI0_29/d__7_ DECAP_INV_G11
XG15850 XI11_0/XI0/XI0_29/d_6_ XI11_0/XI0/XI0_29/d__6_ DECAP_INV_G11
XG15851 XI11_0/XI0/XI0_29/d_5_ XI11_0/XI0/XI0_29/d__5_ DECAP_INV_G11
XG15852 XI11_0/XI0/XI0_29/d_4_ XI11_0/XI0/XI0_29/d__4_ DECAP_INV_G11
XG15853 XI11_0/XI0/XI0_29/d_3_ XI11_0/XI0/XI0_29/d__3_ DECAP_INV_G11
XG15854 XI11_0/XI0/XI0_29/d_2_ XI11_0/XI0/XI0_29/d__2_ DECAP_INV_G11
XG15855 XI11_0/XI0/XI0_29/d_1_ XI11_0/XI0/XI0_29/d__1_ DECAP_INV_G11
XG15856 XI11_0/XI0/XI0_29/d_0_ XI11_0/XI0/XI0_29/d__0_ DECAP_INV_G11
XG15857 XI11_0/XI0/XI0_28/d__15_ XI11_0/XI0/XI0_28/d_15_ DECAP_INV_G11
XG15858 XI11_0/XI0/XI0_28/d__14_ XI11_0/XI0/XI0_28/d_14_ DECAP_INV_G11
XG15859 XI11_0/XI0/XI0_28/d__13_ XI11_0/XI0/XI0_28/d_13_ DECAP_INV_G11
XG15860 XI11_0/XI0/XI0_28/d__12_ XI11_0/XI0/XI0_28/d_12_ DECAP_INV_G11
XG15861 XI11_0/XI0/XI0_28/d__11_ XI11_0/XI0/XI0_28/d_11_ DECAP_INV_G11
XG15862 XI11_0/XI0/XI0_28/d__10_ XI11_0/XI0/XI0_28/d_10_ DECAP_INV_G11
XG15863 XI11_0/XI0/XI0_28/d__9_ XI11_0/XI0/XI0_28/d_9_ DECAP_INV_G11
XG15864 XI11_0/XI0/XI0_28/d__8_ XI11_0/XI0/XI0_28/d_8_ DECAP_INV_G11
XG15865 XI11_0/XI0/XI0_28/d__7_ XI11_0/XI0/XI0_28/d_7_ DECAP_INV_G11
XG15866 XI11_0/XI0/XI0_28/d__6_ XI11_0/XI0/XI0_28/d_6_ DECAP_INV_G11
XG15867 XI11_0/XI0/XI0_28/d__5_ XI11_0/XI0/XI0_28/d_5_ DECAP_INV_G11
XG15868 XI11_0/XI0/XI0_28/d__4_ XI11_0/XI0/XI0_28/d_4_ DECAP_INV_G11
XG15869 XI11_0/XI0/XI0_28/d__3_ XI11_0/XI0/XI0_28/d_3_ DECAP_INV_G11
XG15870 XI11_0/XI0/XI0_28/d__2_ XI11_0/XI0/XI0_28/d_2_ DECAP_INV_G11
XG15871 XI11_0/XI0/XI0_28/d__1_ XI11_0/XI0/XI0_28/d_1_ DECAP_INV_G11
XG15872 XI11_0/XI0/XI0_28/d__0_ XI11_0/XI0/XI0_28/d_0_ DECAP_INV_G11
XG15873 XI11_0/XI0/XI0_28/d_15_ XI11_0/XI0/XI0_28/d__15_ DECAP_INV_G11
XG15874 XI11_0/XI0/XI0_28/d_14_ XI11_0/XI0/XI0_28/d__14_ DECAP_INV_G11
XG15875 XI11_0/XI0/XI0_28/d_13_ XI11_0/XI0/XI0_28/d__13_ DECAP_INV_G11
XG15876 XI11_0/XI0/XI0_28/d_12_ XI11_0/XI0/XI0_28/d__12_ DECAP_INV_G11
XG15877 XI11_0/XI0/XI0_28/d_11_ XI11_0/XI0/XI0_28/d__11_ DECAP_INV_G11
XG15878 XI11_0/XI0/XI0_28/d_10_ XI11_0/XI0/XI0_28/d__10_ DECAP_INV_G11
XG15879 XI11_0/XI0/XI0_28/d_9_ XI11_0/XI0/XI0_28/d__9_ DECAP_INV_G11
XG15880 XI11_0/XI0/XI0_28/d_8_ XI11_0/XI0/XI0_28/d__8_ DECAP_INV_G11
XG15881 XI11_0/XI0/XI0_28/d_7_ XI11_0/XI0/XI0_28/d__7_ DECAP_INV_G11
XG15882 XI11_0/XI0/XI0_28/d_6_ XI11_0/XI0/XI0_28/d__6_ DECAP_INV_G11
XG15883 XI11_0/XI0/XI0_28/d_5_ XI11_0/XI0/XI0_28/d__5_ DECAP_INV_G11
XG15884 XI11_0/XI0/XI0_28/d_4_ XI11_0/XI0/XI0_28/d__4_ DECAP_INV_G11
XG15885 XI11_0/XI0/XI0_28/d_3_ XI11_0/XI0/XI0_28/d__3_ DECAP_INV_G11
XG15886 XI11_0/XI0/XI0_28/d_2_ XI11_0/XI0/XI0_28/d__2_ DECAP_INV_G11
XG15887 XI11_0/XI0/XI0_28/d_1_ XI11_0/XI0/XI0_28/d__1_ DECAP_INV_G11
XG15888 XI11_0/XI0/XI0_28/d_0_ XI11_0/XI0/XI0_28/d__0_ DECAP_INV_G11
XG15889 XI11_0/XI0/XI0_27/d__15_ XI11_0/XI0/XI0_27/d_15_ DECAP_INV_G11
XG15890 XI11_0/XI0/XI0_27/d__14_ XI11_0/XI0/XI0_27/d_14_ DECAP_INV_G11
XG15891 XI11_0/XI0/XI0_27/d__13_ XI11_0/XI0/XI0_27/d_13_ DECAP_INV_G11
XG15892 XI11_0/XI0/XI0_27/d__12_ XI11_0/XI0/XI0_27/d_12_ DECAP_INV_G11
XG15893 XI11_0/XI0/XI0_27/d__11_ XI11_0/XI0/XI0_27/d_11_ DECAP_INV_G11
XG15894 XI11_0/XI0/XI0_27/d__10_ XI11_0/XI0/XI0_27/d_10_ DECAP_INV_G11
XG15895 XI11_0/XI0/XI0_27/d__9_ XI11_0/XI0/XI0_27/d_9_ DECAP_INV_G11
XG15896 XI11_0/XI0/XI0_27/d__8_ XI11_0/XI0/XI0_27/d_8_ DECAP_INV_G11
XG15897 XI11_0/XI0/XI0_27/d__7_ XI11_0/XI0/XI0_27/d_7_ DECAP_INV_G11
XG15898 XI11_0/XI0/XI0_27/d__6_ XI11_0/XI0/XI0_27/d_6_ DECAP_INV_G11
XG15899 XI11_0/XI0/XI0_27/d__5_ XI11_0/XI0/XI0_27/d_5_ DECAP_INV_G11
XG15900 XI11_0/XI0/XI0_27/d__4_ XI11_0/XI0/XI0_27/d_4_ DECAP_INV_G11
XG15901 XI11_0/XI0/XI0_27/d__3_ XI11_0/XI0/XI0_27/d_3_ DECAP_INV_G11
XG15902 XI11_0/XI0/XI0_27/d__2_ XI11_0/XI0/XI0_27/d_2_ DECAP_INV_G11
XG15903 XI11_0/XI0/XI0_27/d__1_ XI11_0/XI0/XI0_27/d_1_ DECAP_INV_G11
XG15904 XI11_0/XI0/XI0_27/d__0_ XI11_0/XI0/XI0_27/d_0_ DECAP_INV_G11
XG15905 XI11_0/XI0/XI0_27/d_15_ XI11_0/XI0/XI0_27/d__15_ DECAP_INV_G11
XG15906 XI11_0/XI0/XI0_27/d_14_ XI11_0/XI0/XI0_27/d__14_ DECAP_INV_G11
XG15907 XI11_0/XI0/XI0_27/d_13_ XI11_0/XI0/XI0_27/d__13_ DECAP_INV_G11
XG15908 XI11_0/XI0/XI0_27/d_12_ XI11_0/XI0/XI0_27/d__12_ DECAP_INV_G11
XG15909 XI11_0/XI0/XI0_27/d_11_ XI11_0/XI0/XI0_27/d__11_ DECAP_INV_G11
XG15910 XI11_0/XI0/XI0_27/d_10_ XI11_0/XI0/XI0_27/d__10_ DECAP_INV_G11
XG15911 XI11_0/XI0/XI0_27/d_9_ XI11_0/XI0/XI0_27/d__9_ DECAP_INV_G11
XG15912 XI11_0/XI0/XI0_27/d_8_ XI11_0/XI0/XI0_27/d__8_ DECAP_INV_G11
XG15913 XI11_0/XI0/XI0_27/d_7_ XI11_0/XI0/XI0_27/d__7_ DECAP_INV_G11
XG15914 XI11_0/XI0/XI0_27/d_6_ XI11_0/XI0/XI0_27/d__6_ DECAP_INV_G11
XG15915 XI11_0/XI0/XI0_27/d_5_ XI11_0/XI0/XI0_27/d__5_ DECAP_INV_G11
XG15916 XI11_0/XI0/XI0_27/d_4_ XI11_0/XI0/XI0_27/d__4_ DECAP_INV_G11
XG15917 XI11_0/XI0/XI0_27/d_3_ XI11_0/XI0/XI0_27/d__3_ DECAP_INV_G11
XG15918 XI11_0/XI0/XI0_27/d_2_ XI11_0/XI0/XI0_27/d__2_ DECAP_INV_G11
XG15919 XI11_0/XI0/XI0_27/d_1_ XI11_0/XI0/XI0_27/d__1_ DECAP_INV_G11
XG15920 XI11_0/XI0/XI0_27/d_0_ XI11_0/XI0/XI0_27/d__0_ DECAP_INV_G11
XG15921 XI11_0/XI0/XI0_26/d__15_ XI11_0/XI0/XI0_26/d_15_ DECAP_INV_G11
XG15922 XI11_0/XI0/XI0_26/d__14_ XI11_0/XI0/XI0_26/d_14_ DECAP_INV_G11
XG15923 XI11_0/XI0/XI0_26/d__13_ XI11_0/XI0/XI0_26/d_13_ DECAP_INV_G11
XG15924 XI11_0/XI0/XI0_26/d__12_ XI11_0/XI0/XI0_26/d_12_ DECAP_INV_G11
XG15925 XI11_0/XI0/XI0_26/d__11_ XI11_0/XI0/XI0_26/d_11_ DECAP_INV_G11
XG15926 XI11_0/XI0/XI0_26/d__10_ XI11_0/XI0/XI0_26/d_10_ DECAP_INV_G11
XG15927 XI11_0/XI0/XI0_26/d__9_ XI11_0/XI0/XI0_26/d_9_ DECAP_INV_G11
XG15928 XI11_0/XI0/XI0_26/d__8_ XI11_0/XI0/XI0_26/d_8_ DECAP_INV_G11
XG15929 XI11_0/XI0/XI0_26/d__7_ XI11_0/XI0/XI0_26/d_7_ DECAP_INV_G11
XG15930 XI11_0/XI0/XI0_26/d__6_ XI11_0/XI0/XI0_26/d_6_ DECAP_INV_G11
XG15931 XI11_0/XI0/XI0_26/d__5_ XI11_0/XI0/XI0_26/d_5_ DECAP_INV_G11
XG15932 XI11_0/XI0/XI0_26/d__4_ XI11_0/XI0/XI0_26/d_4_ DECAP_INV_G11
XG15933 XI11_0/XI0/XI0_26/d__3_ XI11_0/XI0/XI0_26/d_3_ DECAP_INV_G11
XG15934 XI11_0/XI0/XI0_26/d__2_ XI11_0/XI0/XI0_26/d_2_ DECAP_INV_G11
XG15935 XI11_0/XI0/XI0_26/d__1_ XI11_0/XI0/XI0_26/d_1_ DECAP_INV_G11
XG15936 XI11_0/XI0/XI0_26/d__0_ XI11_0/XI0/XI0_26/d_0_ DECAP_INV_G11
XG15937 XI11_0/XI0/XI0_26/d_15_ XI11_0/XI0/XI0_26/d__15_ DECAP_INV_G11
XG15938 XI11_0/XI0/XI0_26/d_14_ XI11_0/XI0/XI0_26/d__14_ DECAP_INV_G11
XG15939 XI11_0/XI0/XI0_26/d_13_ XI11_0/XI0/XI0_26/d__13_ DECAP_INV_G11
XG15940 XI11_0/XI0/XI0_26/d_12_ XI11_0/XI0/XI0_26/d__12_ DECAP_INV_G11
XG15941 XI11_0/XI0/XI0_26/d_11_ XI11_0/XI0/XI0_26/d__11_ DECAP_INV_G11
XG15942 XI11_0/XI0/XI0_26/d_10_ XI11_0/XI0/XI0_26/d__10_ DECAP_INV_G11
XG15943 XI11_0/XI0/XI0_26/d_9_ XI11_0/XI0/XI0_26/d__9_ DECAP_INV_G11
XG15944 XI11_0/XI0/XI0_26/d_8_ XI11_0/XI0/XI0_26/d__8_ DECAP_INV_G11
XG15945 XI11_0/XI0/XI0_26/d_7_ XI11_0/XI0/XI0_26/d__7_ DECAP_INV_G11
XG15946 XI11_0/XI0/XI0_26/d_6_ XI11_0/XI0/XI0_26/d__6_ DECAP_INV_G11
XG15947 XI11_0/XI0/XI0_26/d_5_ XI11_0/XI0/XI0_26/d__5_ DECAP_INV_G11
XG15948 XI11_0/XI0/XI0_26/d_4_ XI11_0/XI0/XI0_26/d__4_ DECAP_INV_G11
XG15949 XI11_0/XI0/XI0_26/d_3_ XI11_0/XI0/XI0_26/d__3_ DECAP_INV_G11
XG15950 XI11_0/XI0/XI0_26/d_2_ XI11_0/XI0/XI0_26/d__2_ DECAP_INV_G11
XG15951 XI11_0/XI0/XI0_26/d_1_ XI11_0/XI0/XI0_26/d__1_ DECAP_INV_G11
XG15952 XI11_0/XI0/XI0_26/d_0_ XI11_0/XI0/XI0_26/d__0_ DECAP_INV_G11
XG15953 XI11_0/XI0/XI0_25/d__15_ XI11_0/XI0/XI0_25/d_15_ DECAP_INV_G11
XG15954 XI11_0/XI0/XI0_25/d__14_ XI11_0/XI0/XI0_25/d_14_ DECAP_INV_G11
XG15955 XI11_0/XI0/XI0_25/d__13_ XI11_0/XI0/XI0_25/d_13_ DECAP_INV_G11
XG15956 XI11_0/XI0/XI0_25/d__12_ XI11_0/XI0/XI0_25/d_12_ DECAP_INV_G11
XG15957 XI11_0/XI0/XI0_25/d__11_ XI11_0/XI0/XI0_25/d_11_ DECAP_INV_G11
XG15958 XI11_0/XI0/XI0_25/d__10_ XI11_0/XI0/XI0_25/d_10_ DECAP_INV_G11
XG15959 XI11_0/XI0/XI0_25/d__9_ XI11_0/XI0/XI0_25/d_9_ DECAP_INV_G11
XG15960 XI11_0/XI0/XI0_25/d__8_ XI11_0/XI0/XI0_25/d_8_ DECAP_INV_G11
XG15961 XI11_0/XI0/XI0_25/d__7_ XI11_0/XI0/XI0_25/d_7_ DECAP_INV_G11
XG15962 XI11_0/XI0/XI0_25/d__6_ XI11_0/XI0/XI0_25/d_6_ DECAP_INV_G11
XG15963 XI11_0/XI0/XI0_25/d__5_ XI11_0/XI0/XI0_25/d_5_ DECAP_INV_G11
XG15964 XI11_0/XI0/XI0_25/d__4_ XI11_0/XI0/XI0_25/d_4_ DECAP_INV_G11
XG15965 XI11_0/XI0/XI0_25/d__3_ XI11_0/XI0/XI0_25/d_3_ DECAP_INV_G11
XG15966 XI11_0/XI0/XI0_25/d__2_ XI11_0/XI0/XI0_25/d_2_ DECAP_INV_G11
XG15967 XI11_0/XI0/XI0_25/d__1_ XI11_0/XI0/XI0_25/d_1_ DECAP_INV_G11
XG15968 XI11_0/XI0/XI0_25/d__0_ XI11_0/XI0/XI0_25/d_0_ DECAP_INV_G11
XG15969 XI11_0/XI0/XI0_25/d_15_ XI11_0/XI0/XI0_25/d__15_ DECAP_INV_G11
XG15970 XI11_0/XI0/XI0_25/d_14_ XI11_0/XI0/XI0_25/d__14_ DECAP_INV_G11
XG15971 XI11_0/XI0/XI0_25/d_13_ XI11_0/XI0/XI0_25/d__13_ DECAP_INV_G11
XG15972 XI11_0/XI0/XI0_25/d_12_ XI11_0/XI0/XI0_25/d__12_ DECAP_INV_G11
XG15973 XI11_0/XI0/XI0_25/d_11_ XI11_0/XI0/XI0_25/d__11_ DECAP_INV_G11
XG15974 XI11_0/XI0/XI0_25/d_10_ XI11_0/XI0/XI0_25/d__10_ DECAP_INV_G11
XG15975 XI11_0/XI0/XI0_25/d_9_ XI11_0/XI0/XI0_25/d__9_ DECAP_INV_G11
XG15976 XI11_0/XI0/XI0_25/d_8_ XI11_0/XI0/XI0_25/d__8_ DECAP_INV_G11
XG15977 XI11_0/XI0/XI0_25/d_7_ XI11_0/XI0/XI0_25/d__7_ DECAP_INV_G11
XG15978 XI11_0/XI0/XI0_25/d_6_ XI11_0/XI0/XI0_25/d__6_ DECAP_INV_G11
XG15979 XI11_0/XI0/XI0_25/d_5_ XI11_0/XI0/XI0_25/d__5_ DECAP_INV_G11
XG15980 XI11_0/XI0/XI0_25/d_4_ XI11_0/XI0/XI0_25/d__4_ DECAP_INV_G11
XG15981 XI11_0/XI0/XI0_25/d_3_ XI11_0/XI0/XI0_25/d__3_ DECAP_INV_G11
XG15982 XI11_0/XI0/XI0_25/d_2_ XI11_0/XI0/XI0_25/d__2_ DECAP_INV_G11
XG15983 XI11_0/XI0/XI0_25/d_1_ XI11_0/XI0/XI0_25/d__1_ DECAP_INV_G11
XG15984 XI11_0/XI0/XI0_25/d_0_ XI11_0/XI0/XI0_25/d__0_ DECAP_INV_G11
XG15985 XI11_0/XI0/XI0_24/d__15_ XI11_0/XI0/XI0_24/d_15_ DECAP_INV_G11
XG15986 XI11_0/XI0/XI0_24/d__14_ XI11_0/XI0/XI0_24/d_14_ DECAP_INV_G11
XG15987 XI11_0/XI0/XI0_24/d__13_ XI11_0/XI0/XI0_24/d_13_ DECAP_INV_G11
XG15988 XI11_0/XI0/XI0_24/d__12_ XI11_0/XI0/XI0_24/d_12_ DECAP_INV_G11
XG15989 XI11_0/XI0/XI0_24/d__11_ XI11_0/XI0/XI0_24/d_11_ DECAP_INV_G11
XG15990 XI11_0/XI0/XI0_24/d__10_ XI11_0/XI0/XI0_24/d_10_ DECAP_INV_G11
XG15991 XI11_0/XI0/XI0_24/d__9_ XI11_0/XI0/XI0_24/d_9_ DECAP_INV_G11
XG15992 XI11_0/XI0/XI0_24/d__8_ XI11_0/XI0/XI0_24/d_8_ DECAP_INV_G11
XG15993 XI11_0/XI0/XI0_24/d__7_ XI11_0/XI0/XI0_24/d_7_ DECAP_INV_G11
XG15994 XI11_0/XI0/XI0_24/d__6_ XI11_0/XI0/XI0_24/d_6_ DECAP_INV_G11
XG15995 XI11_0/XI0/XI0_24/d__5_ XI11_0/XI0/XI0_24/d_5_ DECAP_INV_G11
XG15996 XI11_0/XI0/XI0_24/d__4_ XI11_0/XI0/XI0_24/d_4_ DECAP_INV_G11
XG15997 XI11_0/XI0/XI0_24/d__3_ XI11_0/XI0/XI0_24/d_3_ DECAP_INV_G11
XG15998 XI11_0/XI0/XI0_24/d__2_ XI11_0/XI0/XI0_24/d_2_ DECAP_INV_G11
XG15999 XI11_0/XI0/XI0_24/d__1_ XI11_0/XI0/XI0_24/d_1_ DECAP_INV_G11
XG16000 XI11_0/XI0/XI0_24/d__0_ XI11_0/XI0/XI0_24/d_0_ DECAP_INV_G11
XG16001 XI11_0/XI0/XI0_24/d_15_ XI11_0/XI0/XI0_24/d__15_ DECAP_INV_G11
XG16002 XI11_0/XI0/XI0_24/d_14_ XI11_0/XI0/XI0_24/d__14_ DECAP_INV_G11
XG16003 XI11_0/XI0/XI0_24/d_13_ XI11_0/XI0/XI0_24/d__13_ DECAP_INV_G11
XG16004 XI11_0/XI0/XI0_24/d_12_ XI11_0/XI0/XI0_24/d__12_ DECAP_INV_G11
XG16005 XI11_0/XI0/XI0_24/d_11_ XI11_0/XI0/XI0_24/d__11_ DECAP_INV_G11
XG16006 XI11_0/XI0/XI0_24/d_10_ XI11_0/XI0/XI0_24/d__10_ DECAP_INV_G11
XG16007 XI11_0/XI0/XI0_24/d_9_ XI11_0/XI0/XI0_24/d__9_ DECAP_INV_G11
XG16008 XI11_0/XI0/XI0_24/d_8_ XI11_0/XI0/XI0_24/d__8_ DECAP_INV_G11
XG16009 XI11_0/XI0/XI0_24/d_7_ XI11_0/XI0/XI0_24/d__7_ DECAP_INV_G11
XG16010 XI11_0/XI0/XI0_24/d_6_ XI11_0/XI0/XI0_24/d__6_ DECAP_INV_G11
XG16011 XI11_0/XI0/XI0_24/d_5_ XI11_0/XI0/XI0_24/d__5_ DECAP_INV_G11
XG16012 XI11_0/XI0/XI0_24/d_4_ XI11_0/XI0/XI0_24/d__4_ DECAP_INV_G11
XG16013 XI11_0/XI0/XI0_24/d_3_ XI11_0/XI0/XI0_24/d__3_ DECAP_INV_G11
XG16014 XI11_0/XI0/XI0_24/d_2_ XI11_0/XI0/XI0_24/d__2_ DECAP_INV_G11
XG16015 XI11_0/XI0/XI0_24/d_1_ XI11_0/XI0/XI0_24/d__1_ DECAP_INV_G11
XG16016 XI11_0/XI0/XI0_24/d_0_ XI11_0/XI0/XI0_24/d__0_ DECAP_INV_G11
XG16017 XI11_0/XI0/XI0_23/d__15_ XI11_0/XI0/XI0_23/d_15_ DECAP_INV_G11
XG16018 XI11_0/XI0/XI0_23/d__14_ XI11_0/XI0/XI0_23/d_14_ DECAP_INV_G11
XG16019 XI11_0/XI0/XI0_23/d__13_ XI11_0/XI0/XI0_23/d_13_ DECAP_INV_G11
XG16020 XI11_0/XI0/XI0_23/d__12_ XI11_0/XI0/XI0_23/d_12_ DECAP_INV_G11
XG16021 XI11_0/XI0/XI0_23/d__11_ XI11_0/XI0/XI0_23/d_11_ DECAP_INV_G11
XG16022 XI11_0/XI0/XI0_23/d__10_ XI11_0/XI0/XI0_23/d_10_ DECAP_INV_G11
XG16023 XI11_0/XI0/XI0_23/d__9_ XI11_0/XI0/XI0_23/d_9_ DECAP_INV_G11
XG16024 XI11_0/XI0/XI0_23/d__8_ XI11_0/XI0/XI0_23/d_8_ DECAP_INV_G11
XG16025 XI11_0/XI0/XI0_23/d__7_ XI11_0/XI0/XI0_23/d_7_ DECAP_INV_G11
XG16026 XI11_0/XI0/XI0_23/d__6_ XI11_0/XI0/XI0_23/d_6_ DECAP_INV_G11
XG16027 XI11_0/XI0/XI0_23/d__5_ XI11_0/XI0/XI0_23/d_5_ DECAP_INV_G11
XG16028 XI11_0/XI0/XI0_23/d__4_ XI11_0/XI0/XI0_23/d_4_ DECAP_INV_G11
XG16029 XI11_0/XI0/XI0_23/d__3_ XI11_0/XI0/XI0_23/d_3_ DECAP_INV_G11
XG16030 XI11_0/XI0/XI0_23/d__2_ XI11_0/XI0/XI0_23/d_2_ DECAP_INV_G11
XG16031 XI11_0/XI0/XI0_23/d__1_ XI11_0/XI0/XI0_23/d_1_ DECAP_INV_G11
XG16032 XI11_0/XI0/XI0_23/d__0_ XI11_0/XI0/XI0_23/d_0_ DECAP_INV_G11
XG16033 XI11_0/XI0/XI0_23/d_15_ XI11_0/XI0/XI0_23/d__15_ DECAP_INV_G11
XG16034 XI11_0/XI0/XI0_23/d_14_ XI11_0/XI0/XI0_23/d__14_ DECAP_INV_G11
XG16035 XI11_0/XI0/XI0_23/d_13_ XI11_0/XI0/XI0_23/d__13_ DECAP_INV_G11
XG16036 XI11_0/XI0/XI0_23/d_12_ XI11_0/XI0/XI0_23/d__12_ DECAP_INV_G11
XG16037 XI11_0/XI0/XI0_23/d_11_ XI11_0/XI0/XI0_23/d__11_ DECAP_INV_G11
XG16038 XI11_0/XI0/XI0_23/d_10_ XI11_0/XI0/XI0_23/d__10_ DECAP_INV_G11
XG16039 XI11_0/XI0/XI0_23/d_9_ XI11_0/XI0/XI0_23/d__9_ DECAP_INV_G11
XG16040 XI11_0/XI0/XI0_23/d_8_ XI11_0/XI0/XI0_23/d__8_ DECAP_INV_G11
XG16041 XI11_0/XI0/XI0_23/d_7_ XI11_0/XI0/XI0_23/d__7_ DECAP_INV_G11
XG16042 XI11_0/XI0/XI0_23/d_6_ XI11_0/XI0/XI0_23/d__6_ DECAP_INV_G11
XG16043 XI11_0/XI0/XI0_23/d_5_ XI11_0/XI0/XI0_23/d__5_ DECAP_INV_G11
XG16044 XI11_0/XI0/XI0_23/d_4_ XI11_0/XI0/XI0_23/d__4_ DECAP_INV_G11
XG16045 XI11_0/XI0/XI0_23/d_3_ XI11_0/XI0/XI0_23/d__3_ DECAP_INV_G11
XG16046 XI11_0/XI0/XI0_23/d_2_ XI11_0/XI0/XI0_23/d__2_ DECAP_INV_G11
XG16047 XI11_0/XI0/XI0_23/d_1_ XI11_0/XI0/XI0_23/d__1_ DECAP_INV_G11
XG16048 XI11_0/XI0/XI0_23/d_0_ XI11_0/XI0/XI0_23/d__0_ DECAP_INV_G11
XG16049 XI11_0/XI0/XI0_22/d__15_ XI11_0/XI0/XI0_22/d_15_ DECAP_INV_G11
XG16050 XI11_0/XI0/XI0_22/d__14_ XI11_0/XI0/XI0_22/d_14_ DECAP_INV_G11
XG16051 XI11_0/XI0/XI0_22/d__13_ XI11_0/XI0/XI0_22/d_13_ DECAP_INV_G11
XG16052 XI11_0/XI0/XI0_22/d__12_ XI11_0/XI0/XI0_22/d_12_ DECAP_INV_G11
XG16053 XI11_0/XI0/XI0_22/d__11_ XI11_0/XI0/XI0_22/d_11_ DECAP_INV_G11
XG16054 XI11_0/XI0/XI0_22/d__10_ XI11_0/XI0/XI0_22/d_10_ DECAP_INV_G11
XG16055 XI11_0/XI0/XI0_22/d__9_ XI11_0/XI0/XI0_22/d_9_ DECAP_INV_G11
XG16056 XI11_0/XI0/XI0_22/d__8_ XI11_0/XI0/XI0_22/d_8_ DECAP_INV_G11
XG16057 XI11_0/XI0/XI0_22/d__7_ XI11_0/XI0/XI0_22/d_7_ DECAP_INV_G11
XG16058 XI11_0/XI0/XI0_22/d__6_ XI11_0/XI0/XI0_22/d_6_ DECAP_INV_G11
XG16059 XI11_0/XI0/XI0_22/d__5_ XI11_0/XI0/XI0_22/d_5_ DECAP_INV_G11
XG16060 XI11_0/XI0/XI0_22/d__4_ XI11_0/XI0/XI0_22/d_4_ DECAP_INV_G11
XG16061 XI11_0/XI0/XI0_22/d__3_ XI11_0/XI0/XI0_22/d_3_ DECAP_INV_G11
XG16062 XI11_0/XI0/XI0_22/d__2_ XI11_0/XI0/XI0_22/d_2_ DECAP_INV_G11
XG16063 XI11_0/XI0/XI0_22/d__1_ XI11_0/XI0/XI0_22/d_1_ DECAP_INV_G11
XG16064 XI11_0/XI0/XI0_22/d__0_ XI11_0/XI0/XI0_22/d_0_ DECAP_INV_G11
XG16065 XI11_0/XI0/XI0_22/d_15_ XI11_0/XI0/XI0_22/d__15_ DECAP_INV_G11
XG16066 XI11_0/XI0/XI0_22/d_14_ XI11_0/XI0/XI0_22/d__14_ DECAP_INV_G11
XG16067 XI11_0/XI0/XI0_22/d_13_ XI11_0/XI0/XI0_22/d__13_ DECAP_INV_G11
XG16068 XI11_0/XI0/XI0_22/d_12_ XI11_0/XI0/XI0_22/d__12_ DECAP_INV_G11
XG16069 XI11_0/XI0/XI0_22/d_11_ XI11_0/XI0/XI0_22/d__11_ DECAP_INV_G11
XG16070 XI11_0/XI0/XI0_22/d_10_ XI11_0/XI0/XI0_22/d__10_ DECAP_INV_G11
XG16071 XI11_0/XI0/XI0_22/d_9_ XI11_0/XI0/XI0_22/d__9_ DECAP_INV_G11
XG16072 XI11_0/XI0/XI0_22/d_8_ XI11_0/XI0/XI0_22/d__8_ DECAP_INV_G11
XG16073 XI11_0/XI0/XI0_22/d_7_ XI11_0/XI0/XI0_22/d__7_ DECAP_INV_G11
XG16074 XI11_0/XI0/XI0_22/d_6_ XI11_0/XI0/XI0_22/d__6_ DECAP_INV_G11
XG16075 XI11_0/XI0/XI0_22/d_5_ XI11_0/XI0/XI0_22/d__5_ DECAP_INV_G11
XG16076 XI11_0/XI0/XI0_22/d_4_ XI11_0/XI0/XI0_22/d__4_ DECAP_INV_G11
XG16077 XI11_0/XI0/XI0_22/d_3_ XI11_0/XI0/XI0_22/d__3_ DECAP_INV_G11
XG16078 XI11_0/XI0/XI0_22/d_2_ XI11_0/XI0/XI0_22/d__2_ DECAP_INV_G11
XG16079 XI11_0/XI0/XI0_22/d_1_ XI11_0/XI0/XI0_22/d__1_ DECAP_INV_G11
XG16080 XI11_0/XI0/XI0_22/d_0_ XI11_0/XI0/XI0_22/d__0_ DECAP_INV_G11
XG16081 XI11_0/XI0/XI0_21/d__15_ XI11_0/XI0/XI0_21/d_15_ DECAP_INV_G11
XG16082 XI11_0/XI0/XI0_21/d__14_ XI11_0/XI0/XI0_21/d_14_ DECAP_INV_G11
XG16083 XI11_0/XI0/XI0_21/d__13_ XI11_0/XI0/XI0_21/d_13_ DECAP_INV_G11
XG16084 XI11_0/XI0/XI0_21/d__12_ XI11_0/XI0/XI0_21/d_12_ DECAP_INV_G11
XG16085 XI11_0/XI0/XI0_21/d__11_ XI11_0/XI0/XI0_21/d_11_ DECAP_INV_G11
XG16086 XI11_0/XI0/XI0_21/d__10_ XI11_0/XI0/XI0_21/d_10_ DECAP_INV_G11
XG16087 XI11_0/XI0/XI0_21/d__9_ XI11_0/XI0/XI0_21/d_9_ DECAP_INV_G11
XG16088 XI11_0/XI0/XI0_21/d__8_ XI11_0/XI0/XI0_21/d_8_ DECAP_INV_G11
XG16089 XI11_0/XI0/XI0_21/d__7_ XI11_0/XI0/XI0_21/d_7_ DECAP_INV_G11
XG16090 XI11_0/XI0/XI0_21/d__6_ XI11_0/XI0/XI0_21/d_6_ DECAP_INV_G11
XG16091 XI11_0/XI0/XI0_21/d__5_ XI11_0/XI0/XI0_21/d_5_ DECAP_INV_G11
XG16092 XI11_0/XI0/XI0_21/d__4_ XI11_0/XI0/XI0_21/d_4_ DECAP_INV_G11
XG16093 XI11_0/XI0/XI0_21/d__3_ XI11_0/XI0/XI0_21/d_3_ DECAP_INV_G11
XG16094 XI11_0/XI0/XI0_21/d__2_ XI11_0/XI0/XI0_21/d_2_ DECAP_INV_G11
XG16095 XI11_0/XI0/XI0_21/d__1_ XI11_0/XI0/XI0_21/d_1_ DECAP_INV_G11
XG16096 XI11_0/XI0/XI0_21/d__0_ XI11_0/XI0/XI0_21/d_0_ DECAP_INV_G11
XG16097 XI11_0/XI0/XI0_21/d_15_ XI11_0/XI0/XI0_21/d__15_ DECAP_INV_G11
XG16098 XI11_0/XI0/XI0_21/d_14_ XI11_0/XI0/XI0_21/d__14_ DECAP_INV_G11
XG16099 XI11_0/XI0/XI0_21/d_13_ XI11_0/XI0/XI0_21/d__13_ DECAP_INV_G11
XG16100 XI11_0/XI0/XI0_21/d_12_ XI11_0/XI0/XI0_21/d__12_ DECAP_INV_G11
XG16101 XI11_0/XI0/XI0_21/d_11_ XI11_0/XI0/XI0_21/d__11_ DECAP_INV_G11
XG16102 XI11_0/XI0/XI0_21/d_10_ XI11_0/XI0/XI0_21/d__10_ DECAP_INV_G11
XG16103 XI11_0/XI0/XI0_21/d_9_ XI11_0/XI0/XI0_21/d__9_ DECAP_INV_G11
XG16104 XI11_0/XI0/XI0_21/d_8_ XI11_0/XI0/XI0_21/d__8_ DECAP_INV_G11
XG16105 XI11_0/XI0/XI0_21/d_7_ XI11_0/XI0/XI0_21/d__7_ DECAP_INV_G11
XG16106 XI11_0/XI0/XI0_21/d_6_ XI11_0/XI0/XI0_21/d__6_ DECAP_INV_G11
XG16107 XI11_0/XI0/XI0_21/d_5_ XI11_0/XI0/XI0_21/d__5_ DECAP_INV_G11
XG16108 XI11_0/XI0/XI0_21/d_4_ XI11_0/XI0/XI0_21/d__4_ DECAP_INV_G11
XG16109 XI11_0/XI0/XI0_21/d_3_ XI11_0/XI0/XI0_21/d__3_ DECAP_INV_G11
XG16110 XI11_0/XI0/XI0_21/d_2_ XI11_0/XI0/XI0_21/d__2_ DECAP_INV_G11
XG16111 XI11_0/XI0/XI0_21/d_1_ XI11_0/XI0/XI0_21/d__1_ DECAP_INV_G11
XG16112 XI11_0/XI0/XI0_21/d_0_ XI11_0/XI0/XI0_21/d__0_ DECAP_INV_G11
XG16113 XI11_0/XI0/XI0_20/d__15_ XI11_0/XI0/XI0_20/d_15_ DECAP_INV_G11
XG16114 XI11_0/XI0/XI0_20/d__14_ XI11_0/XI0/XI0_20/d_14_ DECAP_INV_G11
XG16115 XI11_0/XI0/XI0_20/d__13_ XI11_0/XI0/XI0_20/d_13_ DECAP_INV_G11
XG16116 XI11_0/XI0/XI0_20/d__12_ XI11_0/XI0/XI0_20/d_12_ DECAP_INV_G11
XG16117 XI11_0/XI0/XI0_20/d__11_ XI11_0/XI0/XI0_20/d_11_ DECAP_INV_G11
XG16118 XI11_0/XI0/XI0_20/d__10_ XI11_0/XI0/XI0_20/d_10_ DECAP_INV_G11
XG16119 XI11_0/XI0/XI0_20/d__9_ XI11_0/XI0/XI0_20/d_9_ DECAP_INV_G11
XG16120 XI11_0/XI0/XI0_20/d__8_ XI11_0/XI0/XI0_20/d_8_ DECAP_INV_G11
XG16121 XI11_0/XI0/XI0_20/d__7_ XI11_0/XI0/XI0_20/d_7_ DECAP_INV_G11
XG16122 XI11_0/XI0/XI0_20/d__6_ XI11_0/XI0/XI0_20/d_6_ DECAP_INV_G11
XG16123 XI11_0/XI0/XI0_20/d__5_ XI11_0/XI0/XI0_20/d_5_ DECAP_INV_G11
XG16124 XI11_0/XI0/XI0_20/d__4_ XI11_0/XI0/XI0_20/d_4_ DECAP_INV_G11
XG16125 XI11_0/XI0/XI0_20/d__3_ XI11_0/XI0/XI0_20/d_3_ DECAP_INV_G11
XG16126 XI11_0/XI0/XI0_20/d__2_ XI11_0/XI0/XI0_20/d_2_ DECAP_INV_G11
XG16127 XI11_0/XI0/XI0_20/d__1_ XI11_0/XI0/XI0_20/d_1_ DECAP_INV_G11
XG16128 XI11_0/XI0/XI0_20/d__0_ XI11_0/XI0/XI0_20/d_0_ DECAP_INV_G11
XG16129 XI11_0/XI0/XI0_20/d_15_ XI11_0/XI0/XI0_20/d__15_ DECAP_INV_G11
XG16130 XI11_0/XI0/XI0_20/d_14_ XI11_0/XI0/XI0_20/d__14_ DECAP_INV_G11
XG16131 XI11_0/XI0/XI0_20/d_13_ XI11_0/XI0/XI0_20/d__13_ DECAP_INV_G11
XG16132 XI11_0/XI0/XI0_20/d_12_ XI11_0/XI0/XI0_20/d__12_ DECAP_INV_G11
XG16133 XI11_0/XI0/XI0_20/d_11_ XI11_0/XI0/XI0_20/d__11_ DECAP_INV_G11
XG16134 XI11_0/XI0/XI0_20/d_10_ XI11_0/XI0/XI0_20/d__10_ DECAP_INV_G11
XG16135 XI11_0/XI0/XI0_20/d_9_ XI11_0/XI0/XI0_20/d__9_ DECAP_INV_G11
XG16136 XI11_0/XI0/XI0_20/d_8_ XI11_0/XI0/XI0_20/d__8_ DECAP_INV_G11
XG16137 XI11_0/XI0/XI0_20/d_7_ XI11_0/XI0/XI0_20/d__7_ DECAP_INV_G11
XG16138 XI11_0/XI0/XI0_20/d_6_ XI11_0/XI0/XI0_20/d__6_ DECAP_INV_G11
XG16139 XI11_0/XI0/XI0_20/d_5_ XI11_0/XI0/XI0_20/d__5_ DECAP_INV_G11
XG16140 XI11_0/XI0/XI0_20/d_4_ XI11_0/XI0/XI0_20/d__4_ DECAP_INV_G11
XG16141 XI11_0/XI0/XI0_20/d_3_ XI11_0/XI0/XI0_20/d__3_ DECAP_INV_G11
XG16142 XI11_0/XI0/XI0_20/d_2_ XI11_0/XI0/XI0_20/d__2_ DECAP_INV_G11
XG16143 XI11_0/XI0/XI0_20/d_1_ XI11_0/XI0/XI0_20/d__1_ DECAP_INV_G11
XG16144 XI11_0/XI0/XI0_20/d_0_ XI11_0/XI0/XI0_20/d__0_ DECAP_INV_G11
XG16145 XI11_0/XI0/XI0_19/d__15_ XI11_0/XI0/XI0_19/d_15_ DECAP_INV_G11
XG16146 XI11_0/XI0/XI0_19/d__14_ XI11_0/XI0/XI0_19/d_14_ DECAP_INV_G11
XG16147 XI11_0/XI0/XI0_19/d__13_ XI11_0/XI0/XI0_19/d_13_ DECAP_INV_G11
XG16148 XI11_0/XI0/XI0_19/d__12_ XI11_0/XI0/XI0_19/d_12_ DECAP_INV_G11
XG16149 XI11_0/XI0/XI0_19/d__11_ XI11_0/XI0/XI0_19/d_11_ DECAP_INV_G11
XG16150 XI11_0/XI0/XI0_19/d__10_ XI11_0/XI0/XI0_19/d_10_ DECAP_INV_G11
XG16151 XI11_0/XI0/XI0_19/d__9_ XI11_0/XI0/XI0_19/d_9_ DECAP_INV_G11
XG16152 XI11_0/XI0/XI0_19/d__8_ XI11_0/XI0/XI0_19/d_8_ DECAP_INV_G11
XG16153 XI11_0/XI0/XI0_19/d__7_ XI11_0/XI0/XI0_19/d_7_ DECAP_INV_G11
XG16154 XI11_0/XI0/XI0_19/d__6_ XI11_0/XI0/XI0_19/d_6_ DECAP_INV_G11
XG16155 XI11_0/XI0/XI0_19/d__5_ XI11_0/XI0/XI0_19/d_5_ DECAP_INV_G11
XG16156 XI11_0/XI0/XI0_19/d__4_ XI11_0/XI0/XI0_19/d_4_ DECAP_INV_G11
XG16157 XI11_0/XI0/XI0_19/d__3_ XI11_0/XI0/XI0_19/d_3_ DECAP_INV_G11
XG16158 XI11_0/XI0/XI0_19/d__2_ XI11_0/XI0/XI0_19/d_2_ DECAP_INV_G11
XG16159 XI11_0/XI0/XI0_19/d__1_ XI11_0/XI0/XI0_19/d_1_ DECAP_INV_G11
XG16160 XI11_0/XI0/XI0_19/d__0_ XI11_0/XI0/XI0_19/d_0_ DECAP_INV_G11
XG16161 XI11_0/XI0/XI0_19/d_15_ XI11_0/XI0/XI0_19/d__15_ DECAP_INV_G11
XG16162 XI11_0/XI0/XI0_19/d_14_ XI11_0/XI0/XI0_19/d__14_ DECAP_INV_G11
XG16163 XI11_0/XI0/XI0_19/d_13_ XI11_0/XI0/XI0_19/d__13_ DECAP_INV_G11
XG16164 XI11_0/XI0/XI0_19/d_12_ XI11_0/XI0/XI0_19/d__12_ DECAP_INV_G11
XG16165 XI11_0/XI0/XI0_19/d_11_ XI11_0/XI0/XI0_19/d__11_ DECAP_INV_G11
XG16166 XI11_0/XI0/XI0_19/d_10_ XI11_0/XI0/XI0_19/d__10_ DECAP_INV_G11
XG16167 XI11_0/XI0/XI0_19/d_9_ XI11_0/XI0/XI0_19/d__9_ DECAP_INV_G11
XG16168 XI11_0/XI0/XI0_19/d_8_ XI11_0/XI0/XI0_19/d__8_ DECAP_INV_G11
XG16169 XI11_0/XI0/XI0_19/d_7_ XI11_0/XI0/XI0_19/d__7_ DECAP_INV_G11
XG16170 XI11_0/XI0/XI0_19/d_6_ XI11_0/XI0/XI0_19/d__6_ DECAP_INV_G11
XG16171 XI11_0/XI0/XI0_19/d_5_ XI11_0/XI0/XI0_19/d__5_ DECAP_INV_G11
XG16172 XI11_0/XI0/XI0_19/d_4_ XI11_0/XI0/XI0_19/d__4_ DECAP_INV_G11
XG16173 XI11_0/XI0/XI0_19/d_3_ XI11_0/XI0/XI0_19/d__3_ DECAP_INV_G11
XG16174 XI11_0/XI0/XI0_19/d_2_ XI11_0/XI0/XI0_19/d__2_ DECAP_INV_G11
XG16175 XI11_0/XI0/XI0_19/d_1_ XI11_0/XI0/XI0_19/d__1_ DECAP_INV_G11
XG16176 XI11_0/XI0/XI0_19/d_0_ XI11_0/XI0/XI0_19/d__0_ DECAP_INV_G11
XG16177 XI11_0/XI0/XI0_18/d__15_ XI11_0/XI0/XI0_18/d_15_ DECAP_INV_G11
XG16178 XI11_0/XI0/XI0_18/d__14_ XI11_0/XI0/XI0_18/d_14_ DECAP_INV_G11
XG16179 XI11_0/XI0/XI0_18/d__13_ XI11_0/XI0/XI0_18/d_13_ DECAP_INV_G11
XG16180 XI11_0/XI0/XI0_18/d__12_ XI11_0/XI0/XI0_18/d_12_ DECAP_INV_G11
XG16181 XI11_0/XI0/XI0_18/d__11_ XI11_0/XI0/XI0_18/d_11_ DECAP_INV_G11
XG16182 XI11_0/XI0/XI0_18/d__10_ XI11_0/XI0/XI0_18/d_10_ DECAP_INV_G11
XG16183 XI11_0/XI0/XI0_18/d__9_ XI11_0/XI0/XI0_18/d_9_ DECAP_INV_G11
XG16184 XI11_0/XI0/XI0_18/d__8_ XI11_0/XI0/XI0_18/d_8_ DECAP_INV_G11
XG16185 XI11_0/XI0/XI0_18/d__7_ XI11_0/XI0/XI0_18/d_7_ DECAP_INV_G11
XG16186 XI11_0/XI0/XI0_18/d__6_ XI11_0/XI0/XI0_18/d_6_ DECAP_INV_G11
XG16187 XI11_0/XI0/XI0_18/d__5_ XI11_0/XI0/XI0_18/d_5_ DECAP_INV_G11
XG16188 XI11_0/XI0/XI0_18/d__4_ XI11_0/XI0/XI0_18/d_4_ DECAP_INV_G11
XG16189 XI11_0/XI0/XI0_18/d__3_ XI11_0/XI0/XI0_18/d_3_ DECAP_INV_G11
XG16190 XI11_0/XI0/XI0_18/d__2_ XI11_0/XI0/XI0_18/d_2_ DECAP_INV_G11
XG16191 XI11_0/XI0/XI0_18/d__1_ XI11_0/XI0/XI0_18/d_1_ DECAP_INV_G11
XG16192 XI11_0/XI0/XI0_18/d__0_ XI11_0/XI0/XI0_18/d_0_ DECAP_INV_G11
XG16193 XI11_0/XI0/XI0_18/d_15_ XI11_0/XI0/XI0_18/d__15_ DECAP_INV_G11
XG16194 XI11_0/XI0/XI0_18/d_14_ XI11_0/XI0/XI0_18/d__14_ DECAP_INV_G11
XG16195 XI11_0/XI0/XI0_18/d_13_ XI11_0/XI0/XI0_18/d__13_ DECAP_INV_G11
XG16196 XI11_0/XI0/XI0_18/d_12_ XI11_0/XI0/XI0_18/d__12_ DECAP_INV_G11
XG16197 XI11_0/XI0/XI0_18/d_11_ XI11_0/XI0/XI0_18/d__11_ DECAP_INV_G11
XG16198 XI11_0/XI0/XI0_18/d_10_ XI11_0/XI0/XI0_18/d__10_ DECAP_INV_G11
XG16199 XI11_0/XI0/XI0_18/d_9_ XI11_0/XI0/XI0_18/d__9_ DECAP_INV_G11
XG16200 XI11_0/XI0/XI0_18/d_8_ XI11_0/XI0/XI0_18/d__8_ DECAP_INV_G11
XG16201 XI11_0/XI0/XI0_18/d_7_ XI11_0/XI0/XI0_18/d__7_ DECAP_INV_G11
XG16202 XI11_0/XI0/XI0_18/d_6_ XI11_0/XI0/XI0_18/d__6_ DECAP_INV_G11
XG16203 XI11_0/XI0/XI0_18/d_5_ XI11_0/XI0/XI0_18/d__5_ DECAP_INV_G11
XG16204 XI11_0/XI0/XI0_18/d_4_ XI11_0/XI0/XI0_18/d__4_ DECAP_INV_G11
XG16205 XI11_0/XI0/XI0_18/d_3_ XI11_0/XI0/XI0_18/d__3_ DECAP_INV_G11
XG16206 XI11_0/XI0/XI0_18/d_2_ XI11_0/XI0/XI0_18/d__2_ DECAP_INV_G11
XG16207 XI11_0/XI0/XI0_18/d_1_ XI11_0/XI0/XI0_18/d__1_ DECAP_INV_G11
XG16208 XI11_0/XI0/XI0_18/d_0_ XI11_0/XI0/XI0_18/d__0_ DECAP_INV_G11
XG16209 XI11_0/XI0/XI0_17/d__15_ XI11_0/XI0/XI0_17/d_15_ DECAP_INV_G11
XG16210 XI11_0/XI0/XI0_17/d__14_ XI11_0/XI0/XI0_17/d_14_ DECAP_INV_G11
XG16211 XI11_0/XI0/XI0_17/d__13_ XI11_0/XI0/XI0_17/d_13_ DECAP_INV_G11
XG16212 XI11_0/XI0/XI0_17/d__12_ XI11_0/XI0/XI0_17/d_12_ DECAP_INV_G11
XG16213 XI11_0/XI0/XI0_17/d__11_ XI11_0/XI0/XI0_17/d_11_ DECAP_INV_G11
XG16214 XI11_0/XI0/XI0_17/d__10_ XI11_0/XI0/XI0_17/d_10_ DECAP_INV_G11
XG16215 XI11_0/XI0/XI0_17/d__9_ XI11_0/XI0/XI0_17/d_9_ DECAP_INV_G11
XG16216 XI11_0/XI0/XI0_17/d__8_ XI11_0/XI0/XI0_17/d_8_ DECAP_INV_G11
XG16217 XI11_0/XI0/XI0_17/d__7_ XI11_0/XI0/XI0_17/d_7_ DECAP_INV_G11
XG16218 XI11_0/XI0/XI0_17/d__6_ XI11_0/XI0/XI0_17/d_6_ DECAP_INV_G11
XG16219 XI11_0/XI0/XI0_17/d__5_ XI11_0/XI0/XI0_17/d_5_ DECAP_INV_G11
XG16220 XI11_0/XI0/XI0_17/d__4_ XI11_0/XI0/XI0_17/d_4_ DECAP_INV_G11
XG16221 XI11_0/XI0/XI0_17/d__3_ XI11_0/XI0/XI0_17/d_3_ DECAP_INV_G11
XG16222 XI11_0/XI0/XI0_17/d__2_ XI11_0/XI0/XI0_17/d_2_ DECAP_INV_G11
XG16223 XI11_0/XI0/XI0_17/d__1_ XI11_0/XI0/XI0_17/d_1_ DECAP_INV_G11
XG16224 XI11_0/XI0/XI0_17/d__0_ XI11_0/XI0/XI0_17/d_0_ DECAP_INV_G11
XG16225 XI11_0/XI0/XI0_17/d_15_ XI11_0/XI0/XI0_17/d__15_ DECAP_INV_G11
XG16226 XI11_0/XI0/XI0_17/d_14_ XI11_0/XI0/XI0_17/d__14_ DECAP_INV_G11
XG16227 XI11_0/XI0/XI0_17/d_13_ XI11_0/XI0/XI0_17/d__13_ DECAP_INV_G11
XG16228 XI11_0/XI0/XI0_17/d_12_ XI11_0/XI0/XI0_17/d__12_ DECAP_INV_G11
XG16229 XI11_0/XI0/XI0_17/d_11_ XI11_0/XI0/XI0_17/d__11_ DECAP_INV_G11
XG16230 XI11_0/XI0/XI0_17/d_10_ XI11_0/XI0/XI0_17/d__10_ DECAP_INV_G11
XG16231 XI11_0/XI0/XI0_17/d_9_ XI11_0/XI0/XI0_17/d__9_ DECAP_INV_G11
XG16232 XI11_0/XI0/XI0_17/d_8_ XI11_0/XI0/XI0_17/d__8_ DECAP_INV_G11
XG16233 XI11_0/XI0/XI0_17/d_7_ XI11_0/XI0/XI0_17/d__7_ DECAP_INV_G11
XG16234 XI11_0/XI0/XI0_17/d_6_ XI11_0/XI0/XI0_17/d__6_ DECAP_INV_G11
XG16235 XI11_0/XI0/XI0_17/d_5_ XI11_0/XI0/XI0_17/d__5_ DECAP_INV_G11
XG16236 XI11_0/XI0/XI0_17/d_4_ XI11_0/XI0/XI0_17/d__4_ DECAP_INV_G11
XG16237 XI11_0/XI0/XI0_17/d_3_ XI11_0/XI0/XI0_17/d__3_ DECAP_INV_G11
XG16238 XI11_0/XI0/XI0_17/d_2_ XI11_0/XI0/XI0_17/d__2_ DECAP_INV_G11
XG16239 XI11_0/XI0/XI0_17/d_1_ XI11_0/XI0/XI0_17/d__1_ DECAP_INV_G11
XG16240 XI11_0/XI0/XI0_17/d_0_ XI11_0/XI0/XI0_17/d__0_ DECAP_INV_G11
XG16241 XI11_0/XI0/XI0_16/d__15_ XI11_0/XI0/XI0_16/d_15_ DECAP_INV_G11
XG16242 XI11_0/XI0/XI0_16/d__14_ XI11_0/XI0/XI0_16/d_14_ DECAP_INV_G11
XG16243 XI11_0/XI0/XI0_16/d__13_ XI11_0/XI0/XI0_16/d_13_ DECAP_INV_G11
XG16244 XI11_0/XI0/XI0_16/d__12_ XI11_0/XI0/XI0_16/d_12_ DECAP_INV_G11
XG16245 XI11_0/XI0/XI0_16/d__11_ XI11_0/XI0/XI0_16/d_11_ DECAP_INV_G11
XG16246 XI11_0/XI0/XI0_16/d__10_ XI11_0/XI0/XI0_16/d_10_ DECAP_INV_G11
XG16247 XI11_0/XI0/XI0_16/d__9_ XI11_0/XI0/XI0_16/d_9_ DECAP_INV_G11
XG16248 XI11_0/XI0/XI0_16/d__8_ XI11_0/XI0/XI0_16/d_8_ DECAP_INV_G11
XG16249 XI11_0/XI0/XI0_16/d__7_ XI11_0/XI0/XI0_16/d_7_ DECAP_INV_G11
XG16250 XI11_0/XI0/XI0_16/d__6_ XI11_0/XI0/XI0_16/d_6_ DECAP_INV_G11
XG16251 XI11_0/XI0/XI0_16/d__5_ XI11_0/XI0/XI0_16/d_5_ DECAP_INV_G11
XG16252 XI11_0/XI0/XI0_16/d__4_ XI11_0/XI0/XI0_16/d_4_ DECAP_INV_G11
XG16253 XI11_0/XI0/XI0_16/d__3_ XI11_0/XI0/XI0_16/d_3_ DECAP_INV_G11
XG16254 XI11_0/XI0/XI0_16/d__2_ XI11_0/XI0/XI0_16/d_2_ DECAP_INV_G11
XG16255 XI11_0/XI0/XI0_16/d__1_ XI11_0/XI0/XI0_16/d_1_ DECAP_INV_G11
XG16256 XI11_0/XI0/XI0_16/d__0_ XI11_0/XI0/XI0_16/d_0_ DECAP_INV_G11
XG16257 XI11_0/XI0/XI0_16/d_15_ XI11_0/XI0/XI0_16/d__15_ DECAP_INV_G11
XG16258 XI11_0/XI0/XI0_16/d_14_ XI11_0/XI0/XI0_16/d__14_ DECAP_INV_G11
XG16259 XI11_0/XI0/XI0_16/d_13_ XI11_0/XI0/XI0_16/d__13_ DECAP_INV_G11
XG16260 XI11_0/XI0/XI0_16/d_12_ XI11_0/XI0/XI0_16/d__12_ DECAP_INV_G11
XG16261 XI11_0/XI0/XI0_16/d_11_ XI11_0/XI0/XI0_16/d__11_ DECAP_INV_G11
XG16262 XI11_0/XI0/XI0_16/d_10_ XI11_0/XI0/XI0_16/d__10_ DECAP_INV_G11
XG16263 XI11_0/XI0/XI0_16/d_9_ XI11_0/XI0/XI0_16/d__9_ DECAP_INV_G11
XG16264 XI11_0/XI0/XI0_16/d_8_ XI11_0/XI0/XI0_16/d__8_ DECAP_INV_G11
XG16265 XI11_0/XI0/XI0_16/d_7_ XI11_0/XI0/XI0_16/d__7_ DECAP_INV_G11
XG16266 XI11_0/XI0/XI0_16/d_6_ XI11_0/XI0/XI0_16/d__6_ DECAP_INV_G11
XG16267 XI11_0/XI0/XI0_16/d_5_ XI11_0/XI0/XI0_16/d__5_ DECAP_INV_G11
XG16268 XI11_0/XI0/XI0_16/d_4_ XI11_0/XI0/XI0_16/d__4_ DECAP_INV_G11
XG16269 XI11_0/XI0/XI0_16/d_3_ XI11_0/XI0/XI0_16/d__3_ DECAP_INV_G11
XG16270 XI11_0/XI0/XI0_16/d_2_ XI11_0/XI0/XI0_16/d__2_ DECAP_INV_G11
XG16271 XI11_0/XI0/XI0_16/d_1_ XI11_0/XI0/XI0_16/d__1_ DECAP_INV_G11
XG16272 XI11_0/XI0/XI0_16/d_0_ XI11_0/XI0/XI0_16/d__0_ DECAP_INV_G11
XG16273 XI11_0/XI0/XI0_15/d__15_ XI11_0/XI0/XI0_15/d_15_ DECAP_INV_G11
XG16274 XI11_0/XI0/XI0_15/d__14_ XI11_0/XI0/XI0_15/d_14_ DECAP_INV_G11
XG16275 XI11_0/XI0/XI0_15/d__13_ XI11_0/XI0/XI0_15/d_13_ DECAP_INV_G11
XG16276 XI11_0/XI0/XI0_15/d__12_ XI11_0/XI0/XI0_15/d_12_ DECAP_INV_G11
XG16277 XI11_0/XI0/XI0_15/d__11_ XI11_0/XI0/XI0_15/d_11_ DECAP_INV_G11
XG16278 XI11_0/XI0/XI0_15/d__10_ XI11_0/XI0/XI0_15/d_10_ DECAP_INV_G11
XG16279 XI11_0/XI0/XI0_15/d__9_ XI11_0/XI0/XI0_15/d_9_ DECAP_INV_G11
XG16280 XI11_0/XI0/XI0_15/d__8_ XI11_0/XI0/XI0_15/d_8_ DECAP_INV_G11
XG16281 XI11_0/XI0/XI0_15/d__7_ XI11_0/XI0/XI0_15/d_7_ DECAP_INV_G11
XG16282 XI11_0/XI0/XI0_15/d__6_ XI11_0/XI0/XI0_15/d_6_ DECAP_INV_G11
XG16283 XI11_0/XI0/XI0_15/d__5_ XI11_0/XI0/XI0_15/d_5_ DECAP_INV_G11
XG16284 XI11_0/XI0/XI0_15/d__4_ XI11_0/XI0/XI0_15/d_4_ DECAP_INV_G11
XG16285 XI11_0/XI0/XI0_15/d__3_ XI11_0/XI0/XI0_15/d_3_ DECAP_INV_G11
XG16286 XI11_0/XI0/XI0_15/d__2_ XI11_0/XI0/XI0_15/d_2_ DECAP_INV_G11
XG16287 XI11_0/XI0/XI0_15/d__1_ XI11_0/XI0/XI0_15/d_1_ DECAP_INV_G11
XG16288 XI11_0/XI0/XI0_15/d__0_ XI11_0/XI0/XI0_15/d_0_ DECAP_INV_G11
XG16289 XI11_0/XI0/XI0_15/d_15_ XI11_0/XI0/XI0_15/d__15_ DECAP_INV_G11
XG16290 XI11_0/XI0/XI0_15/d_14_ XI11_0/XI0/XI0_15/d__14_ DECAP_INV_G11
XG16291 XI11_0/XI0/XI0_15/d_13_ XI11_0/XI0/XI0_15/d__13_ DECAP_INV_G11
XG16292 XI11_0/XI0/XI0_15/d_12_ XI11_0/XI0/XI0_15/d__12_ DECAP_INV_G11
XG16293 XI11_0/XI0/XI0_15/d_11_ XI11_0/XI0/XI0_15/d__11_ DECAP_INV_G11
XG16294 XI11_0/XI0/XI0_15/d_10_ XI11_0/XI0/XI0_15/d__10_ DECAP_INV_G11
XG16295 XI11_0/XI0/XI0_15/d_9_ XI11_0/XI0/XI0_15/d__9_ DECAP_INV_G11
XG16296 XI11_0/XI0/XI0_15/d_8_ XI11_0/XI0/XI0_15/d__8_ DECAP_INV_G11
XG16297 XI11_0/XI0/XI0_15/d_7_ XI11_0/XI0/XI0_15/d__7_ DECAP_INV_G11
XG16298 XI11_0/XI0/XI0_15/d_6_ XI11_0/XI0/XI0_15/d__6_ DECAP_INV_G11
XG16299 XI11_0/XI0/XI0_15/d_5_ XI11_0/XI0/XI0_15/d__5_ DECAP_INV_G11
XG16300 XI11_0/XI0/XI0_15/d_4_ XI11_0/XI0/XI0_15/d__4_ DECAP_INV_G11
XG16301 XI11_0/XI0/XI0_15/d_3_ XI11_0/XI0/XI0_15/d__3_ DECAP_INV_G11
XG16302 XI11_0/XI0/XI0_15/d_2_ XI11_0/XI0/XI0_15/d__2_ DECAP_INV_G11
XG16303 XI11_0/XI0/XI0_15/d_1_ XI11_0/XI0/XI0_15/d__1_ DECAP_INV_G11
XG16304 XI11_0/XI0/XI0_15/d_0_ XI11_0/XI0/XI0_15/d__0_ DECAP_INV_G11
XG16305 XI11_0/XI0/XI0_14/d__15_ XI11_0/XI0/XI0_14/d_15_ DECAP_INV_G11
XG16306 XI11_0/XI0/XI0_14/d__14_ XI11_0/XI0/XI0_14/d_14_ DECAP_INV_G11
XG16307 XI11_0/XI0/XI0_14/d__13_ XI11_0/XI0/XI0_14/d_13_ DECAP_INV_G11
XG16308 XI11_0/XI0/XI0_14/d__12_ XI11_0/XI0/XI0_14/d_12_ DECAP_INV_G11
XG16309 XI11_0/XI0/XI0_14/d__11_ XI11_0/XI0/XI0_14/d_11_ DECAP_INV_G11
XG16310 XI11_0/XI0/XI0_14/d__10_ XI11_0/XI0/XI0_14/d_10_ DECAP_INV_G11
XG16311 XI11_0/XI0/XI0_14/d__9_ XI11_0/XI0/XI0_14/d_9_ DECAP_INV_G11
XG16312 XI11_0/XI0/XI0_14/d__8_ XI11_0/XI0/XI0_14/d_8_ DECAP_INV_G11
XG16313 XI11_0/XI0/XI0_14/d__7_ XI11_0/XI0/XI0_14/d_7_ DECAP_INV_G11
XG16314 XI11_0/XI0/XI0_14/d__6_ XI11_0/XI0/XI0_14/d_6_ DECAP_INV_G11
XG16315 XI11_0/XI0/XI0_14/d__5_ XI11_0/XI0/XI0_14/d_5_ DECAP_INV_G11
XG16316 XI11_0/XI0/XI0_14/d__4_ XI11_0/XI0/XI0_14/d_4_ DECAP_INV_G11
XG16317 XI11_0/XI0/XI0_14/d__3_ XI11_0/XI0/XI0_14/d_3_ DECAP_INV_G11
XG16318 XI11_0/XI0/XI0_14/d__2_ XI11_0/XI0/XI0_14/d_2_ DECAP_INV_G11
XG16319 XI11_0/XI0/XI0_14/d__1_ XI11_0/XI0/XI0_14/d_1_ DECAP_INV_G11
XG16320 XI11_0/XI0/XI0_14/d__0_ XI11_0/XI0/XI0_14/d_0_ DECAP_INV_G11
XG16321 XI11_0/XI0/XI0_14/d_15_ XI11_0/XI0/XI0_14/d__15_ DECAP_INV_G11
XG16322 XI11_0/XI0/XI0_14/d_14_ XI11_0/XI0/XI0_14/d__14_ DECAP_INV_G11
XG16323 XI11_0/XI0/XI0_14/d_13_ XI11_0/XI0/XI0_14/d__13_ DECAP_INV_G11
XG16324 XI11_0/XI0/XI0_14/d_12_ XI11_0/XI0/XI0_14/d__12_ DECAP_INV_G11
XG16325 XI11_0/XI0/XI0_14/d_11_ XI11_0/XI0/XI0_14/d__11_ DECAP_INV_G11
XG16326 XI11_0/XI0/XI0_14/d_10_ XI11_0/XI0/XI0_14/d__10_ DECAP_INV_G11
XG16327 XI11_0/XI0/XI0_14/d_9_ XI11_0/XI0/XI0_14/d__9_ DECAP_INV_G11
XG16328 XI11_0/XI0/XI0_14/d_8_ XI11_0/XI0/XI0_14/d__8_ DECAP_INV_G11
XG16329 XI11_0/XI0/XI0_14/d_7_ XI11_0/XI0/XI0_14/d__7_ DECAP_INV_G11
XG16330 XI11_0/XI0/XI0_14/d_6_ XI11_0/XI0/XI0_14/d__6_ DECAP_INV_G11
XG16331 XI11_0/XI0/XI0_14/d_5_ XI11_0/XI0/XI0_14/d__5_ DECAP_INV_G11
XG16332 XI11_0/XI0/XI0_14/d_4_ XI11_0/XI0/XI0_14/d__4_ DECAP_INV_G11
XG16333 XI11_0/XI0/XI0_14/d_3_ XI11_0/XI0/XI0_14/d__3_ DECAP_INV_G11
XG16334 XI11_0/XI0/XI0_14/d_2_ XI11_0/XI0/XI0_14/d__2_ DECAP_INV_G11
XG16335 XI11_0/XI0/XI0_14/d_1_ XI11_0/XI0/XI0_14/d__1_ DECAP_INV_G11
XG16336 XI11_0/XI0/XI0_14/d_0_ XI11_0/XI0/XI0_14/d__0_ DECAP_INV_G11
XG16337 XI11_0/XI0/XI0_13/d__15_ XI11_0/XI0/XI0_13/d_15_ DECAP_INV_G11
XG16338 XI11_0/XI0/XI0_13/d__14_ XI11_0/XI0/XI0_13/d_14_ DECAP_INV_G11
XG16339 XI11_0/XI0/XI0_13/d__13_ XI11_0/XI0/XI0_13/d_13_ DECAP_INV_G11
XG16340 XI11_0/XI0/XI0_13/d__12_ XI11_0/XI0/XI0_13/d_12_ DECAP_INV_G11
XG16341 XI11_0/XI0/XI0_13/d__11_ XI11_0/XI0/XI0_13/d_11_ DECAP_INV_G11
XG16342 XI11_0/XI0/XI0_13/d__10_ XI11_0/XI0/XI0_13/d_10_ DECAP_INV_G11
XG16343 XI11_0/XI0/XI0_13/d__9_ XI11_0/XI0/XI0_13/d_9_ DECAP_INV_G11
XG16344 XI11_0/XI0/XI0_13/d__8_ XI11_0/XI0/XI0_13/d_8_ DECAP_INV_G11
XG16345 XI11_0/XI0/XI0_13/d__7_ XI11_0/XI0/XI0_13/d_7_ DECAP_INV_G11
XG16346 XI11_0/XI0/XI0_13/d__6_ XI11_0/XI0/XI0_13/d_6_ DECAP_INV_G11
XG16347 XI11_0/XI0/XI0_13/d__5_ XI11_0/XI0/XI0_13/d_5_ DECAP_INV_G11
XG16348 XI11_0/XI0/XI0_13/d__4_ XI11_0/XI0/XI0_13/d_4_ DECAP_INV_G11
XG16349 XI11_0/XI0/XI0_13/d__3_ XI11_0/XI0/XI0_13/d_3_ DECAP_INV_G11
XG16350 XI11_0/XI0/XI0_13/d__2_ XI11_0/XI0/XI0_13/d_2_ DECAP_INV_G11
XG16351 XI11_0/XI0/XI0_13/d__1_ XI11_0/XI0/XI0_13/d_1_ DECAP_INV_G11
XG16352 XI11_0/XI0/XI0_13/d__0_ XI11_0/XI0/XI0_13/d_0_ DECAP_INV_G11
XG16353 XI11_0/XI0/XI0_13/d_15_ XI11_0/XI0/XI0_13/d__15_ DECAP_INV_G11
XG16354 XI11_0/XI0/XI0_13/d_14_ XI11_0/XI0/XI0_13/d__14_ DECAP_INV_G11
XG16355 XI11_0/XI0/XI0_13/d_13_ XI11_0/XI0/XI0_13/d__13_ DECAP_INV_G11
XG16356 XI11_0/XI0/XI0_13/d_12_ XI11_0/XI0/XI0_13/d__12_ DECAP_INV_G11
XG16357 XI11_0/XI0/XI0_13/d_11_ XI11_0/XI0/XI0_13/d__11_ DECAP_INV_G11
XG16358 XI11_0/XI0/XI0_13/d_10_ XI11_0/XI0/XI0_13/d__10_ DECAP_INV_G11
XG16359 XI11_0/XI0/XI0_13/d_9_ XI11_0/XI0/XI0_13/d__9_ DECAP_INV_G11
XG16360 XI11_0/XI0/XI0_13/d_8_ XI11_0/XI0/XI0_13/d__8_ DECAP_INV_G11
XG16361 XI11_0/XI0/XI0_13/d_7_ XI11_0/XI0/XI0_13/d__7_ DECAP_INV_G11
XG16362 XI11_0/XI0/XI0_13/d_6_ XI11_0/XI0/XI0_13/d__6_ DECAP_INV_G11
XG16363 XI11_0/XI0/XI0_13/d_5_ XI11_0/XI0/XI0_13/d__5_ DECAP_INV_G11
XG16364 XI11_0/XI0/XI0_13/d_4_ XI11_0/XI0/XI0_13/d__4_ DECAP_INV_G11
XG16365 XI11_0/XI0/XI0_13/d_3_ XI11_0/XI0/XI0_13/d__3_ DECAP_INV_G11
XG16366 XI11_0/XI0/XI0_13/d_2_ XI11_0/XI0/XI0_13/d__2_ DECAP_INV_G11
XG16367 XI11_0/XI0/XI0_13/d_1_ XI11_0/XI0/XI0_13/d__1_ DECAP_INV_G11
XG16368 XI11_0/XI0/XI0_13/d_0_ XI11_0/XI0/XI0_13/d__0_ DECAP_INV_G11
XG16369 XI11_0/XI0/XI0_12/d__15_ XI11_0/XI0/XI0_12/d_15_ DECAP_INV_G11
XG16370 XI11_0/XI0/XI0_12/d__14_ XI11_0/XI0/XI0_12/d_14_ DECAP_INV_G11
XG16371 XI11_0/XI0/XI0_12/d__13_ XI11_0/XI0/XI0_12/d_13_ DECAP_INV_G11
XG16372 XI11_0/XI0/XI0_12/d__12_ XI11_0/XI0/XI0_12/d_12_ DECAP_INV_G11
XG16373 XI11_0/XI0/XI0_12/d__11_ XI11_0/XI0/XI0_12/d_11_ DECAP_INV_G11
XG16374 XI11_0/XI0/XI0_12/d__10_ XI11_0/XI0/XI0_12/d_10_ DECAP_INV_G11
XG16375 XI11_0/XI0/XI0_12/d__9_ XI11_0/XI0/XI0_12/d_9_ DECAP_INV_G11
XG16376 XI11_0/XI0/XI0_12/d__8_ XI11_0/XI0/XI0_12/d_8_ DECAP_INV_G11
XG16377 XI11_0/XI0/XI0_12/d__7_ XI11_0/XI0/XI0_12/d_7_ DECAP_INV_G11
XG16378 XI11_0/XI0/XI0_12/d__6_ XI11_0/XI0/XI0_12/d_6_ DECAP_INV_G11
XG16379 XI11_0/XI0/XI0_12/d__5_ XI11_0/XI0/XI0_12/d_5_ DECAP_INV_G11
XG16380 XI11_0/XI0/XI0_12/d__4_ XI11_0/XI0/XI0_12/d_4_ DECAP_INV_G11
XG16381 XI11_0/XI0/XI0_12/d__3_ XI11_0/XI0/XI0_12/d_3_ DECAP_INV_G11
XG16382 XI11_0/XI0/XI0_12/d__2_ XI11_0/XI0/XI0_12/d_2_ DECAP_INV_G11
XG16383 XI11_0/XI0/XI0_12/d__1_ XI11_0/XI0/XI0_12/d_1_ DECAP_INV_G11
XG16384 XI11_0/XI0/XI0_12/d__0_ XI11_0/XI0/XI0_12/d_0_ DECAP_INV_G11
XG16385 XI11_0/XI0/XI0_12/d_15_ XI11_0/XI0/XI0_12/d__15_ DECAP_INV_G11
XG16386 XI11_0/XI0/XI0_12/d_14_ XI11_0/XI0/XI0_12/d__14_ DECAP_INV_G11
XG16387 XI11_0/XI0/XI0_12/d_13_ XI11_0/XI0/XI0_12/d__13_ DECAP_INV_G11
XG16388 XI11_0/XI0/XI0_12/d_12_ XI11_0/XI0/XI0_12/d__12_ DECAP_INV_G11
XG16389 XI11_0/XI0/XI0_12/d_11_ XI11_0/XI0/XI0_12/d__11_ DECAP_INV_G11
XG16390 XI11_0/XI0/XI0_12/d_10_ XI11_0/XI0/XI0_12/d__10_ DECAP_INV_G11
XG16391 XI11_0/XI0/XI0_12/d_9_ XI11_0/XI0/XI0_12/d__9_ DECAP_INV_G11
XG16392 XI11_0/XI0/XI0_12/d_8_ XI11_0/XI0/XI0_12/d__8_ DECAP_INV_G11
XG16393 XI11_0/XI0/XI0_12/d_7_ XI11_0/XI0/XI0_12/d__7_ DECAP_INV_G11
XG16394 XI11_0/XI0/XI0_12/d_6_ XI11_0/XI0/XI0_12/d__6_ DECAP_INV_G11
XG16395 XI11_0/XI0/XI0_12/d_5_ XI11_0/XI0/XI0_12/d__5_ DECAP_INV_G11
XG16396 XI11_0/XI0/XI0_12/d_4_ XI11_0/XI0/XI0_12/d__4_ DECAP_INV_G11
XG16397 XI11_0/XI0/XI0_12/d_3_ XI11_0/XI0/XI0_12/d__3_ DECAP_INV_G11
XG16398 XI11_0/XI0/XI0_12/d_2_ XI11_0/XI0/XI0_12/d__2_ DECAP_INV_G11
XG16399 XI11_0/XI0/XI0_12/d_1_ XI11_0/XI0/XI0_12/d__1_ DECAP_INV_G11
XG16400 XI11_0/XI0/XI0_12/d_0_ XI11_0/XI0/XI0_12/d__0_ DECAP_INV_G11
XG16401 XI11_0/XI0/XI0_11/d__15_ XI11_0/XI0/XI0_11/d_15_ DECAP_INV_G11
XG16402 XI11_0/XI0/XI0_11/d__14_ XI11_0/XI0/XI0_11/d_14_ DECAP_INV_G11
XG16403 XI11_0/XI0/XI0_11/d__13_ XI11_0/XI0/XI0_11/d_13_ DECAP_INV_G11
XG16404 XI11_0/XI0/XI0_11/d__12_ XI11_0/XI0/XI0_11/d_12_ DECAP_INV_G11
XG16405 XI11_0/XI0/XI0_11/d__11_ XI11_0/XI0/XI0_11/d_11_ DECAP_INV_G11
XG16406 XI11_0/XI0/XI0_11/d__10_ XI11_0/XI0/XI0_11/d_10_ DECAP_INV_G11
XG16407 XI11_0/XI0/XI0_11/d__9_ XI11_0/XI0/XI0_11/d_9_ DECAP_INV_G11
XG16408 XI11_0/XI0/XI0_11/d__8_ XI11_0/XI0/XI0_11/d_8_ DECAP_INV_G11
XG16409 XI11_0/XI0/XI0_11/d__7_ XI11_0/XI0/XI0_11/d_7_ DECAP_INV_G11
XG16410 XI11_0/XI0/XI0_11/d__6_ XI11_0/XI0/XI0_11/d_6_ DECAP_INV_G11
XG16411 XI11_0/XI0/XI0_11/d__5_ XI11_0/XI0/XI0_11/d_5_ DECAP_INV_G11
XG16412 XI11_0/XI0/XI0_11/d__4_ XI11_0/XI0/XI0_11/d_4_ DECAP_INV_G11
XG16413 XI11_0/XI0/XI0_11/d__3_ XI11_0/XI0/XI0_11/d_3_ DECAP_INV_G11
XG16414 XI11_0/XI0/XI0_11/d__2_ XI11_0/XI0/XI0_11/d_2_ DECAP_INV_G11
XG16415 XI11_0/XI0/XI0_11/d__1_ XI11_0/XI0/XI0_11/d_1_ DECAP_INV_G11
XG16416 XI11_0/XI0/XI0_11/d__0_ XI11_0/XI0/XI0_11/d_0_ DECAP_INV_G11
XG16417 XI11_0/XI0/XI0_11/d_15_ XI11_0/XI0/XI0_11/d__15_ DECAP_INV_G11
XG16418 XI11_0/XI0/XI0_11/d_14_ XI11_0/XI0/XI0_11/d__14_ DECAP_INV_G11
XG16419 XI11_0/XI0/XI0_11/d_13_ XI11_0/XI0/XI0_11/d__13_ DECAP_INV_G11
XG16420 XI11_0/XI0/XI0_11/d_12_ XI11_0/XI0/XI0_11/d__12_ DECAP_INV_G11
XG16421 XI11_0/XI0/XI0_11/d_11_ XI11_0/XI0/XI0_11/d__11_ DECAP_INV_G11
XG16422 XI11_0/XI0/XI0_11/d_10_ XI11_0/XI0/XI0_11/d__10_ DECAP_INV_G11
XG16423 XI11_0/XI0/XI0_11/d_9_ XI11_0/XI0/XI0_11/d__9_ DECAP_INV_G11
XG16424 XI11_0/XI0/XI0_11/d_8_ XI11_0/XI0/XI0_11/d__8_ DECAP_INV_G11
XG16425 XI11_0/XI0/XI0_11/d_7_ XI11_0/XI0/XI0_11/d__7_ DECAP_INV_G11
XG16426 XI11_0/XI0/XI0_11/d_6_ XI11_0/XI0/XI0_11/d__6_ DECAP_INV_G11
XG16427 XI11_0/XI0/XI0_11/d_5_ XI11_0/XI0/XI0_11/d__5_ DECAP_INV_G11
XG16428 XI11_0/XI0/XI0_11/d_4_ XI11_0/XI0/XI0_11/d__4_ DECAP_INV_G11
XG16429 XI11_0/XI0/XI0_11/d_3_ XI11_0/XI0/XI0_11/d__3_ DECAP_INV_G11
XG16430 XI11_0/XI0/XI0_11/d_2_ XI11_0/XI0/XI0_11/d__2_ DECAP_INV_G11
XG16431 XI11_0/XI0/XI0_11/d_1_ XI11_0/XI0/XI0_11/d__1_ DECAP_INV_G11
XG16432 XI11_0/XI0/XI0_11/d_0_ XI11_0/XI0/XI0_11/d__0_ DECAP_INV_G11
XG16433 XI11_0/XI0/XI0_10/d__15_ XI11_0/XI0/XI0_10/d_15_ DECAP_INV_G11
XG16434 XI11_0/XI0/XI0_10/d__14_ XI11_0/XI0/XI0_10/d_14_ DECAP_INV_G11
XG16435 XI11_0/XI0/XI0_10/d__13_ XI11_0/XI0/XI0_10/d_13_ DECAP_INV_G11
XG16436 XI11_0/XI0/XI0_10/d__12_ XI11_0/XI0/XI0_10/d_12_ DECAP_INV_G11
XG16437 XI11_0/XI0/XI0_10/d__11_ XI11_0/XI0/XI0_10/d_11_ DECAP_INV_G11
XG16438 XI11_0/XI0/XI0_10/d__10_ XI11_0/XI0/XI0_10/d_10_ DECAP_INV_G11
XG16439 XI11_0/XI0/XI0_10/d__9_ XI11_0/XI0/XI0_10/d_9_ DECAP_INV_G11
XG16440 XI11_0/XI0/XI0_10/d__8_ XI11_0/XI0/XI0_10/d_8_ DECAP_INV_G11
XG16441 XI11_0/XI0/XI0_10/d__7_ XI11_0/XI0/XI0_10/d_7_ DECAP_INV_G11
XG16442 XI11_0/XI0/XI0_10/d__6_ XI11_0/XI0/XI0_10/d_6_ DECAP_INV_G11
XG16443 XI11_0/XI0/XI0_10/d__5_ XI11_0/XI0/XI0_10/d_5_ DECAP_INV_G11
XG16444 XI11_0/XI0/XI0_10/d__4_ XI11_0/XI0/XI0_10/d_4_ DECAP_INV_G11
XG16445 XI11_0/XI0/XI0_10/d__3_ XI11_0/XI0/XI0_10/d_3_ DECAP_INV_G11
XG16446 XI11_0/XI0/XI0_10/d__2_ XI11_0/XI0/XI0_10/d_2_ DECAP_INV_G11
XG16447 XI11_0/XI0/XI0_10/d__1_ XI11_0/XI0/XI0_10/d_1_ DECAP_INV_G11
XG16448 XI11_0/XI0/XI0_10/d__0_ XI11_0/XI0/XI0_10/d_0_ DECAP_INV_G11
XG16449 XI11_0/XI0/XI0_10/d_15_ XI11_0/XI0/XI0_10/d__15_ DECAP_INV_G11
XG16450 XI11_0/XI0/XI0_10/d_14_ XI11_0/XI0/XI0_10/d__14_ DECAP_INV_G11
XG16451 XI11_0/XI0/XI0_10/d_13_ XI11_0/XI0/XI0_10/d__13_ DECAP_INV_G11
XG16452 XI11_0/XI0/XI0_10/d_12_ XI11_0/XI0/XI0_10/d__12_ DECAP_INV_G11
XG16453 XI11_0/XI0/XI0_10/d_11_ XI11_0/XI0/XI0_10/d__11_ DECAP_INV_G11
XG16454 XI11_0/XI0/XI0_10/d_10_ XI11_0/XI0/XI0_10/d__10_ DECAP_INV_G11
XG16455 XI11_0/XI0/XI0_10/d_9_ XI11_0/XI0/XI0_10/d__9_ DECAP_INV_G11
XG16456 XI11_0/XI0/XI0_10/d_8_ XI11_0/XI0/XI0_10/d__8_ DECAP_INV_G11
XG16457 XI11_0/XI0/XI0_10/d_7_ XI11_0/XI0/XI0_10/d__7_ DECAP_INV_G11
XG16458 XI11_0/XI0/XI0_10/d_6_ XI11_0/XI0/XI0_10/d__6_ DECAP_INV_G11
XG16459 XI11_0/XI0/XI0_10/d_5_ XI11_0/XI0/XI0_10/d__5_ DECAP_INV_G11
XG16460 XI11_0/XI0/XI0_10/d_4_ XI11_0/XI0/XI0_10/d__4_ DECAP_INV_G11
XG16461 XI11_0/XI0/XI0_10/d_3_ XI11_0/XI0/XI0_10/d__3_ DECAP_INV_G11
XG16462 XI11_0/XI0/XI0_10/d_2_ XI11_0/XI0/XI0_10/d__2_ DECAP_INV_G11
XG16463 XI11_0/XI0/XI0_10/d_1_ XI11_0/XI0/XI0_10/d__1_ DECAP_INV_G11
XG16464 XI11_0/XI0/XI0_10/d_0_ XI11_0/XI0/XI0_10/d__0_ DECAP_INV_G11
XG16465 XI11_0/XI0/XI0_9/d__15_ XI11_0/XI0/XI0_9/d_15_ DECAP_INV_G11
XG16466 XI11_0/XI0/XI0_9/d__14_ XI11_0/XI0/XI0_9/d_14_ DECAP_INV_G11
XG16467 XI11_0/XI0/XI0_9/d__13_ XI11_0/XI0/XI0_9/d_13_ DECAP_INV_G11
XG16468 XI11_0/XI0/XI0_9/d__12_ XI11_0/XI0/XI0_9/d_12_ DECAP_INV_G11
XG16469 XI11_0/XI0/XI0_9/d__11_ XI11_0/XI0/XI0_9/d_11_ DECAP_INV_G11
XG16470 XI11_0/XI0/XI0_9/d__10_ XI11_0/XI0/XI0_9/d_10_ DECAP_INV_G11
XG16471 XI11_0/XI0/XI0_9/d__9_ XI11_0/XI0/XI0_9/d_9_ DECAP_INV_G11
XG16472 XI11_0/XI0/XI0_9/d__8_ XI11_0/XI0/XI0_9/d_8_ DECAP_INV_G11
XG16473 XI11_0/XI0/XI0_9/d__7_ XI11_0/XI0/XI0_9/d_7_ DECAP_INV_G11
XG16474 XI11_0/XI0/XI0_9/d__6_ XI11_0/XI0/XI0_9/d_6_ DECAP_INV_G11
XG16475 XI11_0/XI0/XI0_9/d__5_ XI11_0/XI0/XI0_9/d_5_ DECAP_INV_G11
XG16476 XI11_0/XI0/XI0_9/d__4_ XI11_0/XI0/XI0_9/d_4_ DECAP_INV_G11
XG16477 XI11_0/XI0/XI0_9/d__3_ XI11_0/XI0/XI0_9/d_3_ DECAP_INV_G11
XG16478 XI11_0/XI0/XI0_9/d__2_ XI11_0/XI0/XI0_9/d_2_ DECAP_INV_G11
XG16479 XI11_0/XI0/XI0_9/d__1_ XI11_0/XI0/XI0_9/d_1_ DECAP_INV_G11
XG16480 XI11_0/XI0/XI0_9/d__0_ XI11_0/XI0/XI0_9/d_0_ DECAP_INV_G11
XG16481 XI11_0/XI0/XI0_9/d_15_ XI11_0/XI0/XI0_9/d__15_ DECAP_INV_G11
XG16482 XI11_0/XI0/XI0_9/d_14_ XI11_0/XI0/XI0_9/d__14_ DECAP_INV_G11
XG16483 XI11_0/XI0/XI0_9/d_13_ XI11_0/XI0/XI0_9/d__13_ DECAP_INV_G11
XG16484 XI11_0/XI0/XI0_9/d_12_ XI11_0/XI0/XI0_9/d__12_ DECAP_INV_G11
XG16485 XI11_0/XI0/XI0_9/d_11_ XI11_0/XI0/XI0_9/d__11_ DECAP_INV_G11
XG16486 XI11_0/XI0/XI0_9/d_10_ XI11_0/XI0/XI0_9/d__10_ DECAP_INV_G11
XG16487 XI11_0/XI0/XI0_9/d_9_ XI11_0/XI0/XI0_9/d__9_ DECAP_INV_G11
XG16488 XI11_0/XI0/XI0_9/d_8_ XI11_0/XI0/XI0_9/d__8_ DECAP_INV_G11
XG16489 XI11_0/XI0/XI0_9/d_7_ XI11_0/XI0/XI0_9/d__7_ DECAP_INV_G11
XG16490 XI11_0/XI0/XI0_9/d_6_ XI11_0/XI0/XI0_9/d__6_ DECAP_INV_G11
XG16491 XI11_0/XI0/XI0_9/d_5_ XI11_0/XI0/XI0_9/d__5_ DECAP_INV_G11
XG16492 XI11_0/XI0/XI0_9/d_4_ XI11_0/XI0/XI0_9/d__4_ DECAP_INV_G11
XG16493 XI11_0/XI0/XI0_9/d_3_ XI11_0/XI0/XI0_9/d__3_ DECAP_INV_G11
XG16494 XI11_0/XI0/XI0_9/d_2_ XI11_0/XI0/XI0_9/d__2_ DECAP_INV_G11
XG16495 XI11_0/XI0/XI0_9/d_1_ XI11_0/XI0/XI0_9/d__1_ DECAP_INV_G11
XG16496 XI11_0/XI0/XI0_9/d_0_ XI11_0/XI0/XI0_9/d__0_ DECAP_INV_G11
XG16497 XI11_0/XI0/XI0_8/d__15_ XI11_0/XI0/XI0_8/d_15_ DECAP_INV_G11
XG16498 XI11_0/XI0/XI0_8/d__14_ XI11_0/XI0/XI0_8/d_14_ DECAP_INV_G11
XG16499 XI11_0/XI0/XI0_8/d__13_ XI11_0/XI0/XI0_8/d_13_ DECAP_INV_G11
XG16500 XI11_0/XI0/XI0_8/d__12_ XI11_0/XI0/XI0_8/d_12_ DECAP_INV_G11
XG16501 XI11_0/XI0/XI0_8/d__11_ XI11_0/XI0/XI0_8/d_11_ DECAP_INV_G11
XG16502 XI11_0/XI0/XI0_8/d__10_ XI11_0/XI0/XI0_8/d_10_ DECAP_INV_G11
XG16503 XI11_0/XI0/XI0_8/d__9_ XI11_0/XI0/XI0_8/d_9_ DECAP_INV_G11
XG16504 XI11_0/XI0/XI0_8/d__8_ XI11_0/XI0/XI0_8/d_8_ DECAP_INV_G11
XG16505 XI11_0/XI0/XI0_8/d__7_ XI11_0/XI0/XI0_8/d_7_ DECAP_INV_G11
XG16506 XI11_0/XI0/XI0_8/d__6_ XI11_0/XI0/XI0_8/d_6_ DECAP_INV_G11
XG16507 XI11_0/XI0/XI0_8/d__5_ XI11_0/XI0/XI0_8/d_5_ DECAP_INV_G11
XG16508 XI11_0/XI0/XI0_8/d__4_ XI11_0/XI0/XI0_8/d_4_ DECAP_INV_G11
XG16509 XI11_0/XI0/XI0_8/d__3_ XI11_0/XI0/XI0_8/d_3_ DECAP_INV_G11
XG16510 XI11_0/XI0/XI0_8/d__2_ XI11_0/XI0/XI0_8/d_2_ DECAP_INV_G11
XG16511 XI11_0/XI0/XI0_8/d__1_ XI11_0/XI0/XI0_8/d_1_ DECAP_INV_G11
XG16512 XI11_0/XI0/XI0_8/d__0_ XI11_0/XI0/XI0_8/d_0_ DECAP_INV_G11
XG16513 XI11_0/XI0/XI0_8/d_15_ XI11_0/XI0/XI0_8/d__15_ DECAP_INV_G11
XG16514 XI11_0/XI0/XI0_8/d_14_ XI11_0/XI0/XI0_8/d__14_ DECAP_INV_G11
XG16515 XI11_0/XI0/XI0_8/d_13_ XI11_0/XI0/XI0_8/d__13_ DECAP_INV_G11
XG16516 XI11_0/XI0/XI0_8/d_12_ XI11_0/XI0/XI0_8/d__12_ DECAP_INV_G11
XG16517 XI11_0/XI0/XI0_8/d_11_ XI11_0/XI0/XI0_8/d__11_ DECAP_INV_G11
XG16518 XI11_0/XI0/XI0_8/d_10_ XI11_0/XI0/XI0_8/d__10_ DECAP_INV_G11
XG16519 XI11_0/XI0/XI0_8/d_9_ XI11_0/XI0/XI0_8/d__9_ DECAP_INV_G11
XG16520 XI11_0/XI0/XI0_8/d_8_ XI11_0/XI0/XI0_8/d__8_ DECAP_INV_G11
XG16521 XI11_0/XI0/XI0_8/d_7_ XI11_0/XI0/XI0_8/d__7_ DECAP_INV_G11
XG16522 XI11_0/XI0/XI0_8/d_6_ XI11_0/XI0/XI0_8/d__6_ DECAP_INV_G11
XG16523 XI11_0/XI0/XI0_8/d_5_ XI11_0/XI0/XI0_8/d__5_ DECAP_INV_G11
XG16524 XI11_0/XI0/XI0_8/d_4_ XI11_0/XI0/XI0_8/d__4_ DECAP_INV_G11
XG16525 XI11_0/XI0/XI0_8/d_3_ XI11_0/XI0/XI0_8/d__3_ DECAP_INV_G11
XG16526 XI11_0/XI0/XI0_8/d_2_ XI11_0/XI0/XI0_8/d__2_ DECAP_INV_G11
XG16527 XI11_0/XI0/XI0_8/d_1_ XI11_0/XI0/XI0_8/d__1_ DECAP_INV_G11
XG16528 XI11_0/XI0/XI0_8/d_0_ XI11_0/XI0/XI0_8/d__0_ DECAP_INV_G11
XG16529 XI11_0/XI0/XI0_7/d__15_ XI11_0/XI0/XI0_7/d_15_ DECAP_INV_G11
XG16530 XI11_0/XI0/XI0_7/d__14_ XI11_0/XI0/XI0_7/d_14_ DECAP_INV_G11
XG16531 XI11_0/XI0/XI0_7/d__13_ XI11_0/XI0/XI0_7/d_13_ DECAP_INV_G11
XG16532 XI11_0/XI0/XI0_7/d__12_ XI11_0/XI0/XI0_7/d_12_ DECAP_INV_G11
XG16533 XI11_0/XI0/XI0_7/d__11_ XI11_0/XI0/XI0_7/d_11_ DECAP_INV_G11
XG16534 XI11_0/XI0/XI0_7/d__10_ XI11_0/XI0/XI0_7/d_10_ DECAP_INV_G11
XG16535 XI11_0/XI0/XI0_7/d__9_ XI11_0/XI0/XI0_7/d_9_ DECAP_INV_G11
XG16536 XI11_0/XI0/XI0_7/d__8_ XI11_0/XI0/XI0_7/d_8_ DECAP_INV_G11
XG16537 XI11_0/XI0/XI0_7/d__7_ XI11_0/XI0/XI0_7/d_7_ DECAP_INV_G11
XG16538 XI11_0/XI0/XI0_7/d__6_ XI11_0/XI0/XI0_7/d_6_ DECAP_INV_G11
XG16539 XI11_0/XI0/XI0_7/d__5_ XI11_0/XI0/XI0_7/d_5_ DECAP_INV_G11
XG16540 XI11_0/XI0/XI0_7/d__4_ XI11_0/XI0/XI0_7/d_4_ DECAP_INV_G11
XG16541 XI11_0/XI0/XI0_7/d__3_ XI11_0/XI0/XI0_7/d_3_ DECAP_INV_G11
XG16542 XI11_0/XI0/XI0_7/d__2_ XI11_0/XI0/XI0_7/d_2_ DECAP_INV_G11
XG16543 XI11_0/XI0/XI0_7/d__1_ XI11_0/XI0/XI0_7/d_1_ DECAP_INV_G11
XG16544 XI11_0/XI0/XI0_7/d__0_ XI11_0/XI0/XI0_7/d_0_ DECAP_INV_G11
XG16545 XI11_0/XI0/XI0_7/d_15_ XI11_0/XI0/XI0_7/d__15_ DECAP_INV_G11
XG16546 XI11_0/XI0/XI0_7/d_14_ XI11_0/XI0/XI0_7/d__14_ DECAP_INV_G11
XG16547 XI11_0/XI0/XI0_7/d_13_ XI11_0/XI0/XI0_7/d__13_ DECAP_INV_G11
XG16548 XI11_0/XI0/XI0_7/d_12_ XI11_0/XI0/XI0_7/d__12_ DECAP_INV_G11
XG16549 XI11_0/XI0/XI0_7/d_11_ XI11_0/XI0/XI0_7/d__11_ DECAP_INV_G11
XG16550 XI11_0/XI0/XI0_7/d_10_ XI11_0/XI0/XI0_7/d__10_ DECAP_INV_G11
XG16551 XI11_0/XI0/XI0_7/d_9_ XI11_0/XI0/XI0_7/d__9_ DECAP_INV_G11
XG16552 XI11_0/XI0/XI0_7/d_8_ XI11_0/XI0/XI0_7/d__8_ DECAP_INV_G11
XG16553 XI11_0/XI0/XI0_7/d_7_ XI11_0/XI0/XI0_7/d__7_ DECAP_INV_G11
XG16554 XI11_0/XI0/XI0_7/d_6_ XI11_0/XI0/XI0_7/d__6_ DECAP_INV_G11
XG16555 XI11_0/XI0/XI0_7/d_5_ XI11_0/XI0/XI0_7/d__5_ DECAP_INV_G11
XG16556 XI11_0/XI0/XI0_7/d_4_ XI11_0/XI0/XI0_7/d__4_ DECAP_INV_G11
XG16557 XI11_0/XI0/XI0_7/d_3_ XI11_0/XI0/XI0_7/d__3_ DECAP_INV_G11
XG16558 XI11_0/XI0/XI0_7/d_2_ XI11_0/XI0/XI0_7/d__2_ DECAP_INV_G11
XG16559 XI11_0/XI0/XI0_7/d_1_ XI11_0/XI0/XI0_7/d__1_ DECAP_INV_G11
XG16560 XI11_0/XI0/XI0_7/d_0_ XI11_0/XI0/XI0_7/d__0_ DECAP_INV_G11
XG16561 XI11_0/XI0/XI0_6/d__15_ XI11_0/XI0/XI0_6/d_15_ DECAP_INV_G11
XG16562 XI11_0/XI0/XI0_6/d__14_ XI11_0/XI0/XI0_6/d_14_ DECAP_INV_G11
XG16563 XI11_0/XI0/XI0_6/d__13_ XI11_0/XI0/XI0_6/d_13_ DECAP_INV_G11
XG16564 XI11_0/XI0/XI0_6/d__12_ XI11_0/XI0/XI0_6/d_12_ DECAP_INV_G11
XG16565 XI11_0/XI0/XI0_6/d__11_ XI11_0/XI0/XI0_6/d_11_ DECAP_INV_G11
XG16566 XI11_0/XI0/XI0_6/d__10_ XI11_0/XI0/XI0_6/d_10_ DECAP_INV_G11
XG16567 XI11_0/XI0/XI0_6/d__9_ XI11_0/XI0/XI0_6/d_9_ DECAP_INV_G11
XG16568 XI11_0/XI0/XI0_6/d__8_ XI11_0/XI0/XI0_6/d_8_ DECAP_INV_G11
XG16569 XI11_0/XI0/XI0_6/d__7_ XI11_0/XI0/XI0_6/d_7_ DECAP_INV_G11
XG16570 XI11_0/XI0/XI0_6/d__6_ XI11_0/XI0/XI0_6/d_6_ DECAP_INV_G11
XG16571 XI11_0/XI0/XI0_6/d__5_ XI11_0/XI0/XI0_6/d_5_ DECAP_INV_G11
XG16572 XI11_0/XI0/XI0_6/d__4_ XI11_0/XI0/XI0_6/d_4_ DECAP_INV_G11
XG16573 XI11_0/XI0/XI0_6/d__3_ XI11_0/XI0/XI0_6/d_3_ DECAP_INV_G11
XG16574 XI11_0/XI0/XI0_6/d__2_ XI11_0/XI0/XI0_6/d_2_ DECAP_INV_G11
XG16575 XI11_0/XI0/XI0_6/d__1_ XI11_0/XI0/XI0_6/d_1_ DECAP_INV_G11
XG16576 XI11_0/XI0/XI0_6/d__0_ XI11_0/XI0/XI0_6/d_0_ DECAP_INV_G11
XG16577 XI11_0/XI0/XI0_6/d_15_ XI11_0/XI0/XI0_6/d__15_ DECAP_INV_G11
XG16578 XI11_0/XI0/XI0_6/d_14_ XI11_0/XI0/XI0_6/d__14_ DECAP_INV_G11
XG16579 XI11_0/XI0/XI0_6/d_13_ XI11_0/XI0/XI0_6/d__13_ DECAP_INV_G11
XG16580 XI11_0/XI0/XI0_6/d_12_ XI11_0/XI0/XI0_6/d__12_ DECAP_INV_G11
XG16581 XI11_0/XI0/XI0_6/d_11_ XI11_0/XI0/XI0_6/d__11_ DECAP_INV_G11
XG16582 XI11_0/XI0/XI0_6/d_10_ XI11_0/XI0/XI0_6/d__10_ DECAP_INV_G11
XG16583 XI11_0/XI0/XI0_6/d_9_ XI11_0/XI0/XI0_6/d__9_ DECAP_INV_G11
XG16584 XI11_0/XI0/XI0_6/d_8_ XI11_0/XI0/XI0_6/d__8_ DECAP_INV_G11
XG16585 XI11_0/XI0/XI0_6/d_7_ XI11_0/XI0/XI0_6/d__7_ DECAP_INV_G11
XG16586 XI11_0/XI0/XI0_6/d_6_ XI11_0/XI0/XI0_6/d__6_ DECAP_INV_G11
XG16587 XI11_0/XI0/XI0_6/d_5_ XI11_0/XI0/XI0_6/d__5_ DECAP_INV_G11
XG16588 XI11_0/XI0/XI0_6/d_4_ XI11_0/XI0/XI0_6/d__4_ DECAP_INV_G11
XG16589 XI11_0/XI0/XI0_6/d_3_ XI11_0/XI0/XI0_6/d__3_ DECAP_INV_G11
XG16590 XI11_0/XI0/XI0_6/d_2_ XI11_0/XI0/XI0_6/d__2_ DECAP_INV_G11
XG16591 XI11_0/XI0/XI0_6/d_1_ XI11_0/XI0/XI0_6/d__1_ DECAP_INV_G11
XG16592 XI11_0/XI0/XI0_6/d_0_ XI11_0/XI0/XI0_6/d__0_ DECAP_INV_G11
XG16593 XI11_0/XI0/XI0_5/d__15_ XI11_0/XI0/XI0_5/d_15_ DECAP_INV_G11
XG16594 XI11_0/XI0/XI0_5/d__14_ XI11_0/XI0/XI0_5/d_14_ DECAP_INV_G11
XG16595 XI11_0/XI0/XI0_5/d__13_ XI11_0/XI0/XI0_5/d_13_ DECAP_INV_G11
XG16596 XI11_0/XI0/XI0_5/d__12_ XI11_0/XI0/XI0_5/d_12_ DECAP_INV_G11
XG16597 XI11_0/XI0/XI0_5/d__11_ XI11_0/XI0/XI0_5/d_11_ DECAP_INV_G11
XG16598 XI11_0/XI0/XI0_5/d__10_ XI11_0/XI0/XI0_5/d_10_ DECAP_INV_G11
XG16599 XI11_0/XI0/XI0_5/d__9_ XI11_0/XI0/XI0_5/d_9_ DECAP_INV_G11
XG16600 XI11_0/XI0/XI0_5/d__8_ XI11_0/XI0/XI0_5/d_8_ DECAP_INV_G11
XG16601 XI11_0/XI0/XI0_5/d__7_ XI11_0/XI0/XI0_5/d_7_ DECAP_INV_G11
XG16602 XI11_0/XI0/XI0_5/d__6_ XI11_0/XI0/XI0_5/d_6_ DECAP_INV_G11
XG16603 XI11_0/XI0/XI0_5/d__5_ XI11_0/XI0/XI0_5/d_5_ DECAP_INV_G11
XG16604 XI11_0/XI0/XI0_5/d__4_ XI11_0/XI0/XI0_5/d_4_ DECAP_INV_G11
XG16605 XI11_0/XI0/XI0_5/d__3_ XI11_0/XI0/XI0_5/d_3_ DECAP_INV_G11
XG16606 XI11_0/XI0/XI0_5/d__2_ XI11_0/XI0/XI0_5/d_2_ DECAP_INV_G11
XG16607 XI11_0/XI0/XI0_5/d__1_ XI11_0/XI0/XI0_5/d_1_ DECAP_INV_G11
XG16608 XI11_0/XI0/XI0_5/d__0_ XI11_0/XI0/XI0_5/d_0_ DECAP_INV_G11
XG16609 XI11_0/XI0/XI0_5/d_15_ XI11_0/XI0/XI0_5/d__15_ DECAP_INV_G11
XG16610 XI11_0/XI0/XI0_5/d_14_ XI11_0/XI0/XI0_5/d__14_ DECAP_INV_G11
XG16611 XI11_0/XI0/XI0_5/d_13_ XI11_0/XI0/XI0_5/d__13_ DECAP_INV_G11
XG16612 XI11_0/XI0/XI0_5/d_12_ XI11_0/XI0/XI0_5/d__12_ DECAP_INV_G11
XG16613 XI11_0/XI0/XI0_5/d_11_ XI11_0/XI0/XI0_5/d__11_ DECAP_INV_G11
XG16614 XI11_0/XI0/XI0_5/d_10_ XI11_0/XI0/XI0_5/d__10_ DECAP_INV_G11
XG16615 XI11_0/XI0/XI0_5/d_9_ XI11_0/XI0/XI0_5/d__9_ DECAP_INV_G11
XG16616 XI11_0/XI0/XI0_5/d_8_ XI11_0/XI0/XI0_5/d__8_ DECAP_INV_G11
XG16617 XI11_0/XI0/XI0_5/d_7_ XI11_0/XI0/XI0_5/d__7_ DECAP_INV_G11
XG16618 XI11_0/XI0/XI0_5/d_6_ XI11_0/XI0/XI0_5/d__6_ DECAP_INV_G11
XG16619 XI11_0/XI0/XI0_5/d_5_ XI11_0/XI0/XI0_5/d__5_ DECAP_INV_G11
XG16620 XI11_0/XI0/XI0_5/d_4_ XI11_0/XI0/XI0_5/d__4_ DECAP_INV_G11
XG16621 XI11_0/XI0/XI0_5/d_3_ XI11_0/XI0/XI0_5/d__3_ DECAP_INV_G11
XG16622 XI11_0/XI0/XI0_5/d_2_ XI11_0/XI0/XI0_5/d__2_ DECAP_INV_G11
XG16623 XI11_0/XI0/XI0_5/d_1_ XI11_0/XI0/XI0_5/d__1_ DECAP_INV_G11
XG16624 XI11_0/XI0/XI0_5/d_0_ XI11_0/XI0/XI0_5/d__0_ DECAP_INV_G11
XG16625 XI11_0/XI0/XI0_4/d__15_ XI11_0/XI0/XI0_4/d_15_ DECAP_INV_G11
XG16626 XI11_0/XI0/XI0_4/d__14_ XI11_0/XI0/XI0_4/d_14_ DECAP_INV_G11
XG16627 XI11_0/XI0/XI0_4/d__13_ XI11_0/XI0/XI0_4/d_13_ DECAP_INV_G11
XG16628 XI11_0/XI0/XI0_4/d__12_ XI11_0/XI0/XI0_4/d_12_ DECAP_INV_G11
XG16629 XI11_0/XI0/XI0_4/d__11_ XI11_0/XI0/XI0_4/d_11_ DECAP_INV_G11
XG16630 XI11_0/XI0/XI0_4/d__10_ XI11_0/XI0/XI0_4/d_10_ DECAP_INV_G11
XG16631 XI11_0/XI0/XI0_4/d__9_ XI11_0/XI0/XI0_4/d_9_ DECAP_INV_G11
XG16632 XI11_0/XI0/XI0_4/d__8_ XI11_0/XI0/XI0_4/d_8_ DECAP_INV_G11
XG16633 XI11_0/XI0/XI0_4/d__7_ XI11_0/XI0/XI0_4/d_7_ DECAP_INV_G11
XG16634 XI11_0/XI0/XI0_4/d__6_ XI11_0/XI0/XI0_4/d_6_ DECAP_INV_G11
XG16635 XI11_0/XI0/XI0_4/d__5_ XI11_0/XI0/XI0_4/d_5_ DECAP_INV_G11
XG16636 XI11_0/XI0/XI0_4/d__4_ XI11_0/XI0/XI0_4/d_4_ DECAP_INV_G11
XG16637 XI11_0/XI0/XI0_4/d__3_ XI11_0/XI0/XI0_4/d_3_ DECAP_INV_G11
XG16638 XI11_0/XI0/XI0_4/d__2_ XI11_0/XI0/XI0_4/d_2_ DECAP_INV_G11
XG16639 XI11_0/XI0/XI0_4/d__1_ XI11_0/XI0/XI0_4/d_1_ DECAP_INV_G11
XG16640 XI11_0/XI0/XI0_4/d__0_ XI11_0/XI0/XI0_4/d_0_ DECAP_INV_G11
XG16641 XI11_0/XI0/XI0_4/d_15_ XI11_0/XI0/XI0_4/d__15_ DECAP_INV_G11
XG16642 XI11_0/XI0/XI0_4/d_14_ XI11_0/XI0/XI0_4/d__14_ DECAP_INV_G11
XG16643 XI11_0/XI0/XI0_4/d_13_ XI11_0/XI0/XI0_4/d__13_ DECAP_INV_G11
XG16644 XI11_0/XI0/XI0_4/d_12_ XI11_0/XI0/XI0_4/d__12_ DECAP_INV_G11
XG16645 XI11_0/XI0/XI0_4/d_11_ XI11_0/XI0/XI0_4/d__11_ DECAP_INV_G11
XG16646 XI11_0/XI0/XI0_4/d_10_ XI11_0/XI0/XI0_4/d__10_ DECAP_INV_G11
XG16647 XI11_0/XI0/XI0_4/d_9_ XI11_0/XI0/XI0_4/d__9_ DECAP_INV_G11
XG16648 XI11_0/XI0/XI0_4/d_8_ XI11_0/XI0/XI0_4/d__8_ DECAP_INV_G11
XG16649 XI11_0/XI0/XI0_4/d_7_ XI11_0/XI0/XI0_4/d__7_ DECAP_INV_G11
XG16650 XI11_0/XI0/XI0_4/d_6_ XI11_0/XI0/XI0_4/d__6_ DECAP_INV_G11
XG16651 XI11_0/XI0/XI0_4/d_5_ XI11_0/XI0/XI0_4/d__5_ DECAP_INV_G11
XG16652 XI11_0/XI0/XI0_4/d_4_ XI11_0/XI0/XI0_4/d__4_ DECAP_INV_G11
XG16653 XI11_0/XI0/XI0_4/d_3_ XI11_0/XI0/XI0_4/d__3_ DECAP_INV_G11
XG16654 XI11_0/XI0/XI0_4/d_2_ XI11_0/XI0/XI0_4/d__2_ DECAP_INV_G11
XG16655 XI11_0/XI0/XI0_4/d_1_ XI11_0/XI0/XI0_4/d__1_ DECAP_INV_G11
XG16656 XI11_0/XI0/XI0_4/d_0_ XI11_0/XI0/XI0_4/d__0_ DECAP_INV_G11
XG16657 XI11_0/XI0/XI0_3/d__15_ XI11_0/XI0/XI0_3/d_15_ DECAP_INV_G11
XG16658 XI11_0/XI0/XI0_3/d__14_ XI11_0/XI0/XI0_3/d_14_ DECAP_INV_G11
XG16659 XI11_0/XI0/XI0_3/d__13_ XI11_0/XI0/XI0_3/d_13_ DECAP_INV_G11
XG16660 XI11_0/XI0/XI0_3/d__12_ XI11_0/XI0/XI0_3/d_12_ DECAP_INV_G11
XG16661 XI11_0/XI0/XI0_3/d__11_ XI11_0/XI0/XI0_3/d_11_ DECAP_INV_G11
XG16662 XI11_0/XI0/XI0_3/d__10_ XI11_0/XI0/XI0_3/d_10_ DECAP_INV_G11
XG16663 XI11_0/XI0/XI0_3/d__9_ XI11_0/XI0/XI0_3/d_9_ DECAP_INV_G11
XG16664 XI11_0/XI0/XI0_3/d__8_ XI11_0/XI0/XI0_3/d_8_ DECAP_INV_G11
XG16665 XI11_0/XI0/XI0_3/d__7_ XI11_0/XI0/XI0_3/d_7_ DECAP_INV_G11
XG16666 XI11_0/XI0/XI0_3/d__6_ XI11_0/XI0/XI0_3/d_6_ DECAP_INV_G11
XG16667 XI11_0/XI0/XI0_3/d__5_ XI11_0/XI0/XI0_3/d_5_ DECAP_INV_G11
XG16668 XI11_0/XI0/XI0_3/d__4_ XI11_0/XI0/XI0_3/d_4_ DECAP_INV_G11
XG16669 XI11_0/XI0/XI0_3/d__3_ XI11_0/XI0/XI0_3/d_3_ DECAP_INV_G11
XG16670 XI11_0/XI0/XI0_3/d__2_ XI11_0/XI0/XI0_3/d_2_ DECAP_INV_G11
XG16671 XI11_0/XI0/XI0_3/d__1_ XI11_0/XI0/XI0_3/d_1_ DECAP_INV_G11
XG16672 XI11_0/XI0/XI0_3/d__0_ XI11_0/XI0/XI0_3/d_0_ DECAP_INV_G11
XG16673 XI11_0/XI0/XI0_3/d_15_ XI11_0/XI0/XI0_3/d__15_ DECAP_INV_G11
XG16674 XI11_0/XI0/XI0_3/d_14_ XI11_0/XI0/XI0_3/d__14_ DECAP_INV_G11
XG16675 XI11_0/XI0/XI0_3/d_13_ XI11_0/XI0/XI0_3/d__13_ DECAP_INV_G11
XG16676 XI11_0/XI0/XI0_3/d_12_ XI11_0/XI0/XI0_3/d__12_ DECAP_INV_G11
XG16677 XI11_0/XI0/XI0_3/d_11_ XI11_0/XI0/XI0_3/d__11_ DECAP_INV_G11
XG16678 XI11_0/XI0/XI0_3/d_10_ XI11_0/XI0/XI0_3/d__10_ DECAP_INV_G11
XG16679 XI11_0/XI0/XI0_3/d_9_ XI11_0/XI0/XI0_3/d__9_ DECAP_INV_G11
XG16680 XI11_0/XI0/XI0_3/d_8_ XI11_0/XI0/XI0_3/d__8_ DECAP_INV_G11
XG16681 XI11_0/XI0/XI0_3/d_7_ XI11_0/XI0/XI0_3/d__7_ DECAP_INV_G11
XG16682 XI11_0/XI0/XI0_3/d_6_ XI11_0/XI0/XI0_3/d__6_ DECAP_INV_G11
XG16683 XI11_0/XI0/XI0_3/d_5_ XI11_0/XI0/XI0_3/d__5_ DECAP_INV_G11
XG16684 XI11_0/XI0/XI0_3/d_4_ XI11_0/XI0/XI0_3/d__4_ DECAP_INV_G11
XG16685 XI11_0/XI0/XI0_3/d_3_ XI11_0/XI0/XI0_3/d__3_ DECAP_INV_G11
XG16686 XI11_0/XI0/XI0_3/d_2_ XI11_0/XI0/XI0_3/d__2_ DECAP_INV_G11
XG16687 XI11_0/XI0/XI0_3/d_1_ XI11_0/XI0/XI0_3/d__1_ DECAP_INV_G11
XG16688 XI11_0/XI0/XI0_3/d_0_ XI11_0/XI0/XI0_3/d__0_ DECAP_INV_G11
XG16689 XI11_0/XI0/XI0_2/d__15_ XI11_0/XI0/XI0_2/d_15_ DECAP_INV_G11
XG16690 XI11_0/XI0/XI0_2/d__14_ XI11_0/XI0/XI0_2/d_14_ DECAP_INV_G11
XG16691 XI11_0/XI0/XI0_2/d__13_ XI11_0/XI0/XI0_2/d_13_ DECAP_INV_G11
XG16692 XI11_0/XI0/XI0_2/d__12_ XI11_0/XI0/XI0_2/d_12_ DECAP_INV_G11
XG16693 XI11_0/XI0/XI0_2/d__11_ XI11_0/XI0/XI0_2/d_11_ DECAP_INV_G11
XG16694 XI11_0/XI0/XI0_2/d__10_ XI11_0/XI0/XI0_2/d_10_ DECAP_INV_G11
XG16695 XI11_0/XI0/XI0_2/d__9_ XI11_0/XI0/XI0_2/d_9_ DECAP_INV_G11
XG16696 XI11_0/XI0/XI0_2/d__8_ XI11_0/XI0/XI0_2/d_8_ DECAP_INV_G11
XG16697 XI11_0/XI0/XI0_2/d__7_ XI11_0/XI0/XI0_2/d_7_ DECAP_INV_G11
XG16698 XI11_0/XI0/XI0_2/d__6_ XI11_0/XI0/XI0_2/d_6_ DECAP_INV_G11
XG16699 XI11_0/XI0/XI0_2/d__5_ XI11_0/XI0/XI0_2/d_5_ DECAP_INV_G11
XG16700 XI11_0/XI0/XI0_2/d__4_ XI11_0/XI0/XI0_2/d_4_ DECAP_INV_G11
XG16701 XI11_0/XI0/XI0_2/d__3_ XI11_0/XI0/XI0_2/d_3_ DECAP_INV_G11
XG16702 XI11_0/XI0/XI0_2/d__2_ XI11_0/XI0/XI0_2/d_2_ DECAP_INV_G11
XG16703 XI11_0/XI0/XI0_2/d__1_ XI11_0/XI0/XI0_2/d_1_ DECAP_INV_G11
XG16704 XI11_0/XI0/XI0_2/d__0_ XI11_0/XI0/XI0_2/d_0_ DECAP_INV_G11
XG16705 XI11_0/XI0/XI0_2/d_15_ XI11_0/XI0/XI0_2/d__15_ DECAP_INV_G11
XG16706 XI11_0/XI0/XI0_2/d_14_ XI11_0/XI0/XI0_2/d__14_ DECAP_INV_G11
XG16707 XI11_0/XI0/XI0_2/d_13_ XI11_0/XI0/XI0_2/d__13_ DECAP_INV_G11
XG16708 XI11_0/XI0/XI0_2/d_12_ XI11_0/XI0/XI0_2/d__12_ DECAP_INV_G11
XG16709 XI11_0/XI0/XI0_2/d_11_ XI11_0/XI0/XI0_2/d__11_ DECAP_INV_G11
XG16710 XI11_0/XI0/XI0_2/d_10_ XI11_0/XI0/XI0_2/d__10_ DECAP_INV_G11
XG16711 XI11_0/XI0/XI0_2/d_9_ XI11_0/XI0/XI0_2/d__9_ DECAP_INV_G11
XG16712 XI11_0/XI0/XI0_2/d_8_ XI11_0/XI0/XI0_2/d__8_ DECAP_INV_G11
XG16713 XI11_0/XI0/XI0_2/d_7_ XI11_0/XI0/XI0_2/d__7_ DECAP_INV_G11
XG16714 XI11_0/XI0/XI0_2/d_6_ XI11_0/XI0/XI0_2/d__6_ DECAP_INV_G11
XG16715 XI11_0/XI0/XI0_2/d_5_ XI11_0/XI0/XI0_2/d__5_ DECAP_INV_G11
XG16716 XI11_0/XI0/XI0_2/d_4_ XI11_0/XI0/XI0_2/d__4_ DECAP_INV_G11
XG16717 XI11_0/XI0/XI0_2/d_3_ XI11_0/XI0/XI0_2/d__3_ DECAP_INV_G11
XG16718 XI11_0/XI0/XI0_2/d_2_ XI11_0/XI0/XI0_2/d__2_ DECAP_INV_G11
XG16719 XI11_0/XI0/XI0_2/d_1_ XI11_0/XI0/XI0_2/d__1_ DECAP_INV_G11
XG16720 XI11_0/XI0/XI0_2/d_0_ XI11_0/XI0/XI0_2/d__0_ DECAP_INV_G11
XG16721 XI11_0/XI0/XI0_1/d__15_ XI11_0/XI0/XI0_1/d_15_ DECAP_INV_G11
XG16722 XI11_0/XI0/XI0_1/d__14_ XI11_0/XI0/XI0_1/d_14_ DECAP_INV_G11
XG16723 XI11_0/XI0/XI0_1/d__13_ XI11_0/XI0/XI0_1/d_13_ DECAP_INV_G11
XG16724 XI11_0/XI0/XI0_1/d__12_ XI11_0/XI0/XI0_1/d_12_ DECAP_INV_G11
XG16725 XI11_0/XI0/XI0_1/d__11_ XI11_0/XI0/XI0_1/d_11_ DECAP_INV_G11
XG16726 XI11_0/XI0/XI0_1/d__10_ XI11_0/XI0/XI0_1/d_10_ DECAP_INV_G11
XG16727 XI11_0/XI0/XI0_1/d__9_ XI11_0/XI0/XI0_1/d_9_ DECAP_INV_G11
XG16728 XI11_0/XI0/XI0_1/d__8_ XI11_0/XI0/XI0_1/d_8_ DECAP_INV_G11
XG16729 XI11_0/XI0/XI0_1/d__7_ XI11_0/XI0/XI0_1/d_7_ DECAP_INV_G11
XG16730 XI11_0/XI0/XI0_1/d__6_ XI11_0/XI0/XI0_1/d_6_ DECAP_INV_G11
XG16731 XI11_0/XI0/XI0_1/d__5_ XI11_0/XI0/XI0_1/d_5_ DECAP_INV_G11
XG16732 XI11_0/XI0/XI0_1/d__4_ XI11_0/XI0/XI0_1/d_4_ DECAP_INV_G11
XG16733 XI11_0/XI0/XI0_1/d__3_ XI11_0/XI0/XI0_1/d_3_ DECAP_INV_G11
XG16734 XI11_0/XI0/XI0_1/d__2_ XI11_0/XI0/XI0_1/d_2_ DECAP_INV_G11
XG16735 XI11_0/XI0/XI0_1/d__1_ XI11_0/XI0/XI0_1/d_1_ DECAP_INV_G11
XG16736 XI11_0/XI0/XI0_1/d__0_ XI11_0/XI0/XI0_1/d_0_ DECAP_INV_G11
XG16737 XI11_0/XI0/XI0_1/d_15_ XI11_0/XI0/XI0_1/d__15_ DECAP_INV_G11
XG16738 XI11_0/XI0/XI0_1/d_14_ XI11_0/XI0/XI0_1/d__14_ DECAP_INV_G11
XG16739 XI11_0/XI0/XI0_1/d_13_ XI11_0/XI0/XI0_1/d__13_ DECAP_INV_G11
XG16740 XI11_0/XI0/XI0_1/d_12_ XI11_0/XI0/XI0_1/d__12_ DECAP_INV_G11
XG16741 XI11_0/XI0/XI0_1/d_11_ XI11_0/XI0/XI0_1/d__11_ DECAP_INV_G11
XG16742 XI11_0/XI0/XI0_1/d_10_ XI11_0/XI0/XI0_1/d__10_ DECAP_INV_G11
XG16743 XI11_0/XI0/XI0_1/d_9_ XI11_0/XI0/XI0_1/d__9_ DECAP_INV_G11
XG16744 XI11_0/XI0/XI0_1/d_8_ XI11_0/XI0/XI0_1/d__8_ DECAP_INV_G11
XG16745 XI11_0/XI0/XI0_1/d_7_ XI11_0/XI0/XI0_1/d__7_ DECAP_INV_G11
XG16746 XI11_0/XI0/XI0_1/d_6_ XI11_0/XI0/XI0_1/d__6_ DECAP_INV_G11
XG16747 XI11_0/XI0/XI0_1/d_5_ XI11_0/XI0/XI0_1/d__5_ DECAP_INV_G11
XG16748 XI11_0/XI0/XI0_1/d_4_ XI11_0/XI0/XI0_1/d__4_ DECAP_INV_G11
XG16749 XI11_0/XI0/XI0_1/d_3_ XI11_0/XI0/XI0_1/d__3_ DECAP_INV_G11
XG16750 XI11_0/XI0/XI0_1/d_2_ XI11_0/XI0/XI0_1/d__2_ DECAP_INV_G11
XG16751 XI11_0/XI0/XI0_1/d_1_ XI11_0/XI0/XI0_1/d__1_ DECAP_INV_G11
XG16752 XI11_0/XI0/XI0_1/d_0_ XI11_0/XI0/XI0_1/d__0_ DECAP_INV_G11
XG16753 XI11_0/XI0/XI0_0/d__15_ XI11_0/XI0/XI0_0/d_15_ DECAP_INV_G11
XG16754 XI11_0/XI0/XI0_0/d__14_ XI11_0/XI0/XI0_0/d_14_ DECAP_INV_G11
XG16755 XI11_0/XI0/XI0_0/d__13_ XI11_0/XI0/XI0_0/d_13_ DECAP_INV_G11
XG16756 XI11_0/XI0/XI0_0/d__12_ XI11_0/XI0/XI0_0/d_12_ DECAP_INV_G11
XG16757 XI11_0/XI0/XI0_0/d__11_ XI11_0/XI0/XI0_0/d_11_ DECAP_INV_G11
XG16758 XI11_0/XI0/XI0_0/d__10_ XI11_0/XI0/XI0_0/d_10_ DECAP_INV_G11
XG16759 XI11_0/XI0/XI0_0/d__9_ XI11_0/XI0/XI0_0/d_9_ DECAP_INV_G11
XG16760 XI11_0/XI0/XI0_0/d__8_ XI11_0/XI0/XI0_0/d_8_ DECAP_INV_G11
XG16761 XI11_0/XI0/XI0_0/d__7_ XI11_0/XI0/XI0_0/d_7_ DECAP_INV_G11
XG16762 XI11_0/XI0/XI0_0/d__6_ XI11_0/XI0/XI0_0/d_6_ DECAP_INV_G11
XG16763 XI11_0/XI0/XI0_0/d__5_ XI11_0/XI0/XI0_0/d_5_ DECAP_INV_G11
XG16764 XI11_0/XI0/XI0_0/d__4_ XI11_0/XI0/XI0_0/d_4_ DECAP_INV_G11
XG16765 XI11_0/XI0/XI0_0/d__3_ XI11_0/XI0/XI0_0/d_3_ DECAP_INV_G11
XG16766 XI11_0/XI0/XI0_0/d__2_ XI11_0/XI0/XI0_0/d_2_ DECAP_INV_G11
XG16767 XI11_0/XI0/XI0_0/d__1_ XI11_0/XI0/XI0_0/d_1_ DECAP_INV_G11
XG16768 XI11_0/XI0/XI0_0/d__0_ XI11_0/XI0/XI0_0/d_0_ DECAP_INV_G11
XG16769 XI11_0/XI0/XI0_0/d_15_ XI11_0/XI0/XI0_0/d__15_ DECAP_INV_G11
XG16770 XI11_0/XI0/XI0_0/d_14_ XI11_0/XI0/XI0_0/d__14_ DECAP_INV_G11
XG16771 XI11_0/XI0/XI0_0/d_13_ XI11_0/XI0/XI0_0/d__13_ DECAP_INV_G11
XG16772 XI11_0/XI0/XI0_0/d_12_ XI11_0/XI0/XI0_0/d__12_ DECAP_INV_G11
XG16773 XI11_0/XI0/XI0_0/d_11_ XI11_0/XI0/XI0_0/d__11_ DECAP_INV_G11
XG16774 XI11_0/XI0/XI0_0/d_10_ XI11_0/XI0/XI0_0/d__10_ DECAP_INV_G11
XG16775 XI11_0/XI0/XI0_0/d_9_ XI11_0/XI0/XI0_0/d__9_ DECAP_INV_G11
XG16776 XI11_0/XI0/XI0_0/d_8_ XI11_0/XI0/XI0_0/d__8_ DECAP_INV_G11
XG16777 XI11_0/XI0/XI0_0/d_7_ XI11_0/XI0/XI0_0/d__7_ DECAP_INV_G11
XG16778 XI11_0/XI0/XI0_0/d_6_ XI11_0/XI0/XI0_0/d__6_ DECAP_INV_G11
XG16779 XI11_0/XI0/XI0_0/d_5_ XI11_0/XI0/XI0_0/d__5_ DECAP_INV_G11
XG16780 XI11_0/XI0/XI0_0/d_4_ XI11_0/XI0/XI0_0/d__4_ DECAP_INV_G11
XG16781 XI11_0/XI0/XI0_0/d_3_ XI11_0/XI0/XI0_0/d__3_ DECAP_INV_G11
XG16782 XI11_0/XI0/XI0_0/d_2_ XI11_0/XI0/XI0_0/d__2_ DECAP_INV_G11
XG16783 XI11_0/XI0/XI0_0/d_1_ XI11_0/XI0/XI0_0/d__1_ DECAP_INV_G11
XG16784 XI11_0/XI0/XI0_0/d_0_ XI11_0/XI0/XI0_0/d__0_ DECAP_INV_G11
XG16785 XI10/XI0/net095 XI10/net022 DECAP_INV_G12
XG16786 XI10/XI0/net090 XI10/sck DECAP_INV_G12
XG16787 CS XI10/XI0/net044 DECAP_INV_G10
XG16788 XI10/net036 sck_bar DECAP_INV_G13
XG16789 XI10/net030 sck_bar DECAP_INV_G13
XG16790 XI10/net038 XI10/net030 DECAP_INV_G14
XG16791 XI10/net038 XI10/net036 DECAP_INV_G14
XG16792 XI10/sck XI10/net038 DECAP_INV_G14
XG16793 XI5/net028_0_ XI5/net023_0_ DECAP_INV_G15
XG16794 XI5/net028_1_ XI5/net023_1_ DECAP_INV_G15
XG16795 XI5/net028_2_ XI5/net023_2_ DECAP_INV_G15
XG16796 XI5/net028_3_ XI5/net023_3_ DECAP_INV_G15
XG16797 XI5/net028_4_ XI5/net023_4_ DECAP_INV_G15
XG16798 XI5/net028_5_ XI5/net023_5_ DECAP_INV_G15
XG16799 XI5/net028_6_ XI5/net023_6_ DECAP_INV_G15
XG16800 XI5/net028_7_ XI5/net023_7_ DECAP_INV_G15
XG16801 XI5/net023_0_ wrdata_7_ DECAP_INV_G12
XG16802 XI5/net023_1_ wrdata_6_ DECAP_INV_G12
XG16803 XI5/net023_2_ wrdata_5_ DECAP_INV_G12
XG16804 XI5/net023_3_ wrdata_4_ DECAP_INV_G12
XG16805 XI5/net023_4_ wrdata_3_ DECAP_INV_G12
XG16806 XI5/net023_5_ wrdata_2_ DECAP_INV_G12
XG16807 XI5/net023_6_ wrdata_1_ DECAP_INV_G12
XG16808 XI5/net023_7_ wrdata_0_ DECAP_INV_G12
XG16809 XI5/net025_0_ XI5/net017_0_ DECAP_INV_G15
XG16810 XI5/net025_1_ XI5/net017_1_ DECAP_INV_G15
XG16811 XI5/net025_2_ XI5/net017_2_ DECAP_INV_G15
XG16812 XI5/net025_3_ XI5/net017_3_ DECAP_INV_G15
XG16813 XI5/net025_4_ XI5/net017_4_ DECAP_INV_G15
XG16814 XI5/net025_5_ XI5/net017_5_ DECAP_INV_G15
XG16815 XI5/net025_6_ XI5/net017_6_ DECAP_INV_G15
XG16816 XI5/net025_7_ XI5/net017_7_ DECAP_INV_G15
XG16817 XI5/net017_0_ wrdata__7_ DECAP_INV_G12
XG16818 XI5/net017_1_ wrdata__6_ DECAP_INV_G12
XG16819 XI5/net017_2_ wrdata__5_ DECAP_INV_G12
XG16820 XI5/net017_3_ wrdata__4_ DECAP_INV_G12
XG16821 XI5/net017_4_ wrdata__3_ DECAP_INV_G12
XG16822 XI5/net017_5_ wrdata__2_ DECAP_INV_G12
XG16823 XI5/net017_6_ wrdata__1_ DECAP_INV_G12
XG16824 XI5/net017_7_ wrdata__0_ DECAP_INV_G12
XG16825 XI5/XI4_7/net24 XI5/net028_0_ DECAP_INV_G16
XG16826 XI5/XI4_7/s XI5/net025_0_ DECAP_INV_G16
XG16827 XI5/XI4_7/net24 XI5/XI4_7/s DECAP_INV_G17
XG16828 XI5/XI4_7/pm XI5/XI4_7/m DECAP_INV_G18
XG16829 XI5/XI4_7/cn XI5/XI4_7/c DECAP_INV_G19
XG16830 XI5/ck XI5/XI4_7/cn DECAP_INV_G20
XG16831 XI5/XI4_6/net24 XI5/net028_1_ DECAP_INV_G16
XG16832 XI5/XI4_6/s XI5/net025_1_ DECAP_INV_G16
XG16833 XI5/XI4_6/net24 XI5/XI4_6/s DECAP_INV_G17
XG16834 XI5/XI4_6/pm XI5/XI4_6/m DECAP_INV_G18
XG16835 XI5/XI4_6/cn XI5/XI4_6/c DECAP_INV_G19
XG16836 XI5/ck XI5/XI4_6/cn DECAP_INV_G20
XG16837 XI5/XI4_5/net24 XI5/net028_2_ DECAP_INV_G16
XG16838 XI5/XI4_5/s XI5/net025_2_ DECAP_INV_G16
XG16839 XI5/XI4_5/net24 XI5/XI4_5/s DECAP_INV_G17
XG16840 XI5/XI4_5/pm XI5/XI4_5/m DECAP_INV_G18
XG16841 XI5/XI4_5/cn XI5/XI4_5/c DECAP_INV_G19
XG16842 XI5/ck XI5/XI4_5/cn DECAP_INV_G20
XG16843 XI5/XI4_4/net24 XI5/net028_3_ DECAP_INV_G16
XG16844 XI5/XI4_4/s XI5/net025_3_ DECAP_INV_G16
XG16845 XI5/XI4_4/net24 XI5/XI4_4/s DECAP_INV_G17
XG16846 XI5/XI4_4/pm XI5/XI4_4/m DECAP_INV_G18
XG16847 XI5/XI4_4/cn XI5/XI4_4/c DECAP_INV_G19
XG16848 XI5/ck XI5/XI4_4/cn DECAP_INV_G20
XG16849 XI5/XI4_3/net24 XI5/net028_4_ DECAP_INV_G16
XG16850 XI5/XI4_3/s XI5/net025_4_ DECAP_INV_G16
XG16851 XI5/XI4_3/net24 XI5/XI4_3/s DECAP_INV_G17
XG16852 XI5/XI4_3/pm XI5/XI4_3/m DECAP_INV_G18
XG16853 XI5/XI4_3/cn XI5/XI4_3/c DECAP_INV_G19
XG16854 XI5/ck XI5/XI4_3/cn DECAP_INV_G20
XG16855 XI5/XI4_2/net24 XI5/net028_5_ DECAP_INV_G16
XG16856 XI5/XI4_2/s XI5/net025_5_ DECAP_INV_G16
XG16857 XI5/XI4_2/net24 XI5/XI4_2/s DECAP_INV_G17
XG16858 XI5/XI4_2/pm XI5/XI4_2/m DECAP_INV_G18
XG16859 XI5/XI4_2/cn XI5/XI4_2/c DECAP_INV_G19
XG16860 XI5/ck XI5/XI4_2/cn DECAP_INV_G20
XG16861 XI5/XI4_1/net24 XI5/net028_6_ DECAP_INV_G16
XG16862 XI5/XI4_1/s XI5/net025_6_ DECAP_INV_G16
XG16863 XI5/XI4_1/net24 XI5/XI4_1/s DECAP_INV_G17
XG16864 XI5/XI4_1/pm XI5/XI4_1/m DECAP_INV_G18
XG16865 XI5/XI4_1/cn XI5/XI4_1/c DECAP_INV_G19
XG16866 XI5/ck XI5/XI4_1/cn DECAP_INV_G20
XG16867 XI5/XI4_0/net24 XI5/net028_7_ DECAP_INV_G16
XG16868 XI5/XI4_0/s XI5/net025_7_ DECAP_INV_G16
XG16869 XI5/XI4_0/net24 XI5/XI4_0/s DECAP_INV_G17
XG16870 XI5/XI4_0/pm XI5/XI4_0/m DECAP_INV_G18
XG16871 XI5/XI4_0/cn XI5/XI4_0/c DECAP_INV_G19
XG16872 XI5/ck XI5/XI4_0/cn DECAP_INV_G20
XG16873 XI5/XI6/net25 XI5/XI6/net16 DECAP_INV_G21
XG16874 XI5/XI6/net16 XI5/ck DECAP_INV_G22
XG16875 sck_bar XI5/XI6/net25 DECAP_INV_G23
XG16876 XI5/XI2/net095 XI5/net23 DECAP_INV_G12
XG16877 XI5/XI2/net090 rd_en DECAP_INV_G12
XG16878 RD XI5/XI2/net044 DECAP_INV_G10
XG16879 XI5/XI1/net095 XI5/net27 DECAP_INV_G12
XG16880 XI5/XI1/net090 wr_en DECAP_INV_G12
XG16881 WR XI5/XI1/net044 DECAP_INV_G10
XG16882 XI5/XI0_9/net095 addr__9_ DECAP_INV_G12
XG16883 XI5/XI0_9/net090 addr_9_ DECAP_INV_G12
XG16884 A_9_ XI5/XI0_9/net044 DECAP_INV_G10
XG16885 XI5/XI0_8/net095 addr__8_ DECAP_INV_G12
XG16886 XI5/XI0_8/net090 addr_8_ DECAP_INV_G12
XG16887 A_8_ XI5/XI0_8/net044 DECAP_INV_G10
XG16888 XI5/XI0_7/net095 addr__7_ DECAP_INV_G12
XG16889 XI5/XI0_7/net090 addr_7_ DECAP_INV_G12
XG16890 A_7_ XI5/XI0_7/net044 DECAP_INV_G10
XG16891 XI5/XI0_6/net095 addr__6_ DECAP_INV_G12
XG16892 XI5/XI0_6/net090 addr_6_ DECAP_INV_G12
XG16893 A_6_ XI5/XI0_6/net044 DECAP_INV_G10
XG16894 XI5/XI0_5/net095 addr__5_ DECAP_INV_G12
XG16895 XI5/XI0_5/net090 addr_5_ DECAP_INV_G12
XG16896 A_5_ XI5/XI0_5/net044 DECAP_INV_G10
XG16897 XI5/XI0_4/net095 addr__4_ DECAP_INV_G12
XG16898 XI5/XI0_4/net090 addr_4_ DECAP_INV_G12
XG16899 A_4_ XI5/XI0_4/net044 DECAP_INV_G10
XG16900 XI5/XI0_3/net095 addr__3_ DECAP_INV_G12
XG16901 XI5/XI0_3/net090 addr_3_ DECAP_INV_G12
XG16902 A_3_ XI5/XI0_3/net044 DECAP_INV_G10
XG16903 XI5/XI0_2/net095 addr__2_ DECAP_INV_G12
XG16904 XI5/XI0_2/net090 addr_2_ DECAP_INV_G12
XG16905 A_2_ XI5/XI0_2/net044 DECAP_INV_G10
XG16906 XI5/XI0_1/net095 addr__1_ DECAP_INV_G12
XG16907 XI5/XI0_1/net090 addr_1_ DECAP_INV_G12
XG16908 A_1_ XI5/XI0_1/net044 DECAP_INV_G10
XG16909 XI5/XI0_0/net095 addr__0_ DECAP_INV_G12
XG16910 XI5/XI0_0/net090 addr_0_ DECAP_INV_G12
XG16911 A_0_ XI5/XI0_0/net044 DECAP_INV_G10
XG16912 XI2/net020_0_ xsel_63_ DECAP_INV_G24
XG16913 XI2/net020_1_ xsel_62_ DECAP_INV_G24
XG16914 XI2/net020_2_ xsel_61_ DECAP_INV_G24
XG16915 XI2/net020_3_ xsel_60_ DECAP_INV_G24
XG16916 XI2/net020_4_ xsel_59_ DECAP_INV_G24
XG16917 XI2/net020_5_ xsel_58_ DECAP_INV_G24
XG16918 XI2/net020_6_ xsel_57_ DECAP_INV_G24
XG16919 XI2/net020_7_ xsel_56_ DECAP_INV_G24
XG16920 XI2/net020_8_ xsel_55_ DECAP_INV_G24
XG16921 XI2/net020_9_ xsel_54_ DECAP_INV_G24
XG16922 XI2/net020_10_ xsel_53_ DECAP_INV_G24
XG16923 XI2/net020_11_ xsel_52_ DECAP_INV_G24
XG16924 XI2/net020_12_ xsel_51_ DECAP_INV_G24
XG16925 XI2/net020_13_ xsel_50_ DECAP_INV_G24
XG16926 XI2/net020_14_ xsel_49_ DECAP_INV_G24
XG16927 XI2/net020_15_ xsel_48_ DECAP_INV_G24
XG16928 XI2/net020_16_ xsel_47_ DECAP_INV_G24
XG16929 XI2/net020_17_ xsel_46_ DECAP_INV_G24
XG16930 XI2/net020_18_ xsel_45_ DECAP_INV_G24
XG16931 XI2/net020_19_ xsel_44_ DECAP_INV_G24
XG16932 XI2/net020_20_ xsel_43_ DECAP_INV_G24
XG16933 XI2/net020_21_ xsel_42_ DECAP_INV_G24
XG16934 XI2/net020_22_ xsel_41_ DECAP_INV_G24
XG16935 XI2/net020_23_ xsel_40_ DECAP_INV_G24
XG16936 XI2/net020_24_ xsel_39_ DECAP_INV_G24
XG16937 XI2/net020_25_ xsel_38_ DECAP_INV_G24
XG16938 XI2/net020_26_ xsel_37_ DECAP_INV_G24
XG16939 XI2/net020_27_ xsel_36_ DECAP_INV_G24
XG16940 XI2/net020_28_ xsel_35_ DECAP_INV_G24
XG16941 XI2/net020_29_ xsel_34_ DECAP_INV_G24
XG16942 XI2/net020_30_ xsel_33_ DECAP_INV_G24
XG16943 XI2/net020_31_ xsel_32_ DECAP_INV_G24
XG16944 XI2/net020_32_ xsel_31_ DECAP_INV_G24
XG16945 XI2/net020_33_ xsel_30_ DECAP_INV_G24
XG16946 XI2/net020_34_ xsel_29_ DECAP_INV_G24
XG16947 XI2/net020_35_ xsel_28_ DECAP_INV_G24
XG16948 XI2/net020_36_ xsel_27_ DECAP_INV_G24
XG16949 XI2/net020_37_ xsel_26_ DECAP_INV_G24
XG16950 XI2/net020_38_ xsel_25_ DECAP_INV_G24
XG16951 XI2/net020_39_ xsel_24_ DECAP_INV_G24
XG16952 XI2/net020_40_ xsel_23_ DECAP_INV_G24
XG16953 XI2/net020_41_ xsel_22_ DECAP_INV_G24
XG16954 XI2/net020_42_ xsel_21_ DECAP_INV_G24
XG16955 XI2/net020_43_ xsel_20_ DECAP_INV_G24
XG16956 XI2/net020_44_ xsel_19_ DECAP_INV_G24
XG16957 XI2/net020_45_ xsel_18_ DECAP_INV_G24
XG16958 XI2/net020_46_ xsel_17_ DECAP_INV_G24
XG16959 XI2/net020_47_ xsel_16_ DECAP_INV_G24
XG16960 XI2/net020_48_ xsel_15_ DECAP_INV_G24
XG16961 XI2/net020_49_ xsel_14_ DECAP_INV_G24
XG16962 XI2/net020_50_ xsel_13_ DECAP_INV_G24
XG16963 XI2/net020_51_ xsel_12_ DECAP_INV_G24
XG16964 XI2/net020_52_ xsel_11_ DECAP_INV_G24
XG16965 XI2/net020_53_ xsel_10_ DECAP_INV_G24
XG16966 XI2/net020_54_ xsel_9_ DECAP_INV_G24
XG16967 XI2/net020_55_ xsel_8_ DECAP_INV_G24
XG16968 XI2/net020_56_ xsel_7_ DECAP_INV_G24
XG16969 XI2/net020_57_ xsel_6_ DECAP_INV_G24
XG16970 XI2/net020_58_ xsel_5_ DECAP_INV_G24
XG16971 XI2/net020_59_ xsel_4_ DECAP_INV_G24
XG16972 XI2/net020_60_ xsel_3_ DECAP_INV_G24
XG16973 XI2/net020_61_ xsel_2_ DECAP_INV_G24
XG16974 XI2/net020_62_ xsel_1_ DECAP_INV_G24
XG16975 XI2/net020_63_ xsel_0_ DECAP_INV_G24
XG16976 XI2/net024_0_ XI2/net020_0_ DECAP_INV_G12
XG16977 XI2/net024_1_ XI2/net020_1_ DECAP_INV_G12
XG16978 XI2/net024_2_ XI2/net020_2_ DECAP_INV_G12
XG16979 XI2/net024_3_ XI2/net020_3_ DECAP_INV_G12
XG16980 XI2/net024_4_ XI2/net020_4_ DECAP_INV_G12
XG16981 XI2/net024_5_ XI2/net020_5_ DECAP_INV_G12
XG16982 XI2/net024_6_ XI2/net020_6_ DECAP_INV_G12
XG16983 XI2/net024_7_ XI2/net020_7_ DECAP_INV_G12
XG16984 XI2/net024_8_ XI2/net020_8_ DECAP_INV_G12
XG16985 XI2/net024_9_ XI2/net020_9_ DECAP_INV_G12
XG16986 XI2/net024_10_ XI2/net020_10_ DECAP_INV_G12
XG16987 XI2/net024_11_ XI2/net020_11_ DECAP_INV_G12
XG16988 XI2/net024_12_ XI2/net020_12_ DECAP_INV_G12
XG16989 XI2/net024_13_ XI2/net020_13_ DECAP_INV_G12
XG16990 XI2/net024_14_ XI2/net020_14_ DECAP_INV_G12
XG16991 XI2/net024_15_ XI2/net020_15_ DECAP_INV_G12
XG16992 XI2/net024_16_ XI2/net020_16_ DECAP_INV_G12
XG16993 XI2/net024_17_ XI2/net020_17_ DECAP_INV_G12
XG16994 XI2/net024_18_ XI2/net020_18_ DECAP_INV_G12
XG16995 XI2/net024_19_ XI2/net020_19_ DECAP_INV_G12
XG16996 XI2/net024_20_ XI2/net020_20_ DECAP_INV_G12
XG16997 XI2/net024_21_ XI2/net020_21_ DECAP_INV_G12
XG16998 XI2/net024_22_ XI2/net020_22_ DECAP_INV_G12
XG16999 XI2/net024_23_ XI2/net020_23_ DECAP_INV_G12
XG17000 XI2/net024_24_ XI2/net020_24_ DECAP_INV_G12
XG17001 XI2/net024_25_ XI2/net020_25_ DECAP_INV_G12
XG17002 XI2/net024_26_ XI2/net020_26_ DECAP_INV_G12
XG17003 XI2/net024_27_ XI2/net020_27_ DECAP_INV_G12
XG17004 XI2/net024_28_ XI2/net020_28_ DECAP_INV_G12
XG17005 XI2/net024_29_ XI2/net020_29_ DECAP_INV_G12
XG17006 XI2/net024_30_ XI2/net020_30_ DECAP_INV_G12
XG17007 XI2/net024_31_ XI2/net020_31_ DECAP_INV_G12
XG17008 XI2/net024_32_ XI2/net020_32_ DECAP_INV_G12
XG17009 XI2/net024_33_ XI2/net020_33_ DECAP_INV_G12
XG17010 XI2/net024_34_ XI2/net020_34_ DECAP_INV_G12
XG17011 XI2/net024_35_ XI2/net020_35_ DECAP_INV_G12
XG17012 XI2/net024_36_ XI2/net020_36_ DECAP_INV_G12
XG17013 XI2/net024_37_ XI2/net020_37_ DECAP_INV_G12
XG17014 XI2/net024_38_ XI2/net020_38_ DECAP_INV_G12
XG17015 XI2/net024_39_ XI2/net020_39_ DECAP_INV_G12
XG17016 XI2/net024_40_ XI2/net020_40_ DECAP_INV_G12
XG17017 XI2/net024_41_ XI2/net020_41_ DECAP_INV_G12
XG17018 XI2/net024_42_ XI2/net020_42_ DECAP_INV_G12
XG17019 XI2/net024_43_ XI2/net020_43_ DECAP_INV_G12
XG17020 XI2/net024_44_ XI2/net020_44_ DECAP_INV_G12
XG17021 XI2/net024_45_ XI2/net020_45_ DECAP_INV_G12
XG17022 XI2/net024_46_ XI2/net020_46_ DECAP_INV_G12
XG17023 XI2/net024_47_ XI2/net020_47_ DECAP_INV_G12
XG17024 XI2/net024_48_ XI2/net020_48_ DECAP_INV_G12
XG17025 XI2/net024_49_ XI2/net020_49_ DECAP_INV_G12
XG17026 XI2/net024_50_ XI2/net020_50_ DECAP_INV_G12
XG17027 XI2/net024_51_ XI2/net020_51_ DECAP_INV_G12
XG17028 XI2/net024_52_ XI2/net020_52_ DECAP_INV_G12
XG17029 XI2/net024_53_ XI2/net020_53_ DECAP_INV_G12
XG17030 XI2/net024_54_ XI2/net020_54_ DECAP_INV_G12
XG17031 XI2/net024_55_ XI2/net020_55_ DECAP_INV_G12
XG17032 XI2/net024_56_ XI2/net020_56_ DECAP_INV_G12
XG17033 XI2/net024_57_ XI2/net020_57_ DECAP_INV_G12
XG17034 XI2/net024_58_ XI2/net020_58_ DECAP_INV_G12
XG17035 XI2/net024_59_ XI2/net020_59_ DECAP_INV_G12
XG17036 XI2/net024_60_ XI2/net020_60_ DECAP_INV_G12
XG17037 XI2/net024_61_ XI2/net020_61_ DECAP_INV_G12
XG17038 XI2/net024_62_ XI2/net020_62_ DECAP_INV_G12
XG17039 XI2/net024_63_ XI2/net020_63_ DECAP_INV_G12
XG17040 XI6/net014_0_ XI6/net021_0_ DECAP_INV_G12
XG17041 XI6/net014_1_ XI6/net021_1_ DECAP_INV_G12
XG17042 XI6/net014_2_ XI6/net021_2_ DECAP_INV_G12
XG17043 XI6/net014_3_ XI6/net021_3_ DECAP_INV_G12
XG17044 XI6/net014_4_ XI6/net021_4_ DECAP_INV_G12
XG17045 XI6/net014_5_ XI6/net021_5_ DECAP_INV_G12
XG17046 XI6/net014_6_ XI6/net021_6_ DECAP_INV_G12
XG17047 XI6/net014_7_ XI6/net021_7_ DECAP_INV_G12
XG17048 XI6/net014_8_ XI6/net021_8_ DECAP_INV_G12
XG17049 XI6/net014_9_ XI6/net021_9_ DECAP_INV_G12
XG17050 XI6/net014_10_ XI6/net021_10_ DECAP_INV_G12
XG17051 XI6/net014_11_ XI6/net021_11_ DECAP_INV_G12
XG17052 XI6/net014_12_ XI6/net021_12_ DECAP_INV_G12
XG17053 XI6/net014_13_ XI6/net021_13_ DECAP_INV_G12
XG17054 XI6/net014_14_ XI6/net021_14_ DECAP_INV_G12
XG17055 XI6/net014_15_ XI6/net021_15_ DECAP_INV_G12
XG17056 XI6/net021_0_ ysel_15_ DECAP_INV_G24
XG17057 XI6/net021_1_ ysel_14_ DECAP_INV_G24
XG17058 XI6/net021_2_ ysel_13_ DECAP_INV_G24
XG17059 XI6/net021_3_ ysel_12_ DECAP_INV_G24
XG17060 XI6/net021_4_ ysel_11_ DECAP_INV_G24
XG17061 XI6/net021_5_ ysel_10_ DECAP_INV_G24
XG17062 XI6/net021_6_ ysel_9_ DECAP_INV_G24
XG17063 XI6/net021_7_ ysel_8_ DECAP_INV_G24
XG17064 XI6/net021_8_ ysel_7_ DECAP_INV_G24
XG17065 XI6/net021_9_ ysel_6_ DECAP_INV_G24
XG17066 XI6/net021_10_ ysel_5_ DECAP_INV_G24
XG17067 XI6/net021_11_ ysel_4_ DECAP_INV_G24
XG17068 XI6/net021_12_ ysel_3_ DECAP_INV_G24
XG17069 XI6/net021_13_ ysel_2_ DECAP_INV_G24
XG17070 XI6/net021_14_ ysel_1_ DECAP_INV_G24
XG17071 XI6/net021_15_ ysel_0_ DECAP_INV_G24
.ENDS


