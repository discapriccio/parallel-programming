.SUBCKT ram DOUT_7_  DOUT_6_  DOUT_5_  DOUT_4_  DOUT_3_  DOUT_2_  DOUT_1_  DOUT_0_  A_9_  A_8_  A_7_  A_6_  A_5_  A_4_  A_3_  A_2_  A_1_  A_0_  CLK  CS  DIN_7_  DIN_6_  DIN_5_  DIN_4_  DIN_3_  DIN_2_  DIN_1_  DIN_0_  RD  WR  gnd  vdd  
XI11_7/XI2/MN0_15 XI11_7/net21_0_ ysel_15_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll]
XI11_7/XI2/MN0_14 XI11_7/net21_1_ ysel_14_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_13 XI11_7/net21_2_ ysel_13_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_12 XI11_7/net21_3_ ysel_12_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_11 XI11_7/net21_4_ ysel_11_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_10 XI11_7/net21_5_ ysel_10_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_9 XI11_7/net21_6_ ysel_9_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_8 XI11_7/net21_7_ ysel_8_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_7 XI11_7/net21_8_ ysel_7_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_6 XI11_7/net21_9_ ysel_6_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_5 XI11_7/net21_10_ ysel_5_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_4 XI11_7/net21_11_ ysel_4_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_3 XI11_7/net21_12_ ysel_3_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_2 XI11_7/net21_13_ ysel_2_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_1 XI11_7/net21_14_ ysel_1_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN0_0 XI11_7/net21_15_ ysel_0_ XI11_7/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_15 XI11_7/net20_0_ ysel_15_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_14 XI11_7/net20_1_ ysel_14_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_13 XI11_7/net20_2_ ysel_13_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_12 XI11_7/net20_3_ ysel_12_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_11 XI11_7/net20_4_ ysel_11_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_10 XI11_7/net20_5_ ysel_10_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_9 XI11_7/net20_6_ ysel_9_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_8 XI11_7/net20_7_ ysel_8_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_7 XI11_7/net20_8_ ysel_7_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_6 XI11_7/net20_9_ ysel_6_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_5 XI11_7/net20_10_ ysel_5_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_4 XI11_7/net20_11_ ysel_4_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_3 XI11_7/net20_12_ ysel_3_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_2 XI11_7/net20_13_ ysel_2_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_1 XI11_7/net20_14_ ysel_1_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI2/MN1_0 XI11_7/net20_15_ ysel_0_ XI11_7/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_7/XI4/MN8 vdd XI11_7/XI4/net8 XI11_7/net12 vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_7/XI4/MP0 XI11_7/net9 XI11_7/XI4/net23 vdd vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_7/XI4/MP4 XI11_7/net12 XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI4/MP1 XI11_7/net9 XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI4/MP5 XI11_7/net12 XI11_7/preck XI11_7/net9 vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI4/MN7 vdd XI11_7/XI4/net090 DOUT_7_ vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_7/XI4/MP3 gnd XI11_7/XI4/net089 XI11_7/net12 gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_7/XI4/MN5 XI11_7/net9 XI11_7/XI4/net0103 gnd gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_7/XI4/MN4 XI11_7/XI4/data_out_ XI11_7/XI4/net32 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_7/XI4/MN0 XI11_7/XI4/data_out XI11_7/XI4/net52 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_7/XI4/MN9 gnd XI11_7/XI4/net0112 DOUT_7_ gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_7/XI1_15/MP2 XI11_7/net20_0_ XI11_7/preck XI11_7/net21_0_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_15/MP1 XI11_7/net20_0_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_15/MP0 XI11_7/net21_0_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_14/MP2 XI11_7/net20_1_ XI11_7/preck XI11_7/net21_1_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_14/MP1 XI11_7/net20_1_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_14/MP0 XI11_7/net21_1_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_13/MP2 XI11_7/net20_2_ XI11_7/preck XI11_7/net21_2_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_13/MP1 XI11_7/net20_2_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_13/MP0 XI11_7/net21_2_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_12/MP2 XI11_7/net20_3_ XI11_7/preck XI11_7/net21_3_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_12/MP1 XI11_7/net20_3_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_12/MP0 XI11_7/net21_3_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_11/MP2 XI11_7/net20_4_ XI11_7/preck XI11_7/net21_4_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_11/MP1 XI11_7/net20_4_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_11/MP0 XI11_7/net21_4_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_10/MP2 XI11_7/net20_5_ XI11_7/preck XI11_7/net21_5_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_10/MP1 XI11_7/net20_5_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_10/MP0 XI11_7/net21_5_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_9/MP2 XI11_7/net20_6_ XI11_7/preck XI11_7/net21_6_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_9/MP1 XI11_7/net20_6_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_9/MP0 XI11_7/net21_6_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_8/MP2 XI11_7/net20_7_ XI11_7/preck XI11_7/net21_7_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_8/MP1 XI11_7/net20_7_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_8/MP0 XI11_7/net21_7_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_7/MP2 XI11_7/net20_8_ XI11_7/preck XI11_7/net21_8_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_7/MP1 XI11_7/net20_8_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_7/MP0 XI11_7/net21_8_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_6/MP2 XI11_7/net20_9_ XI11_7/preck XI11_7/net21_9_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_6/MP1 XI11_7/net20_9_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_6/MP0 XI11_7/net21_9_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_5/MP2 XI11_7/net20_10_ XI11_7/preck XI11_7/net21_10_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_5/MP1 XI11_7/net20_10_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_5/MP0 XI11_7/net21_10_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_4/MP2 XI11_7/net20_11_ XI11_7/preck XI11_7/net21_11_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_4/MP1 XI11_7/net20_11_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_4/MP0 XI11_7/net21_11_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_3/MP2 XI11_7/net20_12_ XI11_7/preck XI11_7/net21_12_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_3/MP1 XI11_7/net20_12_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_3/MP0 XI11_7/net21_12_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_2/MP2 XI11_7/net20_13_ XI11_7/preck XI11_7/net21_13_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_2/MP1 XI11_7/net20_13_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_2/MP0 XI11_7/net21_13_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_1/MP2 XI11_7/net20_14_ XI11_7/preck XI11_7/net21_14_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_1/MP1 XI11_7/net20_14_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_1/MP0 XI11_7/net21_14_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_0/MP2 XI11_7/net20_15_ XI11_7/preck XI11_7/net21_15_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_7/XI1_0/MP1 XI11_7/net20_15_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI1_0/MP0 XI11_7/net21_15_ XI11_7/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_7/XI0/MN0_15 gnd gnd XI11_7/net21_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_14 gnd gnd XI11_7/net21_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_13 gnd gnd XI11_7/net21_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_12 gnd gnd XI11_7/net21_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_11 gnd gnd XI11_7/net21_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_10 gnd gnd XI11_7/net21_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_9 gnd gnd XI11_7/net21_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_8 gnd gnd XI11_7/net21_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_7 gnd gnd XI11_7/net21_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_6 gnd gnd XI11_7/net21_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_5 gnd gnd XI11_7/net21_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_4 gnd gnd XI11_7/net21_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_3 gnd gnd XI11_7/net21_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_2 gnd gnd XI11_7/net21_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_1 gnd gnd XI11_7/net21_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN0_0 gnd gnd XI11_7/net21_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_15 gnd gnd XI11_7/net20_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_14 gnd gnd XI11_7/net20_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_13 gnd gnd XI11_7/net20_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_12 gnd gnd XI11_7/net20_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_11 gnd gnd XI11_7/net20_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_10 gnd gnd XI11_7/net20_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_9 gnd gnd XI11_7/net20_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_8 gnd gnd XI11_7/net20_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_7 gnd gnd XI11_7/net20_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_6 gnd gnd XI11_7/net20_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_5 gnd gnd XI11_7/net20_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_4 gnd gnd XI11_7/net20_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_3 gnd gnd XI11_7/net20_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_2 gnd gnd XI11_7/net20_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_1 gnd gnd XI11_7/net20_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/MN1_0 gnd gnd XI11_7/net20_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_15 XI11_7/net21_0_ xsel_63_ XI11_7/XI0/XI0_63/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_14 XI11_7/net21_1_ xsel_63_ XI11_7/XI0/XI0_63/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_13 XI11_7/net21_2_ xsel_63_ XI11_7/XI0/XI0_63/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_12 XI11_7/net21_3_ xsel_63_ XI11_7/XI0/XI0_63/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_11 XI11_7/net21_4_ xsel_63_ XI11_7/XI0/XI0_63/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_10 XI11_7/net21_5_ xsel_63_ XI11_7/XI0/XI0_63/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_9 XI11_7/net21_6_ xsel_63_ XI11_7/XI0/XI0_63/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_8 XI11_7/net21_7_ xsel_63_ XI11_7/XI0/XI0_63/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_7 XI11_7/net21_8_ xsel_63_ XI11_7/XI0/XI0_63/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_6 XI11_7/net21_9_ xsel_63_ XI11_7/XI0/XI0_63/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_5 XI11_7/net21_10_ xsel_63_ XI11_7/XI0/XI0_63/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_4 XI11_7/net21_11_ xsel_63_ XI11_7/XI0/XI0_63/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_3 XI11_7/net21_12_ xsel_63_ XI11_7/XI0/XI0_63/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_2 XI11_7/net21_13_ xsel_63_ XI11_7/XI0/XI0_63/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_1 XI11_7/net21_14_ xsel_63_ XI11_7/XI0/XI0_63/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN0_0 XI11_7/net21_15_ xsel_63_ XI11_7/XI0/XI0_63/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_15 XI11_7/XI0/XI0_63/d__15_ xsel_63_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_14 XI11_7/XI0/XI0_63/d__14_ xsel_63_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_13 XI11_7/XI0/XI0_63/d__13_ xsel_63_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_12 XI11_7/XI0/XI0_63/d__12_ xsel_63_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_11 XI11_7/XI0/XI0_63/d__11_ xsel_63_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_10 XI11_7/XI0/XI0_63/d__10_ xsel_63_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_9 XI11_7/XI0/XI0_63/d__9_ xsel_63_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_8 XI11_7/XI0/XI0_63/d__8_ xsel_63_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_7 XI11_7/XI0/XI0_63/d__7_ xsel_63_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_6 XI11_7/XI0/XI0_63/d__6_ xsel_63_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_5 XI11_7/XI0/XI0_63/d__5_ xsel_63_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_4 XI11_7/XI0/XI0_63/d__4_ xsel_63_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_3 XI11_7/XI0/XI0_63/d__3_ xsel_63_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_2 XI11_7/XI0/XI0_63/d__2_ xsel_63_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_1 XI11_7/XI0/XI0_63/d__1_ xsel_63_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_63/MN1_0 XI11_7/XI0/XI0_63/d__0_ xsel_63_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_15 XI11_7/net21_0_ xsel_62_ XI11_7/XI0/XI0_62/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_14 XI11_7/net21_1_ xsel_62_ XI11_7/XI0/XI0_62/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_13 XI11_7/net21_2_ xsel_62_ XI11_7/XI0/XI0_62/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_12 XI11_7/net21_3_ xsel_62_ XI11_7/XI0/XI0_62/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_11 XI11_7/net21_4_ xsel_62_ XI11_7/XI0/XI0_62/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_10 XI11_7/net21_5_ xsel_62_ XI11_7/XI0/XI0_62/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_9 XI11_7/net21_6_ xsel_62_ XI11_7/XI0/XI0_62/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_8 XI11_7/net21_7_ xsel_62_ XI11_7/XI0/XI0_62/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_7 XI11_7/net21_8_ xsel_62_ XI11_7/XI0/XI0_62/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_6 XI11_7/net21_9_ xsel_62_ XI11_7/XI0/XI0_62/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_5 XI11_7/net21_10_ xsel_62_ XI11_7/XI0/XI0_62/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_4 XI11_7/net21_11_ xsel_62_ XI11_7/XI0/XI0_62/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_3 XI11_7/net21_12_ xsel_62_ XI11_7/XI0/XI0_62/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_2 XI11_7/net21_13_ xsel_62_ XI11_7/XI0/XI0_62/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_1 XI11_7/net21_14_ xsel_62_ XI11_7/XI0/XI0_62/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN0_0 XI11_7/net21_15_ xsel_62_ XI11_7/XI0/XI0_62/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_15 XI11_7/XI0/XI0_62/d__15_ xsel_62_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_14 XI11_7/XI0/XI0_62/d__14_ xsel_62_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_13 XI11_7/XI0/XI0_62/d__13_ xsel_62_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_12 XI11_7/XI0/XI0_62/d__12_ xsel_62_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_11 XI11_7/XI0/XI0_62/d__11_ xsel_62_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_10 XI11_7/XI0/XI0_62/d__10_ xsel_62_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_9 XI11_7/XI0/XI0_62/d__9_ xsel_62_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_8 XI11_7/XI0/XI0_62/d__8_ xsel_62_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_7 XI11_7/XI0/XI0_62/d__7_ xsel_62_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_6 XI11_7/XI0/XI0_62/d__6_ xsel_62_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_5 XI11_7/XI0/XI0_62/d__5_ xsel_62_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_4 XI11_7/XI0/XI0_62/d__4_ xsel_62_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_3 XI11_7/XI0/XI0_62/d__3_ xsel_62_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_2 XI11_7/XI0/XI0_62/d__2_ xsel_62_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_1 XI11_7/XI0/XI0_62/d__1_ xsel_62_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_62/MN1_0 XI11_7/XI0/XI0_62/d__0_ xsel_62_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_15 XI11_7/net21_0_ xsel_61_ XI11_7/XI0/XI0_61/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_14 XI11_7/net21_1_ xsel_61_ XI11_7/XI0/XI0_61/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_13 XI11_7/net21_2_ xsel_61_ XI11_7/XI0/XI0_61/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_12 XI11_7/net21_3_ xsel_61_ XI11_7/XI0/XI0_61/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_11 XI11_7/net21_4_ xsel_61_ XI11_7/XI0/XI0_61/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_10 XI11_7/net21_5_ xsel_61_ XI11_7/XI0/XI0_61/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_9 XI11_7/net21_6_ xsel_61_ XI11_7/XI0/XI0_61/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_8 XI11_7/net21_7_ xsel_61_ XI11_7/XI0/XI0_61/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_7 XI11_7/net21_8_ xsel_61_ XI11_7/XI0/XI0_61/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_6 XI11_7/net21_9_ xsel_61_ XI11_7/XI0/XI0_61/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_5 XI11_7/net21_10_ xsel_61_ XI11_7/XI0/XI0_61/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_4 XI11_7/net21_11_ xsel_61_ XI11_7/XI0/XI0_61/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_3 XI11_7/net21_12_ xsel_61_ XI11_7/XI0/XI0_61/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_2 XI11_7/net21_13_ xsel_61_ XI11_7/XI0/XI0_61/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_1 XI11_7/net21_14_ xsel_61_ XI11_7/XI0/XI0_61/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN0_0 XI11_7/net21_15_ xsel_61_ XI11_7/XI0/XI0_61/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_15 XI11_7/XI0/XI0_61/d__15_ xsel_61_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_14 XI11_7/XI0/XI0_61/d__14_ xsel_61_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_13 XI11_7/XI0/XI0_61/d__13_ xsel_61_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_12 XI11_7/XI0/XI0_61/d__12_ xsel_61_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_11 XI11_7/XI0/XI0_61/d__11_ xsel_61_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_10 XI11_7/XI0/XI0_61/d__10_ xsel_61_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_9 XI11_7/XI0/XI0_61/d__9_ xsel_61_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_8 XI11_7/XI0/XI0_61/d__8_ xsel_61_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_7 XI11_7/XI0/XI0_61/d__7_ xsel_61_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_6 XI11_7/XI0/XI0_61/d__6_ xsel_61_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_5 XI11_7/XI0/XI0_61/d__5_ xsel_61_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_4 XI11_7/XI0/XI0_61/d__4_ xsel_61_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_3 XI11_7/XI0/XI0_61/d__3_ xsel_61_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_2 XI11_7/XI0/XI0_61/d__2_ xsel_61_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_1 XI11_7/XI0/XI0_61/d__1_ xsel_61_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_61/MN1_0 XI11_7/XI0/XI0_61/d__0_ xsel_61_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_15 XI11_7/net21_0_ xsel_60_ XI11_7/XI0/XI0_60/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_14 XI11_7/net21_1_ xsel_60_ XI11_7/XI0/XI0_60/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_13 XI11_7/net21_2_ xsel_60_ XI11_7/XI0/XI0_60/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_12 XI11_7/net21_3_ xsel_60_ XI11_7/XI0/XI0_60/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_11 XI11_7/net21_4_ xsel_60_ XI11_7/XI0/XI0_60/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_10 XI11_7/net21_5_ xsel_60_ XI11_7/XI0/XI0_60/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_9 XI11_7/net21_6_ xsel_60_ XI11_7/XI0/XI0_60/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_8 XI11_7/net21_7_ xsel_60_ XI11_7/XI0/XI0_60/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_7 XI11_7/net21_8_ xsel_60_ XI11_7/XI0/XI0_60/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_6 XI11_7/net21_9_ xsel_60_ XI11_7/XI0/XI0_60/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_5 XI11_7/net21_10_ xsel_60_ XI11_7/XI0/XI0_60/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_4 XI11_7/net21_11_ xsel_60_ XI11_7/XI0/XI0_60/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_3 XI11_7/net21_12_ xsel_60_ XI11_7/XI0/XI0_60/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_2 XI11_7/net21_13_ xsel_60_ XI11_7/XI0/XI0_60/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_1 XI11_7/net21_14_ xsel_60_ XI11_7/XI0/XI0_60/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN0_0 XI11_7/net21_15_ xsel_60_ XI11_7/XI0/XI0_60/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_15 XI11_7/XI0/XI0_60/d__15_ xsel_60_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_14 XI11_7/XI0/XI0_60/d__14_ xsel_60_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_13 XI11_7/XI0/XI0_60/d__13_ xsel_60_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_12 XI11_7/XI0/XI0_60/d__12_ xsel_60_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_11 XI11_7/XI0/XI0_60/d__11_ xsel_60_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_10 XI11_7/XI0/XI0_60/d__10_ xsel_60_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_9 XI11_7/XI0/XI0_60/d__9_ xsel_60_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_8 XI11_7/XI0/XI0_60/d__8_ xsel_60_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_7 XI11_7/XI0/XI0_60/d__7_ xsel_60_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_6 XI11_7/XI0/XI0_60/d__6_ xsel_60_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_5 XI11_7/XI0/XI0_60/d__5_ xsel_60_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_4 XI11_7/XI0/XI0_60/d__4_ xsel_60_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_3 XI11_7/XI0/XI0_60/d__3_ xsel_60_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_2 XI11_7/XI0/XI0_60/d__2_ xsel_60_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_1 XI11_7/XI0/XI0_60/d__1_ xsel_60_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_60/MN1_0 XI11_7/XI0/XI0_60/d__0_ xsel_60_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_15 XI11_7/net21_0_ xsel_59_ XI11_7/XI0/XI0_59/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_14 XI11_7/net21_1_ xsel_59_ XI11_7/XI0/XI0_59/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_13 XI11_7/net21_2_ xsel_59_ XI11_7/XI0/XI0_59/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_12 XI11_7/net21_3_ xsel_59_ XI11_7/XI0/XI0_59/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_11 XI11_7/net21_4_ xsel_59_ XI11_7/XI0/XI0_59/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_10 XI11_7/net21_5_ xsel_59_ XI11_7/XI0/XI0_59/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_9 XI11_7/net21_6_ xsel_59_ XI11_7/XI0/XI0_59/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_8 XI11_7/net21_7_ xsel_59_ XI11_7/XI0/XI0_59/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_7 XI11_7/net21_8_ xsel_59_ XI11_7/XI0/XI0_59/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_6 XI11_7/net21_9_ xsel_59_ XI11_7/XI0/XI0_59/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_5 XI11_7/net21_10_ xsel_59_ XI11_7/XI0/XI0_59/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_4 XI11_7/net21_11_ xsel_59_ XI11_7/XI0/XI0_59/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_3 XI11_7/net21_12_ xsel_59_ XI11_7/XI0/XI0_59/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_2 XI11_7/net21_13_ xsel_59_ XI11_7/XI0/XI0_59/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_1 XI11_7/net21_14_ xsel_59_ XI11_7/XI0/XI0_59/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN0_0 XI11_7/net21_15_ xsel_59_ XI11_7/XI0/XI0_59/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_15 XI11_7/XI0/XI0_59/d__15_ xsel_59_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_14 XI11_7/XI0/XI0_59/d__14_ xsel_59_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_13 XI11_7/XI0/XI0_59/d__13_ xsel_59_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_12 XI11_7/XI0/XI0_59/d__12_ xsel_59_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_11 XI11_7/XI0/XI0_59/d__11_ xsel_59_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_10 XI11_7/XI0/XI0_59/d__10_ xsel_59_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_9 XI11_7/XI0/XI0_59/d__9_ xsel_59_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_8 XI11_7/XI0/XI0_59/d__8_ xsel_59_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_7 XI11_7/XI0/XI0_59/d__7_ xsel_59_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_6 XI11_7/XI0/XI0_59/d__6_ xsel_59_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_5 XI11_7/XI0/XI0_59/d__5_ xsel_59_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_4 XI11_7/XI0/XI0_59/d__4_ xsel_59_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_3 XI11_7/XI0/XI0_59/d__3_ xsel_59_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_2 XI11_7/XI0/XI0_59/d__2_ xsel_59_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_1 XI11_7/XI0/XI0_59/d__1_ xsel_59_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_59/MN1_0 XI11_7/XI0/XI0_59/d__0_ xsel_59_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_15 XI11_7/net21_0_ xsel_58_ XI11_7/XI0/XI0_58/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_14 XI11_7/net21_1_ xsel_58_ XI11_7/XI0/XI0_58/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_13 XI11_7/net21_2_ xsel_58_ XI11_7/XI0/XI0_58/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_12 XI11_7/net21_3_ xsel_58_ XI11_7/XI0/XI0_58/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_11 XI11_7/net21_4_ xsel_58_ XI11_7/XI0/XI0_58/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_10 XI11_7/net21_5_ xsel_58_ XI11_7/XI0/XI0_58/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_9 XI11_7/net21_6_ xsel_58_ XI11_7/XI0/XI0_58/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_8 XI11_7/net21_7_ xsel_58_ XI11_7/XI0/XI0_58/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_7 XI11_7/net21_8_ xsel_58_ XI11_7/XI0/XI0_58/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_6 XI11_7/net21_9_ xsel_58_ XI11_7/XI0/XI0_58/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_5 XI11_7/net21_10_ xsel_58_ XI11_7/XI0/XI0_58/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_4 XI11_7/net21_11_ xsel_58_ XI11_7/XI0/XI0_58/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_3 XI11_7/net21_12_ xsel_58_ XI11_7/XI0/XI0_58/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_2 XI11_7/net21_13_ xsel_58_ XI11_7/XI0/XI0_58/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_1 XI11_7/net21_14_ xsel_58_ XI11_7/XI0/XI0_58/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN0_0 XI11_7/net21_15_ xsel_58_ XI11_7/XI0/XI0_58/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_15 XI11_7/XI0/XI0_58/d__15_ xsel_58_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_14 XI11_7/XI0/XI0_58/d__14_ xsel_58_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_13 XI11_7/XI0/XI0_58/d__13_ xsel_58_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_12 XI11_7/XI0/XI0_58/d__12_ xsel_58_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_11 XI11_7/XI0/XI0_58/d__11_ xsel_58_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_10 XI11_7/XI0/XI0_58/d__10_ xsel_58_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_9 XI11_7/XI0/XI0_58/d__9_ xsel_58_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_8 XI11_7/XI0/XI0_58/d__8_ xsel_58_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_7 XI11_7/XI0/XI0_58/d__7_ xsel_58_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_6 XI11_7/XI0/XI0_58/d__6_ xsel_58_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_5 XI11_7/XI0/XI0_58/d__5_ xsel_58_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_4 XI11_7/XI0/XI0_58/d__4_ xsel_58_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_3 XI11_7/XI0/XI0_58/d__3_ xsel_58_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_2 XI11_7/XI0/XI0_58/d__2_ xsel_58_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_1 XI11_7/XI0/XI0_58/d__1_ xsel_58_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_58/MN1_0 XI11_7/XI0/XI0_58/d__0_ xsel_58_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_15 XI11_7/net21_0_ xsel_57_ XI11_7/XI0/XI0_57/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_14 XI11_7/net21_1_ xsel_57_ XI11_7/XI0/XI0_57/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_13 XI11_7/net21_2_ xsel_57_ XI11_7/XI0/XI0_57/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_12 XI11_7/net21_3_ xsel_57_ XI11_7/XI0/XI0_57/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_11 XI11_7/net21_4_ xsel_57_ XI11_7/XI0/XI0_57/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_10 XI11_7/net21_5_ xsel_57_ XI11_7/XI0/XI0_57/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_9 XI11_7/net21_6_ xsel_57_ XI11_7/XI0/XI0_57/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_8 XI11_7/net21_7_ xsel_57_ XI11_7/XI0/XI0_57/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_7 XI11_7/net21_8_ xsel_57_ XI11_7/XI0/XI0_57/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_6 XI11_7/net21_9_ xsel_57_ XI11_7/XI0/XI0_57/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_5 XI11_7/net21_10_ xsel_57_ XI11_7/XI0/XI0_57/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_4 XI11_7/net21_11_ xsel_57_ XI11_7/XI0/XI0_57/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_3 XI11_7/net21_12_ xsel_57_ XI11_7/XI0/XI0_57/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_2 XI11_7/net21_13_ xsel_57_ XI11_7/XI0/XI0_57/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_1 XI11_7/net21_14_ xsel_57_ XI11_7/XI0/XI0_57/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN0_0 XI11_7/net21_15_ xsel_57_ XI11_7/XI0/XI0_57/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_15 XI11_7/XI0/XI0_57/d__15_ xsel_57_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_14 XI11_7/XI0/XI0_57/d__14_ xsel_57_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_13 XI11_7/XI0/XI0_57/d__13_ xsel_57_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_12 XI11_7/XI0/XI0_57/d__12_ xsel_57_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_11 XI11_7/XI0/XI0_57/d__11_ xsel_57_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_10 XI11_7/XI0/XI0_57/d__10_ xsel_57_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_9 XI11_7/XI0/XI0_57/d__9_ xsel_57_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_8 XI11_7/XI0/XI0_57/d__8_ xsel_57_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_7 XI11_7/XI0/XI0_57/d__7_ xsel_57_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_6 XI11_7/XI0/XI0_57/d__6_ xsel_57_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_5 XI11_7/XI0/XI0_57/d__5_ xsel_57_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_4 XI11_7/XI0/XI0_57/d__4_ xsel_57_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_3 XI11_7/XI0/XI0_57/d__3_ xsel_57_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_2 XI11_7/XI0/XI0_57/d__2_ xsel_57_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_1 XI11_7/XI0/XI0_57/d__1_ xsel_57_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_57/MN1_0 XI11_7/XI0/XI0_57/d__0_ xsel_57_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_15 XI11_7/net21_0_ xsel_56_ XI11_7/XI0/XI0_56/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_14 XI11_7/net21_1_ xsel_56_ XI11_7/XI0/XI0_56/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_13 XI11_7/net21_2_ xsel_56_ XI11_7/XI0/XI0_56/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_12 XI11_7/net21_3_ xsel_56_ XI11_7/XI0/XI0_56/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_11 XI11_7/net21_4_ xsel_56_ XI11_7/XI0/XI0_56/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_10 XI11_7/net21_5_ xsel_56_ XI11_7/XI0/XI0_56/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_9 XI11_7/net21_6_ xsel_56_ XI11_7/XI0/XI0_56/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_8 XI11_7/net21_7_ xsel_56_ XI11_7/XI0/XI0_56/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_7 XI11_7/net21_8_ xsel_56_ XI11_7/XI0/XI0_56/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_6 XI11_7/net21_9_ xsel_56_ XI11_7/XI0/XI0_56/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_5 XI11_7/net21_10_ xsel_56_ XI11_7/XI0/XI0_56/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_4 XI11_7/net21_11_ xsel_56_ XI11_7/XI0/XI0_56/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_3 XI11_7/net21_12_ xsel_56_ XI11_7/XI0/XI0_56/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_2 XI11_7/net21_13_ xsel_56_ XI11_7/XI0/XI0_56/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_1 XI11_7/net21_14_ xsel_56_ XI11_7/XI0/XI0_56/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN0_0 XI11_7/net21_15_ xsel_56_ XI11_7/XI0/XI0_56/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_15 XI11_7/XI0/XI0_56/d__15_ xsel_56_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_14 XI11_7/XI0/XI0_56/d__14_ xsel_56_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_13 XI11_7/XI0/XI0_56/d__13_ xsel_56_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_12 XI11_7/XI0/XI0_56/d__12_ xsel_56_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_11 XI11_7/XI0/XI0_56/d__11_ xsel_56_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_10 XI11_7/XI0/XI0_56/d__10_ xsel_56_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_9 XI11_7/XI0/XI0_56/d__9_ xsel_56_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_8 XI11_7/XI0/XI0_56/d__8_ xsel_56_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_7 XI11_7/XI0/XI0_56/d__7_ xsel_56_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_6 XI11_7/XI0/XI0_56/d__6_ xsel_56_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_5 XI11_7/XI0/XI0_56/d__5_ xsel_56_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_4 XI11_7/XI0/XI0_56/d__4_ xsel_56_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_3 XI11_7/XI0/XI0_56/d__3_ xsel_56_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_2 XI11_7/XI0/XI0_56/d__2_ xsel_56_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_1 XI11_7/XI0/XI0_56/d__1_ xsel_56_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_56/MN1_0 XI11_7/XI0/XI0_56/d__0_ xsel_56_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_15 XI11_7/net21_0_ xsel_55_ XI11_7/XI0/XI0_55/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_14 XI11_7/net21_1_ xsel_55_ XI11_7/XI0/XI0_55/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_13 XI11_7/net21_2_ xsel_55_ XI11_7/XI0/XI0_55/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_12 XI11_7/net21_3_ xsel_55_ XI11_7/XI0/XI0_55/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_11 XI11_7/net21_4_ xsel_55_ XI11_7/XI0/XI0_55/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_10 XI11_7/net21_5_ xsel_55_ XI11_7/XI0/XI0_55/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_9 XI11_7/net21_6_ xsel_55_ XI11_7/XI0/XI0_55/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_8 XI11_7/net21_7_ xsel_55_ XI11_7/XI0/XI0_55/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_7 XI11_7/net21_8_ xsel_55_ XI11_7/XI0/XI0_55/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_6 XI11_7/net21_9_ xsel_55_ XI11_7/XI0/XI0_55/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_5 XI11_7/net21_10_ xsel_55_ XI11_7/XI0/XI0_55/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_4 XI11_7/net21_11_ xsel_55_ XI11_7/XI0/XI0_55/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_3 XI11_7/net21_12_ xsel_55_ XI11_7/XI0/XI0_55/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_2 XI11_7/net21_13_ xsel_55_ XI11_7/XI0/XI0_55/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_1 XI11_7/net21_14_ xsel_55_ XI11_7/XI0/XI0_55/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN0_0 XI11_7/net21_15_ xsel_55_ XI11_7/XI0/XI0_55/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_15 XI11_7/XI0/XI0_55/d__15_ xsel_55_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_14 XI11_7/XI0/XI0_55/d__14_ xsel_55_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_13 XI11_7/XI0/XI0_55/d__13_ xsel_55_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_12 XI11_7/XI0/XI0_55/d__12_ xsel_55_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_11 XI11_7/XI0/XI0_55/d__11_ xsel_55_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_10 XI11_7/XI0/XI0_55/d__10_ xsel_55_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_9 XI11_7/XI0/XI0_55/d__9_ xsel_55_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_8 XI11_7/XI0/XI0_55/d__8_ xsel_55_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_7 XI11_7/XI0/XI0_55/d__7_ xsel_55_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_6 XI11_7/XI0/XI0_55/d__6_ xsel_55_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_5 XI11_7/XI0/XI0_55/d__5_ xsel_55_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_4 XI11_7/XI0/XI0_55/d__4_ xsel_55_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_3 XI11_7/XI0/XI0_55/d__3_ xsel_55_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_2 XI11_7/XI0/XI0_55/d__2_ xsel_55_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_1 XI11_7/XI0/XI0_55/d__1_ xsel_55_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_55/MN1_0 XI11_7/XI0/XI0_55/d__0_ xsel_55_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_15 XI11_7/net21_0_ xsel_54_ XI11_7/XI0/XI0_54/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_14 XI11_7/net21_1_ xsel_54_ XI11_7/XI0/XI0_54/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_13 XI11_7/net21_2_ xsel_54_ XI11_7/XI0/XI0_54/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_12 XI11_7/net21_3_ xsel_54_ XI11_7/XI0/XI0_54/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_11 XI11_7/net21_4_ xsel_54_ XI11_7/XI0/XI0_54/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_10 XI11_7/net21_5_ xsel_54_ XI11_7/XI0/XI0_54/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_9 XI11_7/net21_6_ xsel_54_ XI11_7/XI0/XI0_54/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_8 XI11_7/net21_7_ xsel_54_ XI11_7/XI0/XI0_54/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_7 XI11_7/net21_8_ xsel_54_ XI11_7/XI0/XI0_54/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_6 XI11_7/net21_9_ xsel_54_ XI11_7/XI0/XI0_54/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_5 XI11_7/net21_10_ xsel_54_ XI11_7/XI0/XI0_54/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_4 XI11_7/net21_11_ xsel_54_ XI11_7/XI0/XI0_54/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_3 XI11_7/net21_12_ xsel_54_ XI11_7/XI0/XI0_54/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_2 XI11_7/net21_13_ xsel_54_ XI11_7/XI0/XI0_54/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_1 XI11_7/net21_14_ xsel_54_ XI11_7/XI0/XI0_54/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN0_0 XI11_7/net21_15_ xsel_54_ XI11_7/XI0/XI0_54/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_15 XI11_7/XI0/XI0_54/d__15_ xsel_54_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_14 XI11_7/XI0/XI0_54/d__14_ xsel_54_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_13 XI11_7/XI0/XI0_54/d__13_ xsel_54_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_12 XI11_7/XI0/XI0_54/d__12_ xsel_54_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_11 XI11_7/XI0/XI0_54/d__11_ xsel_54_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_10 XI11_7/XI0/XI0_54/d__10_ xsel_54_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_9 XI11_7/XI0/XI0_54/d__9_ xsel_54_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_8 XI11_7/XI0/XI0_54/d__8_ xsel_54_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_7 XI11_7/XI0/XI0_54/d__7_ xsel_54_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_6 XI11_7/XI0/XI0_54/d__6_ xsel_54_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_5 XI11_7/XI0/XI0_54/d__5_ xsel_54_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_4 XI11_7/XI0/XI0_54/d__4_ xsel_54_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_3 XI11_7/XI0/XI0_54/d__3_ xsel_54_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_2 XI11_7/XI0/XI0_54/d__2_ xsel_54_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_1 XI11_7/XI0/XI0_54/d__1_ xsel_54_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_54/MN1_0 XI11_7/XI0/XI0_54/d__0_ xsel_54_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_15 XI11_7/net21_0_ xsel_53_ XI11_7/XI0/XI0_53/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_14 XI11_7/net21_1_ xsel_53_ XI11_7/XI0/XI0_53/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_13 XI11_7/net21_2_ xsel_53_ XI11_7/XI0/XI0_53/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_12 XI11_7/net21_3_ xsel_53_ XI11_7/XI0/XI0_53/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_11 XI11_7/net21_4_ xsel_53_ XI11_7/XI0/XI0_53/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_10 XI11_7/net21_5_ xsel_53_ XI11_7/XI0/XI0_53/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_9 XI11_7/net21_6_ xsel_53_ XI11_7/XI0/XI0_53/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_8 XI11_7/net21_7_ xsel_53_ XI11_7/XI0/XI0_53/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_7 XI11_7/net21_8_ xsel_53_ XI11_7/XI0/XI0_53/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_6 XI11_7/net21_9_ xsel_53_ XI11_7/XI0/XI0_53/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_5 XI11_7/net21_10_ xsel_53_ XI11_7/XI0/XI0_53/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_4 XI11_7/net21_11_ xsel_53_ XI11_7/XI0/XI0_53/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_3 XI11_7/net21_12_ xsel_53_ XI11_7/XI0/XI0_53/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_2 XI11_7/net21_13_ xsel_53_ XI11_7/XI0/XI0_53/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_1 XI11_7/net21_14_ xsel_53_ XI11_7/XI0/XI0_53/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN0_0 XI11_7/net21_15_ xsel_53_ XI11_7/XI0/XI0_53/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_15 XI11_7/XI0/XI0_53/d__15_ xsel_53_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_14 XI11_7/XI0/XI0_53/d__14_ xsel_53_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_13 XI11_7/XI0/XI0_53/d__13_ xsel_53_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_12 XI11_7/XI0/XI0_53/d__12_ xsel_53_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_11 XI11_7/XI0/XI0_53/d__11_ xsel_53_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_10 XI11_7/XI0/XI0_53/d__10_ xsel_53_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_9 XI11_7/XI0/XI0_53/d__9_ xsel_53_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_8 XI11_7/XI0/XI0_53/d__8_ xsel_53_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_7 XI11_7/XI0/XI0_53/d__7_ xsel_53_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_6 XI11_7/XI0/XI0_53/d__6_ xsel_53_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_5 XI11_7/XI0/XI0_53/d__5_ xsel_53_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_4 XI11_7/XI0/XI0_53/d__4_ xsel_53_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_3 XI11_7/XI0/XI0_53/d__3_ xsel_53_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_2 XI11_7/XI0/XI0_53/d__2_ xsel_53_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_1 XI11_7/XI0/XI0_53/d__1_ xsel_53_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_53/MN1_0 XI11_7/XI0/XI0_53/d__0_ xsel_53_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_15 XI11_7/net21_0_ xsel_52_ XI11_7/XI0/XI0_52/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_14 XI11_7/net21_1_ xsel_52_ XI11_7/XI0/XI0_52/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_13 XI11_7/net21_2_ xsel_52_ XI11_7/XI0/XI0_52/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_12 XI11_7/net21_3_ xsel_52_ XI11_7/XI0/XI0_52/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_11 XI11_7/net21_4_ xsel_52_ XI11_7/XI0/XI0_52/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_10 XI11_7/net21_5_ xsel_52_ XI11_7/XI0/XI0_52/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_9 XI11_7/net21_6_ xsel_52_ XI11_7/XI0/XI0_52/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_8 XI11_7/net21_7_ xsel_52_ XI11_7/XI0/XI0_52/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_7 XI11_7/net21_8_ xsel_52_ XI11_7/XI0/XI0_52/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_6 XI11_7/net21_9_ xsel_52_ XI11_7/XI0/XI0_52/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_5 XI11_7/net21_10_ xsel_52_ XI11_7/XI0/XI0_52/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_4 XI11_7/net21_11_ xsel_52_ XI11_7/XI0/XI0_52/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_3 XI11_7/net21_12_ xsel_52_ XI11_7/XI0/XI0_52/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_2 XI11_7/net21_13_ xsel_52_ XI11_7/XI0/XI0_52/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_1 XI11_7/net21_14_ xsel_52_ XI11_7/XI0/XI0_52/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN0_0 XI11_7/net21_15_ xsel_52_ XI11_7/XI0/XI0_52/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_15 XI11_7/XI0/XI0_52/d__15_ xsel_52_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_14 XI11_7/XI0/XI0_52/d__14_ xsel_52_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_13 XI11_7/XI0/XI0_52/d__13_ xsel_52_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_12 XI11_7/XI0/XI0_52/d__12_ xsel_52_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_11 XI11_7/XI0/XI0_52/d__11_ xsel_52_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_10 XI11_7/XI0/XI0_52/d__10_ xsel_52_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_9 XI11_7/XI0/XI0_52/d__9_ xsel_52_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_8 XI11_7/XI0/XI0_52/d__8_ xsel_52_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_7 XI11_7/XI0/XI0_52/d__7_ xsel_52_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_6 XI11_7/XI0/XI0_52/d__6_ xsel_52_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_5 XI11_7/XI0/XI0_52/d__5_ xsel_52_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_4 XI11_7/XI0/XI0_52/d__4_ xsel_52_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_3 XI11_7/XI0/XI0_52/d__3_ xsel_52_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_2 XI11_7/XI0/XI0_52/d__2_ xsel_52_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_1 XI11_7/XI0/XI0_52/d__1_ xsel_52_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_52/MN1_0 XI11_7/XI0/XI0_52/d__0_ xsel_52_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_15 XI11_7/net21_0_ xsel_51_ XI11_7/XI0/XI0_51/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_14 XI11_7/net21_1_ xsel_51_ XI11_7/XI0/XI0_51/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_13 XI11_7/net21_2_ xsel_51_ XI11_7/XI0/XI0_51/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_12 XI11_7/net21_3_ xsel_51_ XI11_7/XI0/XI0_51/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_11 XI11_7/net21_4_ xsel_51_ XI11_7/XI0/XI0_51/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_10 XI11_7/net21_5_ xsel_51_ XI11_7/XI0/XI0_51/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_9 XI11_7/net21_6_ xsel_51_ XI11_7/XI0/XI0_51/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_8 XI11_7/net21_7_ xsel_51_ XI11_7/XI0/XI0_51/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_7 XI11_7/net21_8_ xsel_51_ XI11_7/XI0/XI0_51/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_6 XI11_7/net21_9_ xsel_51_ XI11_7/XI0/XI0_51/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_5 XI11_7/net21_10_ xsel_51_ XI11_7/XI0/XI0_51/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_4 XI11_7/net21_11_ xsel_51_ XI11_7/XI0/XI0_51/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_3 XI11_7/net21_12_ xsel_51_ XI11_7/XI0/XI0_51/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_2 XI11_7/net21_13_ xsel_51_ XI11_7/XI0/XI0_51/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_1 XI11_7/net21_14_ xsel_51_ XI11_7/XI0/XI0_51/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN0_0 XI11_7/net21_15_ xsel_51_ XI11_7/XI0/XI0_51/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_15 XI11_7/XI0/XI0_51/d__15_ xsel_51_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_14 XI11_7/XI0/XI0_51/d__14_ xsel_51_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_13 XI11_7/XI0/XI0_51/d__13_ xsel_51_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_12 XI11_7/XI0/XI0_51/d__12_ xsel_51_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_11 XI11_7/XI0/XI0_51/d__11_ xsel_51_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_10 XI11_7/XI0/XI0_51/d__10_ xsel_51_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_9 XI11_7/XI0/XI0_51/d__9_ xsel_51_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_8 XI11_7/XI0/XI0_51/d__8_ xsel_51_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_7 XI11_7/XI0/XI0_51/d__7_ xsel_51_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_6 XI11_7/XI0/XI0_51/d__6_ xsel_51_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_5 XI11_7/XI0/XI0_51/d__5_ xsel_51_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_4 XI11_7/XI0/XI0_51/d__4_ xsel_51_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_3 XI11_7/XI0/XI0_51/d__3_ xsel_51_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_2 XI11_7/XI0/XI0_51/d__2_ xsel_51_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_1 XI11_7/XI0/XI0_51/d__1_ xsel_51_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_51/MN1_0 XI11_7/XI0/XI0_51/d__0_ xsel_51_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_15 XI11_7/net21_0_ xsel_50_ XI11_7/XI0/XI0_50/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_14 XI11_7/net21_1_ xsel_50_ XI11_7/XI0/XI0_50/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_13 XI11_7/net21_2_ xsel_50_ XI11_7/XI0/XI0_50/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_12 XI11_7/net21_3_ xsel_50_ XI11_7/XI0/XI0_50/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_11 XI11_7/net21_4_ xsel_50_ XI11_7/XI0/XI0_50/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_10 XI11_7/net21_5_ xsel_50_ XI11_7/XI0/XI0_50/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_9 XI11_7/net21_6_ xsel_50_ XI11_7/XI0/XI0_50/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_8 XI11_7/net21_7_ xsel_50_ XI11_7/XI0/XI0_50/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_7 XI11_7/net21_8_ xsel_50_ XI11_7/XI0/XI0_50/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_6 XI11_7/net21_9_ xsel_50_ XI11_7/XI0/XI0_50/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_5 XI11_7/net21_10_ xsel_50_ XI11_7/XI0/XI0_50/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_4 XI11_7/net21_11_ xsel_50_ XI11_7/XI0/XI0_50/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_3 XI11_7/net21_12_ xsel_50_ XI11_7/XI0/XI0_50/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_2 XI11_7/net21_13_ xsel_50_ XI11_7/XI0/XI0_50/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_1 XI11_7/net21_14_ xsel_50_ XI11_7/XI0/XI0_50/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN0_0 XI11_7/net21_15_ xsel_50_ XI11_7/XI0/XI0_50/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_15 XI11_7/XI0/XI0_50/d__15_ xsel_50_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_14 XI11_7/XI0/XI0_50/d__14_ xsel_50_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_13 XI11_7/XI0/XI0_50/d__13_ xsel_50_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_12 XI11_7/XI0/XI0_50/d__12_ xsel_50_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_11 XI11_7/XI0/XI0_50/d__11_ xsel_50_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_10 XI11_7/XI0/XI0_50/d__10_ xsel_50_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_9 XI11_7/XI0/XI0_50/d__9_ xsel_50_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_8 XI11_7/XI0/XI0_50/d__8_ xsel_50_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_7 XI11_7/XI0/XI0_50/d__7_ xsel_50_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_6 XI11_7/XI0/XI0_50/d__6_ xsel_50_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_5 XI11_7/XI0/XI0_50/d__5_ xsel_50_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_4 XI11_7/XI0/XI0_50/d__4_ xsel_50_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_3 XI11_7/XI0/XI0_50/d__3_ xsel_50_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_2 XI11_7/XI0/XI0_50/d__2_ xsel_50_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_1 XI11_7/XI0/XI0_50/d__1_ xsel_50_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_50/MN1_0 XI11_7/XI0/XI0_50/d__0_ xsel_50_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_15 XI11_7/net21_0_ xsel_49_ XI11_7/XI0/XI0_49/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_14 XI11_7/net21_1_ xsel_49_ XI11_7/XI0/XI0_49/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_13 XI11_7/net21_2_ xsel_49_ XI11_7/XI0/XI0_49/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_12 XI11_7/net21_3_ xsel_49_ XI11_7/XI0/XI0_49/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_11 XI11_7/net21_4_ xsel_49_ XI11_7/XI0/XI0_49/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_10 XI11_7/net21_5_ xsel_49_ XI11_7/XI0/XI0_49/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_9 XI11_7/net21_6_ xsel_49_ XI11_7/XI0/XI0_49/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_8 XI11_7/net21_7_ xsel_49_ XI11_7/XI0/XI0_49/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_7 XI11_7/net21_8_ xsel_49_ XI11_7/XI0/XI0_49/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_6 XI11_7/net21_9_ xsel_49_ XI11_7/XI0/XI0_49/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_5 XI11_7/net21_10_ xsel_49_ XI11_7/XI0/XI0_49/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_4 XI11_7/net21_11_ xsel_49_ XI11_7/XI0/XI0_49/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_3 XI11_7/net21_12_ xsel_49_ XI11_7/XI0/XI0_49/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_2 XI11_7/net21_13_ xsel_49_ XI11_7/XI0/XI0_49/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_1 XI11_7/net21_14_ xsel_49_ XI11_7/XI0/XI0_49/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN0_0 XI11_7/net21_15_ xsel_49_ XI11_7/XI0/XI0_49/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_15 XI11_7/XI0/XI0_49/d__15_ xsel_49_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_14 XI11_7/XI0/XI0_49/d__14_ xsel_49_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_13 XI11_7/XI0/XI0_49/d__13_ xsel_49_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_12 XI11_7/XI0/XI0_49/d__12_ xsel_49_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_11 XI11_7/XI0/XI0_49/d__11_ xsel_49_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_10 XI11_7/XI0/XI0_49/d__10_ xsel_49_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_9 XI11_7/XI0/XI0_49/d__9_ xsel_49_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_8 XI11_7/XI0/XI0_49/d__8_ xsel_49_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_7 XI11_7/XI0/XI0_49/d__7_ xsel_49_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_6 XI11_7/XI0/XI0_49/d__6_ xsel_49_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_5 XI11_7/XI0/XI0_49/d__5_ xsel_49_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_4 XI11_7/XI0/XI0_49/d__4_ xsel_49_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_3 XI11_7/XI0/XI0_49/d__3_ xsel_49_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_2 XI11_7/XI0/XI0_49/d__2_ xsel_49_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_1 XI11_7/XI0/XI0_49/d__1_ xsel_49_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_49/MN1_0 XI11_7/XI0/XI0_49/d__0_ xsel_49_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_15 XI11_7/net21_0_ xsel_48_ XI11_7/XI0/XI0_48/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_14 XI11_7/net21_1_ xsel_48_ XI11_7/XI0/XI0_48/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_13 XI11_7/net21_2_ xsel_48_ XI11_7/XI0/XI0_48/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_12 XI11_7/net21_3_ xsel_48_ XI11_7/XI0/XI0_48/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_11 XI11_7/net21_4_ xsel_48_ XI11_7/XI0/XI0_48/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_10 XI11_7/net21_5_ xsel_48_ XI11_7/XI0/XI0_48/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_9 XI11_7/net21_6_ xsel_48_ XI11_7/XI0/XI0_48/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_8 XI11_7/net21_7_ xsel_48_ XI11_7/XI0/XI0_48/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_7 XI11_7/net21_8_ xsel_48_ XI11_7/XI0/XI0_48/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_6 XI11_7/net21_9_ xsel_48_ XI11_7/XI0/XI0_48/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_5 XI11_7/net21_10_ xsel_48_ XI11_7/XI0/XI0_48/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_4 XI11_7/net21_11_ xsel_48_ XI11_7/XI0/XI0_48/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_3 XI11_7/net21_12_ xsel_48_ XI11_7/XI0/XI0_48/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_2 XI11_7/net21_13_ xsel_48_ XI11_7/XI0/XI0_48/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_1 XI11_7/net21_14_ xsel_48_ XI11_7/XI0/XI0_48/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN0_0 XI11_7/net21_15_ xsel_48_ XI11_7/XI0/XI0_48/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_15 XI11_7/XI0/XI0_48/d__15_ xsel_48_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_14 XI11_7/XI0/XI0_48/d__14_ xsel_48_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_13 XI11_7/XI0/XI0_48/d__13_ xsel_48_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_12 XI11_7/XI0/XI0_48/d__12_ xsel_48_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_11 XI11_7/XI0/XI0_48/d__11_ xsel_48_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_10 XI11_7/XI0/XI0_48/d__10_ xsel_48_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_9 XI11_7/XI0/XI0_48/d__9_ xsel_48_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_8 XI11_7/XI0/XI0_48/d__8_ xsel_48_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_7 XI11_7/XI0/XI0_48/d__7_ xsel_48_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_6 XI11_7/XI0/XI0_48/d__6_ xsel_48_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_5 XI11_7/XI0/XI0_48/d__5_ xsel_48_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_4 XI11_7/XI0/XI0_48/d__4_ xsel_48_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_3 XI11_7/XI0/XI0_48/d__3_ xsel_48_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_2 XI11_7/XI0/XI0_48/d__2_ xsel_48_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_1 XI11_7/XI0/XI0_48/d__1_ xsel_48_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_48/MN1_0 XI11_7/XI0/XI0_48/d__0_ xsel_48_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_15 XI11_7/net21_0_ xsel_47_ XI11_7/XI0/XI0_47/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_14 XI11_7/net21_1_ xsel_47_ XI11_7/XI0/XI0_47/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_13 XI11_7/net21_2_ xsel_47_ XI11_7/XI0/XI0_47/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_12 XI11_7/net21_3_ xsel_47_ XI11_7/XI0/XI0_47/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_11 XI11_7/net21_4_ xsel_47_ XI11_7/XI0/XI0_47/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_10 XI11_7/net21_5_ xsel_47_ XI11_7/XI0/XI0_47/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_9 XI11_7/net21_6_ xsel_47_ XI11_7/XI0/XI0_47/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_8 XI11_7/net21_7_ xsel_47_ XI11_7/XI0/XI0_47/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_7 XI11_7/net21_8_ xsel_47_ XI11_7/XI0/XI0_47/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_6 XI11_7/net21_9_ xsel_47_ XI11_7/XI0/XI0_47/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_5 XI11_7/net21_10_ xsel_47_ XI11_7/XI0/XI0_47/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_4 XI11_7/net21_11_ xsel_47_ XI11_7/XI0/XI0_47/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_3 XI11_7/net21_12_ xsel_47_ XI11_7/XI0/XI0_47/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_2 XI11_7/net21_13_ xsel_47_ XI11_7/XI0/XI0_47/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_1 XI11_7/net21_14_ xsel_47_ XI11_7/XI0/XI0_47/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN0_0 XI11_7/net21_15_ xsel_47_ XI11_7/XI0/XI0_47/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_15 XI11_7/XI0/XI0_47/d__15_ xsel_47_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_14 XI11_7/XI0/XI0_47/d__14_ xsel_47_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_13 XI11_7/XI0/XI0_47/d__13_ xsel_47_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_12 XI11_7/XI0/XI0_47/d__12_ xsel_47_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_11 XI11_7/XI0/XI0_47/d__11_ xsel_47_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_10 XI11_7/XI0/XI0_47/d__10_ xsel_47_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_9 XI11_7/XI0/XI0_47/d__9_ xsel_47_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_8 XI11_7/XI0/XI0_47/d__8_ xsel_47_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_7 XI11_7/XI0/XI0_47/d__7_ xsel_47_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_6 XI11_7/XI0/XI0_47/d__6_ xsel_47_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_5 XI11_7/XI0/XI0_47/d__5_ xsel_47_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_4 XI11_7/XI0/XI0_47/d__4_ xsel_47_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_3 XI11_7/XI0/XI0_47/d__3_ xsel_47_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_2 XI11_7/XI0/XI0_47/d__2_ xsel_47_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_1 XI11_7/XI0/XI0_47/d__1_ xsel_47_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_47/MN1_0 XI11_7/XI0/XI0_47/d__0_ xsel_47_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_15 XI11_7/net21_0_ xsel_46_ XI11_7/XI0/XI0_46/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_14 XI11_7/net21_1_ xsel_46_ XI11_7/XI0/XI0_46/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_13 XI11_7/net21_2_ xsel_46_ XI11_7/XI0/XI0_46/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_12 XI11_7/net21_3_ xsel_46_ XI11_7/XI0/XI0_46/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_11 XI11_7/net21_4_ xsel_46_ XI11_7/XI0/XI0_46/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_10 XI11_7/net21_5_ xsel_46_ XI11_7/XI0/XI0_46/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_9 XI11_7/net21_6_ xsel_46_ XI11_7/XI0/XI0_46/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_8 XI11_7/net21_7_ xsel_46_ XI11_7/XI0/XI0_46/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_7 XI11_7/net21_8_ xsel_46_ XI11_7/XI0/XI0_46/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_6 XI11_7/net21_9_ xsel_46_ XI11_7/XI0/XI0_46/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_5 XI11_7/net21_10_ xsel_46_ XI11_7/XI0/XI0_46/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_4 XI11_7/net21_11_ xsel_46_ XI11_7/XI0/XI0_46/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_3 XI11_7/net21_12_ xsel_46_ XI11_7/XI0/XI0_46/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_2 XI11_7/net21_13_ xsel_46_ XI11_7/XI0/XI0_46/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_1 XI11_7/net21_14_ xsel_46_ XI11_7/XI0/XI0_46/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN0_0 XI11_7/net21_15_ xsel_46_ XI11_7/XI0/XI0_46/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_15 XI11_7/XI0/XI0_46/d__15_ xsel_46_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_14 XI11_7/XI0/XI0_46/d__14_ xsel_46_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_13 XI11_7/XI0/XI0_46/d__13_ xsel_46_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_12 XI11_7/XI0/XI0_46/d__12_ xsel_46_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_11 XI11_7/XI0/XI0_46/d__11_ xsel_46_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_10 XI11_7/XI0/XI0_46/d__10_ xsel_46_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_9 XI11_7/XI0/XI0_46/d__9_ xsel_46_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_8 XI11_7/XI0/XI0_46/d__8_ xsel_46_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_7 XI11_7/XI0/XI0_46/d__7_ xsel_46_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_6 XI11_7/XI0/XI0_46/d__6_ xsel_46_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_5 XI11_7/XI0/XI0_46/d__5_ xsel_46_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_4 XI11_7/XI0/XI0_46/d__4_ xsel_46_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_3 XI11_7/XI0/XI0_46/d__3_ xsel_46_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_2 XI11_7/XI0/XI0_46/d__2_ xsel_46_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_1 XI11_7/XI0/XI0_46/d__1_ xsel_46_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_46/MN1_0 XI11_7/XI0/XI0_46/d__0_ xsel_46_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_15 XI11_7/net21_0_ xsel_45_ XI11_7/XI0/XI0_45/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_14 XI11_7/net21_1_ xsel_45_ XI11_7/XI0/XI0_45/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_13 XI11_7/net21_2_ xsel_45_ XI11_7/XI0/XI0_45/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_12 XI11_7/net21_3_ xsel_45_ XI11_7/XI0/XI0_45/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_11 XI11_7/net21_4_ xsel_45_ XI11_7/XI0/XI0_45/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_10 XI11_7/net21_5_ xsel_45_ XI11_7/XI0/XI0_45/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_9 XI11_7/net21_6_ xsel_45_ XI11_7/XI0/XI0_45/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_8 XI11_7/net21_7_ xsel_45_ XI11_7/XI0/XI0_45/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_7 XI11_7/net21_8_ xsel_45_ XI11_7/XI0/XI0_45/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_6 XI11_7/net21_9_ xsel_45_ XI11_7/XI0/XI0_45/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_5 XI11_7/net21_10_ xsel_45_ XI11_7/XI0/XI0_45/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_4 XI11_7/net21_11_ xsel_45_ XI11_7/XI0/XI0_45/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_3 XI11_7/net21_12_ xsel_45_ XI11_7/XI0/XI0_45/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_2 XI11_7/net21_13_ xsel_45_ XI11_7/XI0/XI0_45/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_1 XI11_7/net21_14_ xsel_45_ XI11_7/XI0/XI0_45/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN0_0 XI11_7/net21_15_ xsel_45_ XI11_7/XI0/XI0_45/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_15 XI11_7/XI0/XI0_45/d__15_ xsel_45_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_14 XI11_7/XI0/XI0_45/d__14_ xsel_45_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_13 XI11_7/XI0/XI0_45/d__13_ xsel_45_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_12 XI11_7/XI0/XI0_45/d__12_ xsel_45_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_11 XI11_7/XI0/XI0_45/d__11_ xsel_45_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_10 XI11_7/XI0/XI0_45/d__10_ xsel_45_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_9 XI11_7/XI0/XI0_45/d__9_ xsel_45_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_8 XI11_7/XI0/XI0_45/d__8_ xsel_45_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_7 XI11_7/XI0/XI0_45/d__7_ xsel_45_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_6 XI11_7/XI0/XI0_45/d__6_ xsel_45_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_5 XI11_7/XI0/XI0_45/d__5_ xsel_45_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_4 XI11_7/XI0/XI0_45/d__4_ xsel_45_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_3 XI11_7/XI0/XI0_45/d__3_ xsel_45_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_2 XI11_7/XI0/XI0_45/d__2_ xsel_45_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_1 XI11_7/XI0/XI0_45/d__1_ xsel_45_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_45/MN1_0 XI11_7/XI0/XI0_45/d__0_ xsel_45_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_15 XI11_7/net21_0_ xsel_44_ XI11_7/XI0/XI0_44/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_14 XI11_7/net21_1_ xsel_44_ XI11_7/XI0/XI0_44/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_13 XI11_7/net21_2_ xsel_44_ XI11_7/XI0/XI0_44/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_12 XI11_7/net21_3_ xsel_44_ XI11_7/XI0/XI0_44/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_11 XI11_7/net21_4_ xsel_44_ XI11_7/XI0/XI0_44/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_10 XI11_7/net21_5_ xsel_44_ XI11_7/XI0/XI0_44/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_9 XI11_7/net21_6_ xsel_44_ XI11_7/XI0/XI0_44/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_8 XI11_7/net21_7_ xsel_44_ XI11_7/XI0/XI0_44/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_7 XI11_7/net21_8_ xsel_44_ XI11_7/XI0/XI0_44/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_6 XI11_7/net21_9_ xsel_44_ XI11_7/XI0/XI0_44/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_5 XI11_7/net21_10_ xsel_44_ XI11_7/XI0/XI0_44/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_4 XI11_7/net21_11_ xsel_44_ XI11_7/XI0/XI0_44/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_3 XI11_7/net21_12_ xsel_44_ XI11_7/XI0/XI0_44/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_2 XI11_7/net21_13_ xsel_44_ XI11_7/XI0/XI0_44/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_1 XI11_7/net21_14_ xsel_44_ XI11_7/XI0/XI0_44/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN0_0 XI11_7/net21_15_ xsel_44_ XI11_7/XI0/XI0_44/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_15 XI11_7/XI0/XI0_44/d__15_ xsel_44_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_14 XI11_7/XI0/XI0_44/d__14_ xsel_44_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_13 XI11_7/XI0/XI0_44/d__13_ xsel_44_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_12 XI11_7/XI0/XI0_44/d__12_ xsel_44_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_11 XI11_7/XI0/XI0_44/d__11_ xsel_44_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_10 XI11_7/XI0/XI0_44/d__10_ xsel_44_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_9 XI11_7/XI0/XI0_44/d__9_ xsel_44_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_8 XI11_7/XI0/XI0_44/d__8_ xsel_44_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_7 XI11_7/XI0/XI0_44/d__7_ xsel_44_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_6 XI11_7/XI0/XI0_44/d__6_ xsel_44_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_5 XI11_7/XI0/XI0_44/d__5_ xsel_44_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_4 XI11_7/XI0/XI0_44/d__4_ xsel_44_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_3 XI11_7/XI0/XI0_44/d__3_ xsel_44_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_2 XI11_7/XI0/XI0_44/d__2_ xsel_44_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_1 XI11_7/XI0/XI0_44/d__1_ xsel_44_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_44/MN1_0 XI11_7/XI0/XI0_44/d__0_ xsel_44_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_15 XI11_7/net21_0_ xsel_43_ XI11_7/XI0/XI0_43/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_14 XI11_7/net21_1_ xsel_43_ XI11_7/XI0/XI0_43/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_13 XI11_7/net21_2_ xsel_43_ XI11_7/XI0/XI0_43/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_12 XI11_7/net21_3_ xsel_43_ XI11_7/XI0/XI0_43/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_11 XI11_7/net21_4_ xsel_43_ XI11_7/XI0/XI0_43/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_10 XI11_7/net21_5_ xsel_43_ XI11_7/XI0/XI0_43/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_9 XI11_7/net21_6_ xsel_43_ XI11_7/XI0/XI0_43/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_8 XI11_7/net21_7_ xsel_43_ XI11_7/XI0/XI0_43/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_7 XI11_7/net21_8_ xsel_43_ XI11_7/XI0/XI0_43/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_6 XI11_7/net21_9_ xsel_43_ XI11_7/XI0/XI0_43/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_5 XI11_7/net21_10_ xsel_43_ XI11_7/XI0/XI0_43/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_4 XI11_7/net21_11_ xsel_43_ XI11_7/XI0/XI0_43/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_3 XI11_7/net21_12_ xsel_43_ XI11_7/XI0/XI0_43/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_2 XI11_7/net21_13_ xsel_43_ XI11_7/XI0/XI0_43/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_1 XI11_7/net21_14_ xsel_43_ XI11_7/XI0/XI0_43/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN0_0 XI11_7/net21_15_ xsel_43_ XI11_7/XI0/XI0_43/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_15 XI11_7/XI0/XI0_43/d__15_ xsel_43_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_14 XI11_7/XI0/XI0_43/d__14_ xsel_43_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_13 XI11_7/XI0/XI0_43/d__13_ xsel_43_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_12 XI11_7/XI0/XI0_43/d__12_ xsel_43_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_11 XI11_7/XI0/XI0_43/d__11_ xsel_43_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_10 XI11_7/XI0/XI0_43/d__10_ xsel_43_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_9 XI11_7/XI0/XI0_43/d__9_ xsel_43_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_8 XI11_7/XI0/XI0_43/d__8_ xsel_43_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_7 XI11_7/XI0/XI0_43/d__7_ xsel_43_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_6 XI11_7/XI0/XI0_43/d__6_ xsel_43_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_5 XI11_7/XI0/XI0_43/d__5_ xsel_43_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_4 XI11_7/XI0/XI0_43/d__4_ xsel_43_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_3 XI11_7/XI0/XI0_43/d__3_ xsel_43_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_2 XI11_7/XI0/XI0_43/d__2_ xsel_43_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_1 XI11_7/XI0/XI0_43/d__1_ xsel_43_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_43/MN1_0 XI11_7/XI0/XI0_43/d__0_ xsel_43_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_15 XI11_7/net21_0_ xsel_42_ XI11_7/XI0/XI0_42/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_14 XI11_7/net21_1_ xsel_42_ XI11_7/XI0/XI0_42/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_13 XI11_7/net21_2_ xsel_42_ XI11_7/XI0/XI0_42/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_12 XI11_7/net21_3_ xsel_42_ XI11_7/XI0/XI0_42/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_11 XI11_7/net21_4_ xsel_42_ XI11_7/XI0/XI0_42/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_10 XI11_7/net21_5_ xsel_42_ XI11_7/XI0/XI0_42/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_9 XI11_7/net21_6_ xsel_42_ XI11_7/XI0/XI0_42/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_8 XI11_7/net21_7_ xsel_42_ XI11_7/XI0/XI0_42/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_7 XI11_7/net21_8_ xsel_42_ XI11_7/XI0/XI0_42/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_6 XI11_7/net21_9_ xsel_42_ XI11_7/XI0/XI0_42/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_5 XI11_7/net21_10_ xsel_42_ XI11_7/XI0/XI0_42/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_4 XI11_7/net21_11_ xsel_42_ XI11_7/XI0/XI0_42/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_3 XI11_7/net21_12_ xsel_42_ XI11_7/XI0/XI0_42/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_2 XI11_7/net21_13_ xsel_42_ XI11_7/XI0/XI0_42/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_1 XI11_7/net21_14_ xsel_42_ XI11_7/XI0/XI0_42/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN0_0 XI11_7/net21_15_ xsel_42_ XI11_7/XI0/XI0_42/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_15 XI11_7/XI0/XI0_42/d__15_ xsel_42_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_14 XI11_7/XI0/XI0_42/d__14_ xsel_42_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_13 XI11_7/XI0/XI0_42/d__13_ xsel_42_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_12 XI11_7/XI0/XI0_42/d__12_ xsel_42_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_11 XI11_7/XI0/XI0_42/d__11_ xsel_42_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_10 XI11_7/XI0/XI0_42/d__10_ xsel_42_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_9 XI11_7/XI0/XI0_42/d__9_ xsel_42_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_8 XI11_7/XI0/XI0_42/d__8_ xsel_42_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_7 XI11_7/XI0/XI0_42/d__7_ xsel_42_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_6 XI11_7/XI0/XI0_42/d__6_ xsel_42_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_5 XI11_7/XI0/XI0_42/d__5_ xsel_42_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_4 XI11_7/XI0/XI0_42/d__4_ xsel_42_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_3 XI11_7/XI0/XI0_42/d__3_ xsel_42_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_2 XI11_7/XI0/XI0_42/d__2_ xsel_42_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_1 XI11_7/XI0/XI0_42/d__1_ xsel_42_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_42/MN1_0 XI11_7/XI0/XI0_42/d__0_ xsel_42_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_15 XI11_7/net21_0_ xsel_41_ XI11_7/XI0/XI0_41/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_14 XI11_7/net21_1_ xsel_41_ XI11_7/XI0/XI0_41/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_13 XI11_7/net21_2_ xsel_41_ XI11_7/XI0/XI0_41/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_12 XI11_7/net21_3_ xsel_41_ XI11_7/XI0/XI0_41/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_11 XI11_7/net21_4_ xsel_41_ XI11_7/XI0/XI0_41/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_10 XI11_7/net21_5_ xsel_41_ XI11_7/XI0/XI0_41/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_9 XI11_7/net21_6_ xsel_41_ XI11_7/XI0/XI0_41/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_8 XI11_7/net21_7_ xsel_41_ XI11_7/XI0/XI0_41/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_7 XI11_7/net21_8_ xsel_41_ XI11_7/XI0/XI0_41/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_6 XI11_7/net21_9_ xsel_41_ XI11_7/XI0/XI0_41/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_5 XI11_7/net21_10_ xsel_41_ XI11_7/XI0/XI0_41/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_4 XI11_7/net21_11_ xsel_41_ XI11_7/XI0/XI0_41/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_3 XI11_7/net21_12_ xsel_41_ XI11_7/XI0/XI0_41/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_2 XI11_7/net21_13_ xsel_41_ XI11_7/XI0/XI0_41/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_1 XI11_7/net21_14_ xsel_41_ XI11_7/XI0/XI0_41/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN0_0 XI11_7/net21_15_ xsel_41_ XI11_7/XI0/XI0_41/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_15 XI11_7/XI0/XI0_41/d__15_ xsel_41_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_14 XI11_7/XI0/XI0_41/d__14_ xsel_41_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_13 XI11_7/XI0/XI0_41/d__13_ xsel_41_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_12 XI11_7/XI0/XI0_41/d__12_ xsel_41_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_11 XI11_7/XI0/XI0_41/d__11_ xsel_41_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_10 XI11_7/XI0/XI0_41/d__10_ xsel_41_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_9 XI11_7/XI0/XI0_41/d__9_ xsel_41_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_8 XI11_7/XI0/XI0_41/d__8_ xsel_41_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_7 XI11_7/XI0/XI0_41/d__7_ xsel_41_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_6 XI11_7/XI0/XI0_41/d__6_ xsel_41_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_5 XI11_7/XI0/XI0_41/d__5_ xsel_41_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_4 XI11_7/XI0/XI0_41/d__4_ xsel_41_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_3 XI11_7/XI0/XI0_41/d__3_ xsel_41_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_2 XI11_7/XI0/XI0_41/d__2_ xsel_41_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_1 XI11_7/XI0/XI0_41/d__1_ xsel_41_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_41/MN1_0 XI11_7/XI0/XI0_41/d__0_ xsel_41_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_15 XI11_7/net21_0_ xsel_40_ XI11_7/XI0/XI0_40/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_14 XI11_7/net21_1_ xsel_40_ XI11_7/XI0/XI0_40/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_13 XI11_7/net21_2_ xsel_40_ XI11_7/XI0/XI0_40/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_12 XI11_7/net21_3_ xsel_40_ XI11_7/XI0/XI0_40/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_11 XI11_7/net21_4_ xsel_40_ XI11_7/XI0/XI0_40/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_10 XI11_7/net21_5_ xsel_40_ XI11_7/XI0/XI0_40/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_9 XI11_7/net21_6_ xsel_40_ XI11_7/XI0/XI0_40/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_8 XI11_7/net21_7_ xsel_40_ XI11_7/XI0/XI0_40/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_7 XI11_7/net21_8_ xsel_40_ XI11_7/XI0/XI0_40/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_6 XI11_7/net21_9_ xsel_40_ XI11_7/XI0/XI0_40/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_5 XI11_7/net21_10_ xsel_40_ XI11_7/XI0/XI0_40/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_4 XI11_7/net21_11_ xsel_40_ XI11_7/XI0/XI0_40/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_3 XI11_7/net21_12_ xsel_40_ XI11_7/XI0/XI0_40/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_2 XI11_7/net21_13_ xsel_40_ XI11_7/XI0/XI0_40/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_1 XI11_7/net21_14_ xsel_40_ XI11_7/XI0/XI0_40/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN0_0 XI11_7/net21_15_ xsel_40_ XI11_7/XI0/XI0_40/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_15 XI11_7/XI0/XI0_40/d__15_ xsel_40_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_14 XI11_7/XI0/XI0_40/d__14_ xsel_40_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_13 XI11_7/XI0/XI0_40/d__13_ xsel_40_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_12 XI11_7/XI0/XI0_40/d__12_ xsel_40_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_11 XI11_7/XI0/XI0_40/d__11_ xsel_40_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_10 XI11_7/XI0/XI0_40/d__10_ xsel_40_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_9 XI11_7/XI0/XI0_40/d__9_ xsel_40_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_8 XI11_7/XI0/XI0_40/d__8_ xsel_40_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_7 XI11_7/XI0/XI0_40/d__7_ xsel_40_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_6 XI11_7/XI0/XI0_40/d__6_ xsel_40_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_5 XI11_7/XI0/XI0_40/d__5_ xsel_40_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_4 XI11_7/XI0/XI0_40/d__4_ xsel_40_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_3 XI11_7/XI0/XI0_40/d__3_ xsel_40_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_2 XI11_7/XI0/XI0_40/d__2_ xsel_40_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_1 XI11_7/XI0/XI0_40/d__1_ xsel_40_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_40/MN1_0 XI11_7/XI0/XI0_40/d__0_ xsel_40_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_15 XI11_7/net21_0_ xsel_39_ XI11_7/XI0/XI0_39/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_14 XI11_7/net21_1_ xsel_39_ XI11_7/XI0/XI0_39/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_13 XI11_7/net21_2_ xsel_39_ XI11_7/XI0/XI0_39/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_12 XI11_7/net21_3_ xsel_39_ XI11_7/XI0/XI0_39/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_11 XI11_7/net21_4_ xsel_39_ XI11_7/XI0/XI0_39/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_10 XI11_7/net21_5_ xsel_39_ XI11_7/XI0/XI0_39/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_9 XI11_7/net21_6_ xsel_39_ XI11_7/XI0/XI0_39/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_8 XI11_7/net21_7_ xsel_39_ XI11_7/XI0/XI0_39/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_7 XI11_7/net21_8_ xsel_39_ XI11_7/XI0/XI0_39/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_6 XI11_7/net21_9_ xsel_39_ XI11_7/XI0/XI0_39/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_5 XI11_7/net21_10_ xsel_39_ XI11_7/XI0/XI0_39/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_4 XI11_7/net21_11_ xsel_39_ XI11_7/XI0/XI0_39/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_3 XI11_7/net21_12_ xsel_39_ XI11_7/XI0/XI0_39/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_2 XI11_7/net21_13_ xsel_39_ XI11_7/XI0/XI0_39/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_1 XI11_7/net21_14_ xsel_39_ XI11_7/XI0/XI0_39/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN0_0 XI11_7/net21_15_ xsel_39_ XI11_7/XI0/XI0_39/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_15 XI11_7/XI0/XI0_39/d__15_ xsel_39_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_14 XI11_7/XI0/XI0_39/d__14_ xsel_39_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_13 XI11_7/XI0/XI0_39/d__13_ xsel_39_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_12 XI11_7/XI0/XI0_39/d__12_ xsel_39_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_11 XI11_7/XI0/XI0_39/d__11_ xsel_39_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_10 XI11_7/XI0/XI0_39/d__10_ xsel_39_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_9 XI11_7/XI0/XI0_39/d__9_ xsel_39_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_8 XI11_7/XI0/XI0_39/d__8_ xsel_39_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_7 XI11_7/XI0/XI0_39/d__7_ xsel_39_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_6 XI11_7/XI0/XI0_39/d__6_ xsel_39_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_5 XI11_7/XI0/XI0_39/d__5_ xsel_39_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_4 XI11_7/XI0/XI0_39/d__4_ xsel_39_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_3 XI11_7/XI0/XI0_39/d__3_ xsel_39_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_2 XI11_7/XI0/XI0_39/d__2_ xsel_39_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_1 XI11_7/XI0/XI0_39/d__1_ xsel_39_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_39/MN1_0 XI11_7/XI0/XI0_39/d__0_ xsel_39_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_15 XI11_7/net21_0_ xsel_38_ XI11_7/XI0/XI0_38/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_14 XI11_7/net21_1_ xsel_38_ XI11_7/XI0/XI0_38/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_13 XI11_7/net21_2_ xsel_38_ XI11_7/XI0/XI0_38/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_12 XI11_7/net21_3_ xsel_38_ XI11_7/XI0/XI0_38/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_11 XI11_7/net21_4_ xsel_38_ XI11_7/XI0/XI0_38/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_10 XI11_7/net21_5_ xsel_38_ XI11_7/XI0/XI0_38/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_9 XI11_7/net21_6_ xsel_38_ XI11_7/XI0/XI0_38/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_8 XI11_7/net21_7_ xsel_38_ XI11_7/XI0/XI0_38/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_7 XI11_7/net21_8_ xsel_38_ XI11_7/XI0/XI0_38/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_6 XI11_7/net21_9_ xsel_38_ XI11_7/XI0/XI0_38/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_5 XI11_7/net21_10_ xsel_38_ XI11_7/XI0/XI0_38/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_4 XI11_7/net21_11_ xsel_38_ XI11_7/XI0/XI0_38/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_3 XI11_7/net21_12_ xsel_38_ XI11_7/XI0/XI0_38/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_2 XI11_7/net21_13_ xsel_38_ XI11_7/XI0/XI0_38/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_1 XI11_7/net21_14_ xsel_38_ XI11_7/XI0/XI0_38/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN0_0 XI11_7/net21_15_ xsel_38_ XI11_7/XI0/XI0_38/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_15 XI11_7/XI0/XI0_38/d__15_ xsel_38_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_14 XI11_7/XI0/XI0_38/d__14_ xsel_38_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_13 XI11_7/XI0/XI0_38/d__13_ xsel_38_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_12 XI11_7/XI0/XI0_38/d__12_ xsel_38_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_11 XI11_7/XI0/XI0_38/d__11_ xsel_38_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_10 XI11_7/XI0/XI0_38/d__10_ xsel_38_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_9 XI11_7/XI0/XI0_38/d__9_ xsel_38_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_8 XI11_7/XI0/XI0_38/d__8_ xsel_38_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_7 XI11_7/XI0/XI0_38/d__7_ xsel_38_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_6 XI11_7/XI0/XI0_38/d__6_ xsel_38_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_5 XI11_7/XI0/XI0_38/d__5_ xsel_38_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_4 XI11_7/XI0/XI0_38/d__4_ xsel_38_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_3 XI11_7/XI0/XI0_38/d__3_ xsel_38_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_2 XI11_7/XI0/XI0_38/d__2_ xsel_38_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_1 XI11_7/XI0/XI0_38/d__1_ xsel_38_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_38/MN1_0 XI11_7/XI0/XI0_38/d__0_ xsel_38_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_15 XI11_7/net21_0_ xsel_37_ XI11_7/XI0/XI0_37/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_14 XI11_7/net21_1_ xsel_37_ XI11_7/XI0/XI0_37/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_13 XI11_7/net21_2_ xsel_37_ XI11_7/XI0/XI0_37/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_12 XI11_7/net21_3_ xsel_37_ XI11_7/XI0/XI0_37/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_11 XI11_7/net21_4_ xsel_37_ XI11_7/XI0/XI0_37/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_10 XI11_7/net21_5_ xsel_37_ XI11_7/XI0/XI0_37/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_9 XI11_7/net21_6_ xsel_37_ XI11_7/XI0/XI0_37/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_8 XI11_7/net21_7_ xsel_37_ XI11_7/XI0/XI0_37/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_7 XI11_7/net21_8_ xsel_37_ XI11_7/XI0/XI0_37/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_6 XI11_7/net21_9_ xsel_37_ XI11_7/XI0/XI0_37/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_5 XI11_7/net21_10_ xsel_37_ XI11_7/XI0/XI0_37/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_4 XI11_7/net21_11_ xsel_37_ XI11_7/XI0/XI0_37/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_3 XI11_7/net21_12_ xsel_37_ XI11_7/XI0/XI0_37/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_2 XI11_7/net21_13_ xsel_37_ XI11_7/XI0/XI0_37/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_1 XI11_7/net21_14_ xsel_37_ XI11_7/XI0/XI0_37/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN0_0 XI11_7/net21_15_ xsel_37_ XI11_7/XI0/XI0_37/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_15 XI11_7/XI0/XI0_37/d__15_ xsel_37_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_14 XI11_7/XI0/XI0_37/d__14_ xsel_37_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_13 XI11_7/XI0/XI0_37/d__13_ xsel_37_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_12 XI11_7/XI0/XI0_37/d__12_ xsel_37_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_11 XI11_7/XI0/XI0_37/d__11_ xsel_37_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_10 XI11_7/XI0/XI0_37/d__10_ xsel_37_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_9 XI11_7/XI0/XI0_37/d__9_ xsel_37_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_8 XI11_7/XI0/XI0_37/d__8_ xsel_37_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_7 XI11_7/XI0/XI0_37/d__7_ xsel_37_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_6 XI11_7/XI0/XI0_37/d__6_ xsel_37_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_5 XI11_7/XI0/XI0_37/d__5_ xsel_37_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_4 XI11_7/XI0/XI0_37/d__4_ xsel_37_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_3 XI11_7/XI0/XI0_37/d__3_ xsel_37_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_2 XI11_7/XI0/XI0_37/d__2_ xsel_37_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_1 XI11_7/XI0/XI0_37/d__1_ xsel_37_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_37/MN1_0 XI11_7/XI0/XI0_37/d__0_ xsel_37_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_15 XI11_7/net21_0_ xsel_36_ XI11_7/XI0/XI0_36/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_14 XI11_7/net21_1_ xsel_36_ XI11_7/XI0/XI0_36/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_13 XI11_7/net21_2_ xsel_36_ XI11_7/XI0/XI0_36/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_12 XI11_7/net21_3_ xsel_36_ XI11_7/XI0/XI0_36/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_11 XI11_7/net21_4_ xsel_36_ XI11_7/XI0/XI0_36/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_10 XI11_7/net21_5_ xsel_36_ XI11_7/XI0/XI0_36/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_9 XI11_7/net21_6_ xsel_36_ XI11_7/XI0/XI0_36/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_8 XI11_7/net21_7_ xsel_36_ XI11_7/XI0/XI0_36/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_7 XI11_7/net21_8_ xsel_36_ XI11_7/XI0/XI0_36/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_6 XI11_7/net21_9_ xsel_36_ XI11_7/XI0/XI0_36/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_5 XI11_7/net21_10_ xsel_36_ XI11_7/XI0/XI0_36/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_4 XI11_7/net21_11_ xsel_36_ XI11_7/XI0/XI0_36/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_3 XI11_7/net21_12_ xsel_36_ XI11_7/XI0/XI0_36/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_2 XI11_7/net21_13_ xsel_36_ XI11_7/XI0/XI0_36/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_1 XI11_7/net21_14_ xsel_36_ XI11_7/XI0/XI0_36/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN0_0 XI11_7/net21_15_ xsel_36_ XI11_7/XI0/XI0_36/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_15 XI11_7/XI0/XI0_36/d__15_ xsel_36_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_14 XI11_7/XI0/XI0_36/d__14_ xsel_36_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_13 XI11_7/XI0/XI0_36/d__13_ xsel_36_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_12 XI11_7/XI0/XI0_36/d__12_ xsel_36_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_11 XI11_7/XI0/XI0_36/d__11_ xsel_36_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_10 XI11_7/XI0/XI0_36/d__10_ xsel_36_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_9 XI11_7/XI0/XI0_36/d__9_ xsel_36_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_8 XI11_7/XI0/XI0_36/d__8_ xsel_36_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_7 XI11_7/XI0/XI0_36/d__7_ xsel_36_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_6 XI11_7/XI0/XI0_36/d__6_ xsel_36_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_5 XI11_7/XI0/XI0_36/d__5_ xsel_36_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_4 XI11_7/XI0/XI0_36/d__4_ xsel_36_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_3 XI11_7/XI0/XI0_36/d__3_ xsel_36_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_2 XI11_7/XI0/XI0_36/d__2_ xsel_36_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_1 XI11_7/XI0/XI0_36/d__1_ xsel_36_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_36/MN1_0 XI11_7/XI0/XI0_36/d__0_ xsel_36_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_15 XI11_7/net21_0_ xsel_35_ XI11_7/XI0/XI0_35/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_14 XI11_7/net21_1_ xsel_35_ XI11_7/XI0/XI0_35/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_13 XI11_7/net21_2_ xsel_35_ XI11_7/XI0/XI0_35/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_12 XI11_7/net21_3_ xsel_35_ XI11_7/XI0/XI0_35/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_11 XI11_7/net21_4_ xsel_35_ XI11_7/XI0/XI0_35/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_10 XI11_7/net21_5_ xsel_35_ XI11_7/XI0/XI0_35/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_9 XI11_7/net21_6_ xsel_35_ XI11_7/XI0/XI0_35/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_8 XI11_7/net21_7_ xsel_35_ XI11_7/XI0/XI0_35/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_7 XI11_7/net21_8_ xsel_35_ XI11_7/XI0/XI0_35/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_6 XI11_7/net21_9_ xsel_35_ XI11_7/XI0/XI0_35/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_5 XI11_7/net21_10_ xsel_35_ XI11_7/XI0/XI0_35/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_4 XI11_7/net21_11_ xsel_35_ XI11_7/XI0/XI0_35/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_3 XI11_7/net21_12_ xsel_35_ XI11_7/XI0/XI0_35/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_2 XI11_7/net21_13_ xsel_35_ XI11_7/XI0/XI0_35/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_1 XI11_7/net21_14_ xsel_35_ XI11_7/XI0/XI0_35/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN0_0 XI11_7/net21_15_ xsel_35_ XI11_7/XI0/XI0_35/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_15 XI11_7/XI0/XI0_35/d__15_ xsel_35_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_14 XI11_7/XI0/XI0_35/d__14_ xsel_35_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_13 XI11_7/XI0/XI0_35/d__13_ xsel_35_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_12 XI11_7/XI0/XI0_35/d__12_ xsel_35_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_11 XI11_7/XI0/XI0_35/d__11_ xsel_35_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_10 XI11_7/XI0/XI0_35/d__10_ xsel_35_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_9 XI11_7/XI0/XI0_35/d__9_ xsel_35_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_8 XI11_7/XI0/XI0_35/d__8_ xsel_35_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_7 XI11_7/XI0/XI0_35/d__7_ xsel_35_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_6 XI11_7/XI0/XI0_35/d__6_ xsel_35_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_5 XI11_7/XI0/XI0_35/d__5_ xsel_35_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_4 XI11_7/XI0/XI0_35/d__4_ xsel_35_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_3 XI11_7/XI0/XI0_35/d__3_ xsel_35_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_2 XI11_7/XI0/XI0_35/d__2_ xsel_35_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_1 XI11_7/XI0/XI0_35/d__1_ xsel_35_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_35/MN1_0 XI11_7/XI0/XI0_35/d__0_ xsel_35_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_15 XI11_7/net21_0_ xsel_34_ XI11_7/XI0/XI0_34/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_14 XI11_7/net21_1_ xsel_34_ XI11_7/XI0/XI0_34/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_13 XI11_7/net21_2_ xsel_34_ XI11_7/XI0/XI0_34/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_12 XI11_7/net21_3_ xsel_34_ XI11_7/XI0/XI0_34/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_11 XI11_7/net21_4_ xsel_34_ XI11_7/XI0/XI0_34/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_10 XI11_7/net21_5_ xsel_34_ XI11_7/XI0/XI0_34/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_9 XI11_7/net21_6_ xsel_34_ XI11_7/XI0/XI0_34/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_8 XI11_7/net21_7_ xsel_34_ XI11_7/XI0/XI0_34/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_7 XI11_7/net21_8_ xsel_34_ XI11_7/XI0/XI0_34/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_6 XI11_7/net21_9_ xsel_34_ XI11_7/XI0/XI0_34/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_5 XI11_7/net21_10_ xsel_34_ XI11_7/XI0/XI0_34/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_4 XI11_7/net21_11_ xsel_34_ XI11_7/XI0/XI0_34/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_3 XI11_7/net21_12_ xsel_34_ XI11_7/XI0/XI0_34/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_2 XI11_7/net21_13_ xsel_34_ XI11_7/XI0/XI0_34/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_1 XI11_7/net21_14_ xsel_34_ XI11_7/XI0/XI0_34/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN0_0 XI11_7/net21_15_ xsel_34_ XI11_7/XI0/XI0_34/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_15 XI11_7/XI0/XI0_34/d__15_ xsel_34_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_14 XI11_7/XI0/XI0_34/d__14_ xsel_34_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_13 XI11_7/XI0/XI0_34/d__13_ xsel_34_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_12 XI11_7/XI0/XI0_34/d__12_ xsel_34_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_11 XI11_7/XI0/XI0_34/d__11_ xsel_34_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_10 XI11_7/XI0/XI0_34/d__10_ xsel_34_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_9 XI11_7/XI0/XI0_34/d__9_ xsel_34_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_8 XI11_7/XI0/XI0_34/d__8_ xsel_34_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_7 XI11_7/XI0/XI0_34/d__7_ xsel_34_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_6 XI11_7/XI0/XI0_34/d__6_ xsel_34_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_5 XI11_7/XI0/XI0_34/d__5_ xsel_34_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_4 XI11_7/XI0/XI0_34/d__4_ xsel_34_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_3 XI11_7/XI0/XI0_34/d__3_ xsel_34_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_2 XI11_7/XI0/XI0_34/d__2_ xsel_34_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_1 XI11_7/XI0/XI0_34/d__1_ xsel_34_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_34/MN1_0 XI11_7/XI0/XI0_34/d__0_ xsel_34_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_15 XI11_7/net21_0_ xsel_33_ XI11_7/XI0/XI0_33/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_14 XI11_7/net21_1_ xsel_33_ XI11_7/XI0/XI0_33/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_13 XI11_7/net21_2_ xsel_33_ XI11_7/XI0/XI0_33/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_12 XI11_7/net21_3_ xsel_33_ XI11_7/XI0/XI0_33/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_11 XI11_7/net21_4_ xsel_33_ XI11_7/XI0/XI0_33/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_10 XI11_7/net21_5_ xsel_33_ XI11_7/XI0/XI0_33/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_9 XI11_7/net21_6_ xsel_33_ XI11_7/XI0/XI0_33/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_8 XI11_7/net21_7_ xsel_33_ XI11_7/XI0/XI0_33/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_7 XI11_7/net21_8_ xsel_33_ XI11_7/XI0/XI0_33/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_6 XI11_7/net21_9_ xsel_33_ XI11_7/XI0/XI0_33/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_5 XI11_7/net21_10_ xsel_33_ XI11_7/XI0/XI0_33/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_4 XI11_7/net21_11_ xsel_33_ XI11_7/XI0/XI0_33/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_3 XI11_7/net21_12_ xsel_33_ XI11_7/XI0/XI0_33/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_2 XI11_7/net21_13_ xsel_33_ XI11_7/XI0/XI0_33/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_1 XI11_7/net21_14_ xsel_33_ XI11_7/XI0/XI0_33/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN0_0 XI11_7/net21_15_ xsel_33_ XI11_7/XI0/XI0_33/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_15 XI11_7/XI0/XI0_33/d__15_ xsel_33_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_14 XI11_7/XI0/XI0_33/d__14_ xsel_33_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_13 XI11_7/XI0/XI0_33/d__13_ xsel_33_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_12 XI11_7/XI0/XI0_33/d__12_ xsel_33_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_11 XI11_7/XI0/XI0_33/d__11_ xsel_33_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_10 XI11_7/XI0/XI0_33/d__10_ xsel_33_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_9 XI11_7/XI0/XI0_33/d__9_ xsel_33_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_8 XI11_7/XI0/XI0_33/d__8_ xsel_33_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_7 XI11_7/XI0/XI0_33/d__7_ xsel_33_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_6 XI11_7/XI0/XI0_33/d__6_ xsel_33_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_5 XI11_7/XI0/XI0_33/d__5_ xsel_33_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_4 XI11_7/XI0/XI0_33/d__4_ xsel_33_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_3 XI11_7/XI0/XI0_33/d__3_ xsel_33_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_2 XI11_7/XI0/XI0_33/d__2_ xsel_33_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_1 XI11_7/XI0/XI0_33/d__1_ xsel_33_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_33/MN1_0 XI11_7/XI0/XI0_33/d__0_ xsel_33_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_15 XI11_7/net21_0_ xsel_32_ XI11_7/XI0/XI0_32/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_14 XI11_7/net21_1_ xsel_32_ XI11_7/XI0/XI0_32/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_13 XI11_7/net21_2_ xsel_32_ XI11_7/XI0/XI0_32/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_12 XI11_7/net21_3_ xsel_32_ XI11_7/XI0/XI0_32/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_11 XI11_7/net21_4_ xsel_32_ XI11_7/XI0/XI0_32/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_10 XI11_7/net21_5_ xsel_32_ XI11_7/XI0/XI0_32/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_9 XI11_7/net21_6_ xsel_32_ XI11_7/XI0/XI0_32/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_8 XI11_7/net21_7_ xsel_32_ XI11_7/XI0/XI0_32/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_7 XI11_7/net21_8_ xsel_32_ XI11_7/XI0/XI0_32/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_6 XI11_7/net21_9_ xsel_32_ XI11_7/XI0/XI0_32/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_5 XI11_7/net21_10_ xsel_32_ XI11_7/XI0/XI0_32/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_4 XI11_7/net21_11_ xsel_32_ XI11_7/XI0/XI0_32/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_3 XI11_7/net21_12_ xsel_32_ XI11_7/XI0/XI0_32/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_2 XI11_7/net21_13_ xsel_32_ XI11_7/XI0/XI0_32/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_1 XI11_7/net21_14_ xsel_32_ XI11_7/XI0/XI0_32/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN0_0 XI11_7/net21_15_ xsel_32_ XI11_7/XI0/XI0_32/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_15 XI11_7/XI0/XI0_32/d__15_ xsel_32_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_14 XI11_7/XI0/XI0_32/d__14_ xsel_32_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_13 XI11_7/XI0/XI0_32/d__13_ xsel_32_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_12 XI11_7/XI0/XI0_32/d__12_ xsel_32_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_11 XI11_7/XI0/XI0_32/d__11_ xsel_32_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_10 XI11_7/XI0/XI0_32/d__10_ xsel_32_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_9 XI11_7/XI0/XI0_32/d__9_ xsel_32_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_8 XI11_7/XI0/XI0_32/d__8_ xsel_32_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_7 XI11_7/XI0/XI0_32/d__7_ xsel_32_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_6 XI11_7/XI0/XI0_32/d__6_ xsel_32_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_5 XI11_7/XI0/XI0_32/d__5_ xsel_32_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_4 XI11_7/XI0/XI0_32/d__4_ xsel_32_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_3 XI11_7/XI0/XI0_32/d__3_ xsel_32_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_2 XI11_7/XI0/XI0_32/d__2_ xsel_32_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_1 XI11_7/XI0/XI0_32/d__1_ xsel_32_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_32/MN1_0 XI11_7/XI0/XI0_32/d__0_ xsel_32_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_15 XI11_7/net21_0_ xsel_31_ XI11_7/XI0/XI0_31/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_14 XI11_7/net21_1_ xsel_31_ XI11_7/XI0/XI0_31/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_13 XI11_7/net21_2_ xsel_31_ XI11_7/XI0/XI0_31/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_12 XI11_7/net21_3_ xsel_31_ XI11_7/XI0/XI0_31/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_11 XI11_7/net21_4_ xsel_31_ XI11_7/XI0/XI0_31/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_10 XI11_7/net21_5_ xsel_31_ XI11_7/XI0/XI0_31/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_9 XI11_7/net21_6_ xsel_31_ XI11_7/XI0/XI0_31/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_8 XI11_7/net21_7_ xsel_31_ XI11_7/XI0/XI0_31/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_7 XI11_7/net21_8_ xsel_31_ XI11_7/XI0/XI0_31/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_6 XI11_7/net21_9_ xsel_31_ XI11_7/XI0/XI0_31/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_5 XI11_7/net21_10_ xsel_31_ XI11_7/XI0/XI0_31/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_4 XI11_7/net21_11_ xsel_31_ XI11_7/XI0/XI0_31/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_3 XI11_7/net21_12_ xsel_31_ XI11_7/XI0/XI0_31/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_2 XI11_7/net21_13_ xsel_31_ XI11_7/XI0/XI0_31/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_1 XI11_7/net21_14_ xsel_31_ XI11_7/XI0/XI0_31/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN0_0 XI11_7/net21_15_ xsel_31_ XI11_7/XI0/XI0_31/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_15 XI11_7/XI0/XI0_31/d__15_ xsel_31_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_14 XI11_7/XI0/XI0_31/d__14_ xsel_31_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_13 XI11_7/XI0/XI0_31/d__13_ xsel_31_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_12 XI11_7/XI0/XI0_31/d__12_ xsel_31_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_11 XI11_7/XI0/XI0_31/d__11_ xsel_31_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_10 XI11_7/XI0/XI0_31/d__10_ xsel_31_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_9 XI11_7/XI0/XI0_31/d__9_ xsel_31_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_8 XI11_7/XI0/XI0_31/d__8_ xsel_31_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_7 XI11_7/XI0/XI0_31/d__7_ xsel_31_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_6 XI11_7/XI0/XI0_31/d__6_ xsel_31_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_5 XI11_7/XI0/XI0_31/d__5_ xsel_31_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_4 XI11_7/XI0/XI0_31/d__4_ xsel_31_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_3 XI11_7/XI0/XI0_31/d__3_ xsel_31_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_2 XI11_7/XI0/XI0_31/d__2_ xsel_31_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_1 XI11_7/XI0/XI0_31/d__1_ xsel_31_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_31/MN1_0 XI11_7/XI0/XI0_31/d__0_ xsel_31_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_15 XI11_7/net21_0_ xsel_30_ XI11_7/XI0/XI0_30/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_14 XI11_7/net21_1_ xsel_30_ XI11_7/XI0/XI0_30/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_13 XI11_7/net21_2_ xsel_30_ XI11_7/XI0/XI0_30/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_12 XI11_7/net21_3_ xsel_30_ XI11_7/XI0/XI0_30/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_11 XI11_7/net21_4_ xsel_30_ XI11_7/XI0/XI0_30/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_10 XI11_7/net21_5_ xsel_30_ XI11_7/XI0/XI0_30/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_9 XI11_7/net21_6_ xsel_30_ XI11_7/XI0/XI0_30/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_8 XI11_7/net21_7_ xsel_30_ XI11_7/XI0/XI0_30/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_7 XI11_7/net21_8_ xsel_30_ XI11_7/XI0/XI0_30/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_6 XI11_7/net21_9_ xsel_30_ XI11_7/XI0/XI0_30/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_5 XI11_7/net21_10_ xsel_30_ XI11_7/XI0/XI0_30/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_4 XI11_7/net21_11_ xsel_30_ XI11_7/XI0/XI0_30/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_3 XI11_7/net21_12_ xsel_30_ XI11_7/XI0/XI0_30/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_2 XI11_7/net21_13_ xsel_30_ XI11_7/XI0/XI0_30/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_1 XI11_7/net21_14_ xsel_30_ XI11_7/XI0/XI0_30/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN0_0 XI11_7/net21_15_ xsel_30_ XI11_7/XI0/XI0_30/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_15 XI11_7/XI0/XI0_30/d__15_ xsel_30_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_14 XI11_7/XI0/XI0_30/d__14_ xsel_30_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_13 XI11_7/XI0/XI0_30/d__13_ xsel_30_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_12 XI11_7/XI0/XI0_30/d__12_ xsel_30_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_11 XI11_7/XI0/XI0_30/d__11_ xsel_30_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_10 XI11_7/XI0/XI0_30/d__10_ xsel_30_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_9 XI11_7/XI0/XI0_30/d__9_ xsel_30_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_8 XI11_7/XI0/XI0_30/d__8_ xsel_30_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_7 XI11_7/XI0/XI0_30/d__7_ xsel_30_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_6 XI11_7/XI0/XI0_30/d__6_ xsel_30_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_5 XI11_7/XI0/XI0_30/d__5_ xsel_30_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_4 XI11_7/XI0/XI0_30/d__4_ xsel_30_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_3 XI11_7/XI0/XI0_30/d__3_ xsel_30_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_2 XI11_7/XI0/XI0_30/d__2_ xsel_30_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_1 XI11_7/XI0/XI0_30/d__1_ xsel_30_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_30/MN1_0 XI11_7/XI0/XI0_30/d__0_ xsel_30_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_15 XI11_7/net21_0_ xsel_29_ XI11_7/XI0/XI0_29/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_14 XI11_7/net21_1_ xsel_29_ XI11_7/XI0/XI0_29/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_13 XI11_7/net21_2_ xsel_29_ XI11_7/XI0/XI0_29/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_12 XI11_7/net21_3_ xsel_29_ XI11_7/XI0/XI0_29/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_11 XI11_7/net21_4_ xsel_29_ XI11_7/XI0/XI0_29/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_10 XI11_7/net21_5_ xsel_29_ XI11_7/XI0/XI0_29/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_9 XI11_7/net21_6_ xsel_29_ XI11_7/XI0/XI0_29/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_8 XI11_7/net21_7_ xsel_29_ XI11_7/XI0/XI0_29/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_7 XI11_7/net21_8_ xsel_29_ XI11_7/XI0/XI0_29/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_6 XI11_7/net21_9_ xsel_29_ XI11_7/XI0/XI0_29/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_5 XI11_7/net21_10_ xsel_29_ XI11_7/XI0/XI0_29/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_4 XI11_7/net21_11_ xsel_29_ XI11_7/XI0/XI0_29/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_3 XI11_7/net21_12_ xsel_29_ XI11_7/XI0/XI0_29/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_2 XI11_7/net21_13_ xsel_29_ XI11_7/XI0/XI0_29/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_1 XI11_7/net21_14_ xsel_29_ XI11_7/XI0/XI0_29/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN0_0 XI11_7/net21_15_ xsel_29_ XI11_7/XI0/XI0_29/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_15 XI11_7/XI0/XI0_29/d__15_ xsel_29_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_14 XI11_7/XI0/XI0_29/d__14_ xsel_29_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_13 XI11_7/XI0/XI0_29/d__13_ xsel_29_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_12 XI11_7/XI0/XI0_29/d__12_ xsel_29_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_11 XI11_7/XI0/XI0_29/d__11_ xsel_29_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_10 XI11_7/XI0/XI0_29/d__10_ xsel_29_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_9 XI11_7/XI0/XI0_29/d__9_ xsel_29_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_8 XI11_7/XI0/XI0_29/d__8_ xsel_29_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_7 XI11_7/XI0/XI0_29/d__7_ xsel_29_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_6 XI11_7/XI0/XI0_29/d__6_ xsel_29_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_5 XI11_7/XI0/XI0_29/d__5_ xsel_29_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_4 XI11_7/XI0/XI0_29/d__4_ xsel_29_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_3 XI11_7/XI0/XI0_29/d__3_ xsel_29_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_2 XI11_7/XI0/XI0_29/d__2_ xsel_29_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_1 XI11_7/XI0/XI0_29/d__1_ xsel_29_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_29/MN1_0 XI11_7/XI0/XI0_29/d__0_ xsel_29_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_15 XI11_7/net21_0_ xsel_28_ XI11_7/XI0/XI0_28/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_14 XI11_7/net21_1_ xsel_28_ XI11_7/XI0/XI0_28/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_13 XI11_7/net21_2_ xsel_28_ XI11_7/XI0/XI0_28/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_12 XI11_7/net21_3_ xsel_28_ XI11_7/XI0/XI0_28/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_11 XI11_7/net21_4_ xsel_28_ XI11_7/XI0/XI0_28/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_10 XI11_7/net21_5_ xsel_28_ XI11_7/XI0/XI0_28/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_9 XI11_7/net21_6_ xsel_28_ XI11_7/XI0/XI0_28/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_8 XI11_7/net21_7_ xsel_28_ XI11_7/XI0/XI0_28/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_7 XI11_7/net21_8_ xsel_28_ XI11_7/XI0/XI0_28/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_6 XI11_7/net21_9_ xsel_28_ XI11_7/XI0/XI0_28/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_5 XI11_7/net21_10_ xsel_28_ XI11_7/XI0/XI0_28/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_4 XI11_7/net21_11_ xsel_28_ XI11_7/XI0/XI0_28/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_3 XI11_7/net21_12_ xsel_28_ XI11_7/XI0/XI0_28/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_2 XI11_7/net21_13_ xsel_28_ XI11_7/XI0/XI0_28/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_1 XI11_7/net21_14_ xsel_28_ XI11_7/XI0/XI0_28/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN0_0 XI11_7/net21_15_ xsel_28_ XI11_7/XI0/XI0_28/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_15 XI11_7/XI0/XI0_28/d__15_ xsel_28_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_14 XI11_7/XI0/XI0_28/d__14_ xsel_28_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_13 XI11_7/XI0/XI0_28/d__13_ xsel_28_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_12 XI11_7/XI0/XI0_28/d__12_ xsel_28_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_11 XI11_7/XI0/XI0_28/d__11_ xsel_28_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_10 XI11_7/XI0/XI0_28/d__10_ xsel_28_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_9 XI11_7/XI0/XI0_28/d__9_ xsel_28_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_8 XI11_7/XI0/XI0_28/d__8_ xsel_28_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_7 XI11_7/XI0/XI0_28/d__7_ xsel_28_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_6 XI11_7/XI0/XI0_28/d__6_ xsel_28_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_5 XI11_7/XI0/XI0_28/d__5_ xsel_28_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_4 XI11_7/XI0/XI0_28/d__4_ xsel_28_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_3 XI11_7/XI0/XI0_28/d__3_ xsel_28_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_2 XI11_7/XI0/XI0_28/d__2_ xsel_28_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_1 XI11_7/XI0/XI0_28/d__1_ xsel_28_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_28/MN1_0 XI11_7/XI0/XI0_28/d__0_ xsel_28_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_15 XI11_7/net21_0_ xsel_27_ XI11_7/XI0/XI0_27/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_14 XI11_7/net21_1_ xsel_27_ XI11_7/XI0/XI0_27/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_13 XI11_7/net21_2_ xsel_27_ XI11_7/XI0/XI0_27/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_12 XI11_7/net21_3_ xsel_27_ XI11_7/XI0/XI0_27/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_11 XI11_7/net21_4_ xsel_27_ XI11_7/XI0/XI0_27/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_10 XI11_7/net21_5_ xsel_27_ XI11_7/XI0/XI0_27/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_9 XI11_7/net21_6_ xsel_27_ XI11_7/XI0/XI0_27/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_8 XI11_7/net21_7_ xsel_27_ XI11_7/XI0/XI0_27/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_7 XI11_7/net21_8_ xsel_27_ XI11_7/XI0/XI0_27/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_6 XI11_7/net21_9_ xsel_27_ XI11_7/XI0/XI0_27/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_5 XI11_7/net21_10_ xsel_27_ XI11_7/XI0/XI0_27/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_4 XI11_7/net21_11_ xsel_27_ XI11_7/XI0/XI0_27/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_3 XI11_7/net21_12_ xsel_27_ XI11_7/XI0/XI0_27/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_2 XI11_7/net21_13_ xsel_27_ XI11_7/XI0/XI0_27/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_1 XI11_7/net21_14_ xsel_27_ XI11_7/XI0/XI0_27/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN0_0 XI11_7/net21_15_ xsel_27_ XI11_7/XI0/XI0_27/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_15 XI11_7/XI0/XI0_27/d__15_ xsel_27_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_14 XI11_7/XI0/XI0_27/d__14_ xsel_27_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_13 XI11_7/XI0/XI0_27/d__13_ xsel_27_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_12 XI11_7/XI0/XI0_27/d__12_ xsel_27_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_11 XI11_7/XI0/XI0_27/d__11_ xsel_27_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_10 XI11_7/XI0/XI0_27/d__10_ xsel_27_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_9 XI11_7/XI0/XI0_27/d__9_ xsel_27_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_8 XI11_7/XI0/XI0_27/d__8_ xsel_27_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_7 XI11_7/XI0/XI0_27/d__7_ xsel_27_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_6 XI11_7/XI0/XI0_27/d__6_ xsel_27_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_5 XI11_7/XI0/XI0_27/d__5_ xsel_27_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_4 XI11_7/XI0/XI0_27/d__4_ xsel_27_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_3 XI11_7/XI0/XI0_27/d__3_ xsel_27_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_2 XI11_7/XI0/XI0_27/d__2_ xsel_27_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_1 XI11_7/XI0/XI0_27/d__1_ xsel_27_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_27/MN1_0 XI11_7/XI0/XI0_27/d__0_ xsel_27_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_15 XI11_7/net21_0_ xsel_26_ XI11_7/XI0/XI0_26/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_14 XI11_7/net21_1_ xsel_26_ XI11_7/XI0/XI0_26/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_13 XI11_7/net21_2_ xsel_26_ XI11_7/XI0/XI0_26/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_12 XI11_7/net21_3_ xsel_26_ XI11_7/XI0/XI0_26/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_11 XI11_7/net21_4_ xsel_26_ XI11_7/XI0/XI0_26/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_10 XI11_7/net21_5_ xsel_26_ XI11_7/XI0/XI0_26/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_9 XI11_7/net21_6_ xsel_26_ XI11_7/XI0/XI0_26/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_8 XI11_7/net21_7_ xsel_26_ XI11_7/XI0/XI0_26/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_7 XI11_7/net21_8_ xsel_26_ XI11_7/XI0/XI0_26/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_6 XI11_7/net21_9_ xsel_26_ XI11_7/XI0/XI0_26/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_5 XI11_7/net21_10_ xsel_26_ XI11_7/XI0/XI0_26/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_4 XI11_7/net21_11_ xsel_26_ XI11_7/XI0/XI0_26/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_3 XI11_7/net21_12_ xsel_26_ XI11_7/XI0/XI0_26/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_2 XI11_7/net21_13_ xsel_26_ XI11_7/XI0/XI0_26/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_1 XI11_7/net21_14_ xsel_26_ XI11_7/XI0/XI0_26/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN0_0 XI11_7/net21_15_ xsel_26_ XI11_7/XI0/XI0_26/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_15 XI11_7/XI0/XI0_26/d__15_ xsel_26_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_14 XI11_7/XI0/XI0_26/d__14_ xsel_26_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_13 XI11_7/XI0/XI0_26/d__13_ xsel_26_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_12 XI11_7/XI0/XI0_26/d__12_ xsel_26_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_11 XI11_7/XI0/XI0_26/d__11_ xsel_26_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_10 XI11_7/XI0/XI0_26/d__10_ xsel_26_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_9 XI11_7/XI0/XI0_26/d__9_ xsel_26_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_8 XI11_7/XI0/XI0_26/d__8_ xsel_26_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_7 XI11_7/XI0/XI0_26/d__7_ xsel_26_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_6 XI11_7/XI0/XI0_26/d__6_ xsel_26_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_5 XI11_7/XI0/XI0_26/d__5_ xsel_26_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_4 XI11_7/XI0/XI0_26/d__4_ xsel_26_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_3 XI11_7/XI0/XI0_26/d__3_ xsel_26_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_2 XI11_7/XI0/XI0_26/d__2_ xsel_26_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_1 XI11_7/XI0/XI0_26/d__1_ xsel_26_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_26/MN1_0 XI11_7/XI0/XI0_26/d__0_ xsel_26_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_15 XI11_7/net21_0_ xsel_25_ XI11_7/XI0/XI0_25/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_14 XI11_7/net21_1_ xsel_25_ XI11_7/XI0/XI0_25/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_13 XI11_7/net21_2_ xsel_25_ XI11_7/XI0/XI0_25/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_12 XI11_7/net21_3_ xsel_25_ XI11_7/XI0/XI0_25/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_11 XI11_7/net21_4_ xsel_25_ XI11_7/XI0/XI0_25/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_10 XI11_7/net21_5_ xsel_25_ XI11_7/XI0/XI0_25/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_9 XI11_7/net21_6_ xsel_25_ XI11_7/XI0/XI0_25/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_8 XI11_7/net21_7_ xsel_25_ XI11_7/XI0/XI0_25/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_7 XI11_7/net21_8_ xsel_25_ XI11_7/XI0/XI0_25/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_6 XI11_7/net21_9_ xsel_25_ XI11_7/XI0/XI0_25/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_5 XI11_7/net21_10_ xsel_25_ XI11_7/XI0/XI0_25/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_4 XI11_7/net21_11_ xsel_25_ XI11_7/XI0/XI0_25/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_3 XI11_7/net21_12_ xsel_25_ XI11_7/XI0/XI0_25/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_2 XI11_7/net21_13_ xsel_25_ XI11_7/XI0/XI0_25/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_1 XI11_7/net21_14_ xsel_25_ XI11_7/XI0/XI0_25/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN0_0 XI11_7/net21_15_ xsel_25_ XI11_7/XI0/XI0_25/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_15 XI11_7/XI0/XI0_25/d__15_ xsel_25_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_14 XI11_7/XI0/XI0_25/d__14_ xsel_25_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_13 XI11_7/XI0/XI0_25/d__13_ xsel_25_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_12 XI11_7/XI0/XI0_25/d__12_ xsel_25_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_11 XI11_7/XI0/XI0_25/d__11_ xsel_25_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_10 XI11_7/XI0/XI0_25/d__10_ xsel_25_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_9 XI11_7/XI0/XI0_25/d__9_ xsel_25_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_8 XI11_7/XI0/XI0_25/d__8_ xsel_25_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_7 XI11_7/XI0/XI0_25/d__7_ xsel_25_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_6 XI11_7/XI0/XI0_25/d__6_ xsel_25_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_5 XI11_7/XI0/XI0_25/d__5_ xsel_25_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_4 XI11_7/XI0/XI0_25/d__4_ xsel_25_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_3 XI11_7/XI0/XI0_25/d__3_ xsel_25_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_2 XI11_7/XI0/XI0_25/d__2_ xsel_25_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_1 XI11_7/XI0/XI0_25/d__1_ xsel_25_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_25/MN1_0 XI11_7/XI0/XI0_25/d__0_ xsel_25_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_15 XI11_7/net21_0_ xsel_24_ XI11_7/XI0/XI0_24/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_14 XI11_7/net21_1_ xsel_24_ XI11_7/XI0/XI0_24/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_13 XI11_7/net21_2_ xsel_24_ XI11_7/XI0/XI0_24/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_12 XI11_7/net21_3_ xsel_24_ XI11_7/XI0/XI0_24/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_11 XI11_7/net21_4_ xsel_24_ XI11_7/XI0/XI0_24/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_10 XI11_7/net21_5_ xsel_24_ XI11_7/XI0/XI0_24/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_9 XI11_7/net21_6_ xsel_24_ XI11_7/XI0/XI0_24/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_8 XI11_7/net21_7_ xsel_24_ XI11_7/XI0/XI0_24/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_7 XI11_7/net21_8_ xsel_24_ XI11_7/XI0/XI0_24/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_6 XI11_7/net21_9_ xsel_24_ XI11_7/XI0/XI0_24/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_5 XI11_7/net21_10_ xsel_24_ XI11_7/XI0/XI0_24/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_4 XI11_7/net21_11_ xsel_24_ XI11_7/XI0/XI0_24/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_3 XI11_7/net21_12_ xsel_24_ XI11_7/XI0/XI0_24/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_2 XI11_7/net21_13_ xsel_24_ XI11_7/XI0/XI0_24/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_1 XI11_7/net21_14_ xsel_24_ XI11_7/XI0/XI0_24/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN0_0 XI11_7/net21_15_ xsel_24_ XI11_7/XI0/XI0_24/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_15 XI11_7/XI0/XI0_24/d__15_ xsel_24_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_14 XI11_7/XI0/XI0_24/d__14_ xsel_24_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_13 XI11_7/XI0/XI0_24/d__13_ xsel_24_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_12 XI11_7/XI0/XI0_24/d__12_ xsel_24_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_11 XI11_7/XI0/XI0_24/d__11_ xsel_24_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_10 XI11_7/XI0/XI0_24/d__10_ xsel_24_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_9 XI11_7/XI0/XI0_24/d__9_ xsel_24_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_8 XI11_7/XI0/XI0_24/d__8_ xsel_24_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_7 XI11_7/XI0/XI0_24/d__7_ xsel_24_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_6 XI11_7/XI0/XI0_24/d__6_ xsel_24_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_5 XI11_7/XI0/XI0_24/d__5_ xsel_24_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_4 XI11_7/XI0/XI0_24/d__4_ xsel_24_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_3 XI11_7/XI0/XI0_24/d__3_ xsel_24_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_2 XI11_7/XI0/XI0_24/d__2_ xsel_24_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_1 XI11_7/XI0/XI0_24/d__1_ xsel_24_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_24/MN1_0 XI11_7/XI0/XI0_24/d__0_ xsel_24_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_15 XI11_7/net21_0_ xsel_23_ XI11_7/XI0/XI0_23/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_14 XI11_7/net21_1_ xsel_23_ XI11_7/XI0/XI0_23/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_13 XI11_7/net21_2_ xsel_23_ XI11_7/XI0/XI0_23/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_12 XI11_7/net21_3_ xsel_23_ XI11_7/XI0/XI0_23/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_11 XI11_7/net21_4_ xsel_23_ XI11_7/XI0/XI0_23/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_10 XI11_7/net21_5_ xsel_23_ XI11_7/XI0/XI0_23/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_9 XI11_7/net21_6_ xsel_23_ XI11_7/XI0/XI0_23/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_8 XI11_7/net21_7_ xsel_23_ XI11_7/XI0/XI0_23/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_7 XI11_7/net21_8_ xsel_23_ XI11_7/XI0/XI0_23/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_6 XI11_7/net21_9_ xsel_23_ XI11_7/XI0/XI0_23/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_5 XI11_7/net21_10_ xsel_23_ XI11_7/XI0/XI0_23/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_4 XI11_7/net21_11_ xsel_23_ XI11_7/XI0/XI0_23/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_3 XI11_7/net21_12_ xsel_23_ XI11_7/XI0/XI0_23/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_2 XI11_7/net21_13_ xsel_23_ XI11_7/XI0/XI0_23/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_1 XI11_7/net21_14_ xsel_23_ XI11_7/XI0/XI0_23/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN0_0 XI11_7/net21_15_ xsel_23_ XI11_7/XI0/XI0_23/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_15 XI11_7/XI0/XI0_23/d__15_ xsel_23_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_14 XI11_7/XI0/XI0_23/d__14_ xsel_23_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_13 XI11_7/XI0/XI0_23/d__13_ xsel_23_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_12 XI11_7/XI0/XI0_23/d__12_ xsel_23_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_11 XI11_7/XI0/XI0_23/d__11_ xsel_23_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_10 XI11_7/XI0/XI0_23/d__10_ xsel_23_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_9 XI11_7/XI0/XI0_23/d__9_ xsel_23_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_8 XI11_7/XI0/XI0_23/d__8_ xsel_23_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_7 XI11_7/XI0/XI0_23/d__7_ xsel_23_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_6 XI11_7/XI0/XI0_23/d__6_ xsel_23_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_5 XI11_7/XI0/XI0_23/d__5_ xsel_23_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_4 XI11_7/XI0/XI0_23/d__4_ xsel_23_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_3 XI11_7/XI0/XI0_23/d__3_ xsel_23_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_2 XI11_7/XI0/XI0_23/d__2_ xsel_23_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_1 XI11_7/XI0/XI0_23/d__1_ xsel_23_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_23/MN1_0 XI11_7/XI0/XI0_23/d__0_ xsel_23_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_15 XI11_7/net21_0_ xsel_22_ XI11_7/XI0/XI0_22/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_14 XI11_7/net21_1_ xsel_22_ XI11_7/XI0/XI0_22/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_13 XI11_7/net21_2_ xsel_22_ XI11_7/XI0/XI0_22/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_12 XI11_7/net21_3_ xsel_22_ XI11_7/XI0/XI0_22/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_11 XI11_7/net21_4_ xsel_22_ XI11_7/XI0/XI0_22/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_10 XI11_7/net21_5_ xsel_22_ XI11_7/XI0/XI0_22/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_9 XI11_7/net21_6_ xsel_22_ XI11_7/XI0/XI0_22/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_8 XI11_7/net21_7_ xsel_22_ XI11_7/XI0/XI0_22/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_7 XI11_7/net21_8_ xsel_22_ XI11_7/XI0/XI0_22/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_6 XI11_7/net21_9_ xsel_22_ XI11_7/XI0/XI0_22/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_5 XI11_7/net21_10_ xsel_22_ XI11_7/XI0/XI0_22/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_4 XI11_7/net21_11_ xsel_22_ XI11_7/XI0/XI0_22/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_3 XI11_7/net21_12_ xsel_22_ XI11_7/XI0/XI0_22/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_2 XI11_7/net21_13_ xsel_22_ XI11_7/XI0/XI0_22/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_1 XI11_7/net21_14_ xsel_22_ XI11_7/XI0/XI0_22/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN0_0 XI11_7/net21_15_ xsel_22_ XI11_7/XI0/XI0_22/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_15 XI11_7/XI0/XI0_22/d__15_ xsel_22_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_14 XI11_7/XI0/XI0_22/d__14_ xsel_22_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_13 XI11_7/XI0/XI0_22/d__13_ xsel_22_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_12 XI11_7/XI0/XI0_22/d__12_ xsel_22_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_11 XI11_7/XI0/XI0_22/d__11_ xsel_22_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_10 XI11_7/XI0/XI0_22/d__10_ xsel_22_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_9 XI11_7/XI0/XI0_22/d__9_ xsel_22_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_8 XI11_7/XI0/XI0_22/d__8_ xsel_22_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_7 XI11_7/XI0/XI0_22/d__7_ xsel_22_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_6 XI11_7/XI0/XI0_22/d__6_ xsel_22_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_5 XI11_7/XI0/XI0_22/d__5_ xsel_22_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_4 XI11_7/XI0/XI0_22/d__4_ xsel_22_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_3 XI11_7/XI0/XI0_22/d__3_ xsel_22_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_2 XI11_7/XI0/XI0_22/d__2_ xsel_22_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_1 XI11_7/XI0/XI0_22/d__1_ xsel_22_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_22/MN1_0 XI11_7/XI0/XI0_22/d__0_ xsel_22_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_15 XI11_7/net21_0_ xsel_21_ XI11_7/XI0/XI0_21/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_14 XI11_7/net21_1_ xsel_21_ XI11_7/XI0/XI0_21/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_13 XI11_7/net21_2_ xsel_21_ XI11_7/XI0/XI0_21/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_12 XI11_7/net21_3_ xsel_21_ XI11_7/XI0/XI0_21/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_11 XI11_7/net21_4_ xsel_21_ XI11_7/XI0/XI0_21/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_10 XI11_7/net21_5_ xsel_21_ XI11_7/XI0/XI0_21/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_9 XI11_7/net21_6_ xsel_21_ XI11_7/XI0/XI0_21/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_8 XI11_7/net21_7_ xsel_21_ XI11_7/XI0/XI0_21/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_7 XI11_7/net21_8_ xsel_21_ XI11_7/XI0/XI0_21/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_6 XI11_7/net21_9_ xsel_21_ XI11_7/XI0/XI0_21/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_5 XI11_7/net21_10_ xsel_21_ XI11_7/XI0/XI0_21/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_4 XI11_7/net21_11_ xsel_21_ XI11_7/XI0/XI0_21/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_3 XI11_7/net21_12_ xsel_21_ XI11_7/XI0/XI0_21/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_2 XI11_7/net21_13_ xsel_21_ XI11_7/XI0/XI0_21/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_1 XI11_7/net21_14_ xsel_21_ XI11_7/XI0/XI0_21/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN0_0 XI11_7/net21_15_ xsel_21_ XI11_7/XI0/XI0_21/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_15 XI11_7/XI0/XI0_21/d__15_ xsel_21_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_14 XI11_7/XI0/XI0_21/d__14_ xsel_21_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_13 XI11_7/XI0/XI0_21/d__13_ xsel_21_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_12 XI11_7/XI0/XI0_21/d__12_ xsel_21_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_11 XI11_7/XI0/XI0_21/d__11_ xsel_21_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_10 XI11_7/XI0/XI0_21/d__10_ xsel_21_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_9 XI11_7/XI0/XI0_21/d__9_ xsel_21_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_8 XI11_7/XI0/XI0_21/d__8_ xsel_21_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_7 XI11_7/XI0/XI0_21/d__7_ xsel_21_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_6 XI11_7/XI0/XI0_21/d__6_ xsel_21_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_5 XI11_7/XI0/XI0_21/d__5_ xsel_21_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_4 XI11_7/XI0/XI0_21/d__4_ xsel_21_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_3 XI11_7/XI0/XI0_21/d__3_ xsel_21_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_2 XI11_7/XI0/XI0_21/d__2_ xsel_21_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_1 XI11_7/XI0/XI0_21/d__1_ xsel_21_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_21/MN1_0 XI11_7/XI0/XI0_21/d__0_ xsel_21_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_15 XI11_7/net21_0_ xsel_20_ XI11_7/XI0/XI0_20/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_14 XI11_7/net21_1_ xsel_20_ XI11_7/XI0/XI0_20/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_13 XI11_7/net21_2_ xsel_20_ XI11_7/XI0/XI0_20/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_12 XI11_7/net21_3_ xsel_20_ XI11_7/XI0/XI0_20/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_11 XI11_7/net21_4_ xsel_20_ XI11_7/XI0/XI0_20/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_10 XI11_7/net21_5_ xsel_20_ XI11_7/XI0/XI0_20/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_9 XI11_7/net21_6_ xsel_20_ XI11_7/XI0/XI0_20/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_8 XI11_7/net21_7_ xsel_20_ XI11_7/XI0/XI0_20/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_7 XI11_7/net21_8_ xsel_20_ XI11_7/XI0/XI0_20/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_6 XI11_7/net21_9_ xsel_20_ XI11_7/XI0/XI0_20/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_5 XI11_7/net21_10_ xsel_20_ XI11_7/XI0/XI0_20/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_4 XI11_7/net21_11_ xsel_20_ XI11_7/XI0/XI0_20/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_3 XI11_7/net21_12_ xsel_20_ XI11_7/XI0/XI0_20/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_2 XI11_7/net21_13_ xsel_20_ XI11_7/XI0/XI0_20/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_1 XI11_7/net21_14_ xsel_20_ XI11_7/XI0/XI0_20/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN0_0 XI11_7/net21_15_ xsel_20_ XI11_7/XI0/XI0_20/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_15 XI11_7/XI0/XI0_20/d__15_ xsel_20_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_14 XI11_7/XI0/XI0_20/d__14_ xsel_20_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_13 XI11_7/XI0/XI0_20/d__13_ xsel_20_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_12 XI11_7/XI0/XI0_20/d__12_ xsel_20_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_11 XI11_7/XI0/XI0_20/d__11_ xsel_20_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_10 XI11_7/XI0/XI0_20/d__10_ xsel_20_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_9 XI11_7/XI0/XI0_20/d__9_ xsel_20_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_8 XI11_7/XI0/XI0_20/d__8_ xsel_20_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_7 XI11_7/XI0/XI0_20/d__7_ xsel_20_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_6 XI11_7/XI0/XI0_20/d__6_ xsel_20_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_5 XI11_7/XI0/XI0_20/d__5_ xsel_20_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_4 XI11_7/XI0/XI0_20/d__4_ xsel_20_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_3 XI11_7/XI0/XI0_20/d__3_ xsel_20_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_2 XI11_7/XI0/XI0_20/d__2_ xsel_20_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_1 XI11_7/XI0/XI0_20/d__1_ xsel_20_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_20/MN1_0 XI11_7/XI0/XI0_20/d__0_ xsel_20_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_15 XI11_7/net21_0_ xsel_19_ XI11_7/XI0/XI0_19/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_14 XI11_7/net21_1_ xsel_19_ XI11_7/XI0/XI0_19/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_13 XI11_7/net21_2_ xsel_19_ XI11_7/XI0/XI0_19/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_12 XI11_7/net21_3_ xsel_19_ XI11_7/XI0/XI0_19/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_11 XI11_7/net21_4_ xsel_19_ XI11_7/XI0/XI0_19/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_10 XI11_7/net21_5_ xsel_19_ XI11_7/XI0/XI0_19/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_9 XI11_7/net21_6_ xsel_19_ XI11_7/XI0/XI0_19/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_8 XI11_7/net21_7_ xsel_19_ XI11_7/XI0/XI0_19/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_7 XI11_7/net21_8_ xsel_19_ XI11_7/XI0/XI0_19/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_6 XI11_7/net21_9_ xsel_19_ XI11_7/XI0/XI0_19/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_5 XI11_7/net21_10_ xsel_19_ XI11_7/XI0/XI0_19/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_4 XI11_7/net21_11_ xsel_19_ XI11_7/XI0/XI0_19/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_3 XI11_7/net21_12_ xsel_19_ XI11_7/XI0/XI0_19/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_2 XI11_7/net21_13_ xsel_19_ XI11_7/XI0/XI0_19/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_1 XI11_7/net21_14_ xsel_19_ XI11_7/XI0/XI0_19/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN0_0 XI11_7/net21_15_ xsel_19_ XI11_7/XI0/XI0_19/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_15 XI11_7/XI0/XI0_19/d__15_ xsel_19_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_14 XI11_7/XI0/XI0_19/d__14_ xsel_19_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_13 XI11_7/XI0/XI0_19/d__13_ xsel_19_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_12 XI11_7/XI0/XI0_19/d__12_ xsel_19_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_11 XI11_7/XI0/XI0_19/d__11_ xsel_19_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_10 XI11_7/XI0/XI0_19/d__10_ xsel_19_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_9 XI11_7/XI0/XI0_19/d__9_ xsel_19_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_8 XI11_7/XI0/XI0_19/d__8_ xsel_19_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_7 XI11_7/XI0/XI0_19/d__7_ xsel_19_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_6 XI11_7/XI0/XI0_19/d__6_ xsel_19_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_5 XI11_7/XI0/XI0_19/d__5_ xsel_19_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_4 XI11_7/XI0/XI0_19/d__4_ xsel_19_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_3 XI11_7/XI0/XI0_19/d__3_ xsel_19_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_2 XI11_7/XI0/XI0_19/d__2_ xsel_19_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_1 XI11_7/XI0/XI0_19/d__1_ xsel_19_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_19/MN1_0 XI11_7/XI0/XI0_19/d__0_ xsel_19_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_15 XI11_7/net21_0_ xsel_18_ XI11_7/XI0/XI0_18/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_14 XI11_7/net21_1_ xsel_18_ XI11_7/XI0/XI0_18/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_13 XI11_7/net21_2_ xsel_18_ XI11_7/XI0/XI0_18/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_12 XI11_7/net21_3_ xsel_18_ XI11_7/XI0/XI0_18/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_11 XI11_7/net21_4_ xsel_18_ XI11_7/XI0/XI0_18/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_10 XI11_7/net21_5_ xsel_18_ XI11_7/XI0/XI0_18/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_9 XI11_7/net21_6_ xsel_18_ XI11_7/XI0/XI0_18/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_8 XI11_7/net21_7_ xsel_18_ XI11_7/XI0/XI0_18/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_7 XI11_7/net21_8_ xsel_18_ XI11_7/XI0/XI0_18/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_6 XI11_7/net21_9_ xsel_18_ XI11_7/XI0/XI0_18/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_5 XI11_7/net21_10_ xsel_18_ XI11_7/XI0/XI0_18/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_4 XI11_7/net21_11_ xsel_18_ XI11_7/XI0/XI0_18/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_3 XI11_7/net21_12_ xsel_18_ XI11_7/XI0/XI0_18/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_2 XI11_7/net21_13_ xsel_18_ XI11_7/XI0/XI0_18/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_1 XI11_7/net21_14_ xsel_18_ XI11_7/XI0/XI0_18/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN0_0 XI11_7/net21_15_ xsel_18_ XI11_7/XI0/XI0_18/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_15 XI11_7/XI0/XI0_18/d__15_ xsel_18_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_14 XI11_7/XI0/XI0_18/d__14_ xsel_18_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_13 XI11_7/XI0/XI0_18/d__13_ xsel_18_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_12 XI11_7/XI0/XI0_18/d__12_ xsel_18_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_11 XI11_7/XI0/XI0_18/d__11_ xsel_18_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_10 XI11_7/XI0/XI0_18/d__10_ xsel_18_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_9 XI11_7/XI0/XI0_18/d__9_ xsel_18_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_8 XI11_7/XI0/XI0_18/d__8_ xsel_18_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_7 XI11_7/XI0/XI0_18/d__7_ xsel_18_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_6 XI11_7/XI0/XI0_18/d__6_ xsel_18_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_5 XI11_7/XI0/XI0_18/d__5_ xsel_18_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_4 XI11_7/XI0/XI0_18/d__4_ xsel_18_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_3 XI11_7/XI0/XI0_18/d__3_ xsel_18_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_2 XI11_7/XI0/XI0_18/d__2_ xsel_18_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_1 XI11_7/XI0/XI0_18/d__1_ xsel_18_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_18/MN1_0 XI11_7/XI0/XI0_18/d__0_ xsel_18_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_15 XI11_7/net21_0_ xsel_17_ XI11_7/XI0/XI0_17/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_14 XI11_7/net21_1_ xsel_17_ XI11_7/XI0/XI0_17/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_13 XI11_7/net21_2_ xsel_17_ XI11_7/XI0/XI0_17/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_12 XI11_7/net21_3_ xsel_17_ XI11_7/XI0/XI0_17/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_11 XI11_7/net21_4_ xsel_17_ XI11_7/XI0/XI0_17/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_10 XI11_7/net21_5_ xsel_17_ XI11_7/XI0/XI0_17/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_9 XI11_7/net21_6_ xsel_17_ XI11_7/XI0/XI0_17/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_8 XI11_7/net21_7_ xsel_17_ XI11_7/XI0/XI0_17/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_7 XI11_7/net21_8_ xsel_17_ XI11_7/XI0/XI0_17/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_6 XI11_7/net21_9_ xsel_17_ XI11_7/XI0/XI0_17/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_5 XI11_7/net21_10_ xsel_17_ XI11_7/XI0/XI0_17/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_4 XI11_7/net21_11_ xsel_17_ XI11_7/XI0/XI0_17/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_3 XI11_7/net21_12_ xsel_17_ XI11_7/XI0/XI0_17/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_2 XI11_7/net21_13_ xsel_17_ XI11_7/XI0/XI0_17/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_1 XI11_7/net21_14_ xsel_17_ XI11_7/XI0/XI0_17/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN0_0 XI11_7/net21_15_ xsel_17_ XI11_7/XI0/XI0_17/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_15 XI11_7/XI0/XI0_17/d__15_ xsel_17_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_14 XI11_7/XI0/XI0_17/d__14_ xsel_17_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_13 XI11_7/XI0/XI0_17/d__13_ xsel_17_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_12 XI11_7/XI0/XI0_17/d__12_ xsel_17_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_11 XI11_7/XI0/XI0_17/d__11_ xsel_17_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_10 XI11_7/XI0/XI0_17/d__10_ xsel_17_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_9 XI11_7/XI0/XI0_17/d__9_ xsel_17_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_8 XI11_7/XI0/XI0_17/d__8_ xsel_17_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_7 XI11_7/XI0/XI0_17/d__7_ xsel_17_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_6 XI11_7/XI0/XI0_17/d__6_ xsel_17_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_5 XI11_7/XI0/XI0_17/d__5_ xsel_17_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_4 XI11_7/XI0/XI0_17/d__4_ xsel_17_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_3 XI11_7/XI0/XI0_17/d__3_ xsel_17_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_2 XI11_7/XI0/XI0_17/d__2_ xsel_17_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_1 XI11_7/XI0/XI0_17/d__1_ xsel_17_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_17/MN1_0 XI11_7/XI0/XI0_17/d__0_ xsel_17_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_15 XI11_7/net21_0_ xsel_16_ XI11_7/XI0/XI0_16/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_14 XI11_7/net21_1_ xsel_16_ XI11_7/XI0/XI0_16/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_13 XI11_7/net21_2_ xsel_16_ XI11_7/XI0/XI0_16/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_12 XI11_7/net21_3_ xsel_16_ XI11_7/XI0/XI0_16/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_11 XI11_7/net21_4_ xsel_16_ XI11_7/XI0/XI0_16/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_10 XI11_7/net21_5_ xsel_16_ XI11_7/XI0/XI0_16/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_9 XI11_7/net21_6_ xsel_16_ XI11_7/XI0/XI0_16/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_8 XI11_7/net21_7_ xsel_16_ XI11_7/XI0/XI0_16/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_7 XI11_7/net21_8_ xsel_16_ XI11_7/XI0/XI0_16/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_6 XI11_7/net21_9_ xsel_16_ XI11_7/XI0/XI0_16/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_5 XI11_7/net21_10_ xsel_16_ XI11_7/XI0/XI0_16/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_4 XI11_7/net21_11_ xsel_16_ XI11_7/XI0/XI0_16/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_3 XI11_7/net21_12_ xsel_16_ XI11_7/XI0/XI0_16/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_2 XI11_7/net21_13_ xsel_16_ XI11_7/XI0/XI0_16/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_1 XI11_7/net21_14_ xsel_16_ XI11_7/XI0/XI0_16/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN0_0 XI11_7/net21_15_ xsel_16_ XI11_7/XI0/XI0_16/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_15 XI11_7/XI0/XI0_16/d__15_ xsel_16_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_14 XI11_7/XI0/XI0_16/d__14_ xsel_16_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_13 XI11_7/XI0/XI0_16/d__13_ xsel_16_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_12 XI11_7/XI0/XI0_16/d__12_ xsel_16_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_11 XI11_7/XI0/XI0_16/d__11_ xsel_16_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_10 XI11_7/XI0/XI0_16/d__10_ xsel_16_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_9 XI11_7/XI0/XI0_16/d__9_ xsel_16_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_8 XI11_7/XI0/XI0_16/d__8_ xsel_16_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_7 XI11_7/XI0/XI0_16/d__7_ xsel_16_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_6 XI11_7/XI0/XI0_16/d__6_ xsel_16_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_5 XI11_7/XI0/XI0_16/d__5_ xsel_16_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_4 XI11_7/XI0/XI0_16/d__4_ xsel_16_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_3 XI11_7/XI0/XI0_16/d__3_ xsel_16_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_2 XI11_7/XI0/XI0_16/d__2_ xsel_16_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_1 XI11_7/XI0/XI0_16/d__1_ xsel_16_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_16/MN1_0 XI11_7/XI0/XI0_16/d__0_ xsel_16_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_15 XI11_7/net21_0_ xsel_15_ XI11_7/XI0/XI0_15/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_14 XI11_7/net21_1_ xsel_15_ XI11_7/XI0/XI0_15/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_13 XI11_7/net21_2_ xsel_15_ XI11_7/XI0/XI0_15/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_12 XI11_7/net21_3_ xsel_15_ XI11_7/XI0/XI0_15/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_11 XI11_7/net21_4_ xsel_15_ XI11_7/XI0/XI0_15/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_10 XI11_7/net21_5_ xsel_15_ XI11_7/XI0/XI0_15/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_9 XI11_7/net21_6_ xsel_15_ XI11_7/XI0/XI0_15/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_8 XI11_7/net21_7_ xsel_15_ XI11_7/XI0/XI0_15/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_7 XI11_7/net21_8_ xsel_15_ XI11_7/XI0/XI0_15/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_6 XI11_7/net21_9_ xsel_15_ XI11_7/XI0/XI0_15/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_5 XI11_7/net21_10_ xsel_15_ XI11_7/XI0/XI0_15/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_4 XI11_7/net21_11_ xsel_15_ XI11_7/XI0/XI0_15/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_3 XI11_7/net21_12_ xsel_15_ XI11_7/XI0/XI0_15/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_2 XI11_7/net21_13_ xsel_15_ XI11_7/XI0/XI0_15/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_1 XI11_7/net21_14_ xsel_15_ XI11_7/XI0/XI0_15/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN0_0 XI11_7/net21_15_ xsel_15_ XI11_7/XI0/XI0_15/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_15 XI11_7/XI0/XI0_15/d__15_ xsel_15_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_14 XI11_7/XI0/XI0_15/d__14_ xsel_15_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_13 XI11_7/XI0/XI0_15/d__13_ xsel_15_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_12 XI11_7/XI0/XI0_15/d__12_ xsel_15_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_11 XI11_7/XI0/XI0_15/d__11_ xsel_15_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_10 XI11_7/XI0/XI0_15/d__10_ xsel_15_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_9 XI11_7/XI0/XI0_15/d__9_ xsel_15_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_8 XI11_7/XI0/XI0_15/d__8_ xsel_15_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_7 XI11_7/XI0/XI0_15/d__7_ xsel_15_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_6 XI11_7/XI0/XI0_15/d__6_ xsel_15_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_5 XI11_7/XI0/XI0_15/d__5_ xsel_15_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_4 XI11_7/XI0/XI0_15/d__4_ xsel_15_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_3 XI11_7/XI0/XI0_15/d__3_ xsel_15_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_2 XI11_7/XI0/XI0_15/d__2_ xsel_15_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_1 XI11_7/XI0/XI0_15/d__1_ xsel_15_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_15/MN1_0 XI11_7/XI0/XI0_15/d__0_ xsel_15_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_15 XI11_7/net21_0_ xsel_14_ XI11_7/XI0/XI0_14/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_14 XI11_7/net21_1_ xsel_14_ XI11_7/XI0/XI0_14/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_13 XI11_7/net21_2_ xsel_14_ XI11_7/XI0/XI0_14/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_12 XI11_7/net21_3_ xsel_14_ XI11_7/XI0/XI0_14/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_11 XI11_7/net21_4_ xsel_14_ XI11_7/XI0/XI0_14/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_10 XI11_7/net21_5_ xsel_14_ XI11_7/XI0/XI0_14/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_9 XI11_7/net21_6_ xsel_14_ XI11_7/XI0/XI0_14/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_8 XI11_7/net21_7_ xsel_14_ XI11_7/XI0/XI0_14/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_7 XI11_7/net21_8_ xsel_14_ XI11_7/XI0/XI0_14/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_6 XI11_7/net21_9_ xsel_14_ XI11_7/XI0/XI0_14/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_5 XI11_7/net21_10_ xsel_14_ XI11_7/XI0/XI0_14/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_4 XI11_7/net21_11_ xsel_14_ XI11_7/XI0/XI0_14/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_3 XI11_7/net21_12_ xsel_14_ XI11_7/XI0/XI0_14/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_2 XI11_7/net21_13_ xsel_14_ XI11_7/XI0/XI0_14/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_1 XI11_7/net21_14_ xsel_14_ XI11_7/XI0/XI0_14/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN0_0 XI11_7/net21_15_ xsel_14_ XI11_7/XI0/XI0_14/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_15 XI11_7/XI0/XI0_14/d__15_ xsel_14_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_14 XI11_7/XI0/XI0_14/d__14_ xsel_14_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_13 XI11_7/XI0/XI0_14/d__13_ xsel_14_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_12 XI11_7/XI0/XI0_14/d__12_ xsel_14_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_11 XI11_7/XI0/XI0_14/d__11_ xsel_14_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_10 XI11_7/XI0/XI0_14/d__10_ xsel_14_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_9 XI11_7/XI0/XI0_14/d__9_ xsel_14_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_8 XI11_7/XI0/XI0_14/d__8_ xsel_14_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_7 XI11_7/XI0/XI0_14/d__7_ xsel_14_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_6 XI11_7/XI0/XI0_14/d__6_ xsel_14_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_5 XI11_7/XI0/XI0_14/d__5_ xsel_14_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_4 XI11_7/XI0/XI0_14/d__4_ xsel_14_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_3 XI11_7/XI0/XI0_14/d__3_ xsel_14_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_2 XI11_7/XI0/XI0_14/d__2_ xsel_14_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_1 XI11_7/XI0/XI0_14/d__1_ xsel_14_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_14/MN1_0 XI11_7/XI0/XI0_14/d__0_ xsel_14_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_15 XI11_7/net21_0_ xsel_13_ XI11_7/XI0/XI0_13/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_14 XI11_7/net21_1_ xsel_13_ XI11_7/XI0/XI0_13/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_13 XI11_7/net21_2_ xsel_13_ XI11_7/XI0/XI0_13/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_12 XI11_7/net21_3_ xsel_13_ XI11_7/XI0/XI0_13/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_11 XI11_7/net21_4_ xsel_13_ XI11_7/XI0/XI0_13/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_10 XI11_7/net21_5_ xsel_13_ XI11_7/XI0/XI0_13/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_9 XI11_7/net21_6_ xsel_13_ XI11_7/XI0/XI0_13/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_8 XI11_7/net21_7_ xsel_13_ XI11_7/XI0/XI0_13/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_7 XI11_7/net21_8_ xsel_13_ XI11_7/XI0/XI0_13/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_6 XI11_7/net21_9_ xsel_13_ XI11_7/XI0/XI0_13/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_5 XI11_7/net21_10_ xsel_13_ XI11_7/XI0/XI0_13/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_4 XI11_7/net21_11_ xsel_13_ XI11_7/XI0/XI0_13/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_3 XI11_7/net21_12_ xsel_13_ XI11_7/XI0/XI0_13/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_2 XI11_7/net21_13_ xsel_13_ XI11_7/XI0/XI0_13/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_1 XI11_7/net21_14_ xsel_13_ XI11_7/XI0/XI0_13/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN0_0 XI11_7/net21_15_ xsel_13_ XI11_7/XI0/XI0_13/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_15 XI11_7/XI0/XI0_13/d__15_ xsel_13_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_14 XI11_7/XI0/XI0_13/d__14_ xsel_13_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_13 XI11_7/XI0/XI0_13/d__13_ xsel_13_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_12 XI11_7/XI0/XI0_13/d__12_ xsel_13_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_11 XI11_7/XI0/XI0_13/d__11_ xsel_13_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_10 XI11_7/XI0/XI0_13/d__10_ xsel_13_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_9 XI11_7/XI0/XI0_13/d__9_ xsel_13_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_8 XI11_7/XI0/XI0_13/d__8_ xsel_13_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_7 XI11_7/XI0/XI0_13/d__7_ xsel_13_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_6 XI11_7/XI0/XI0_13/d__6_ xsel_13_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_5 XI11_7/XI0/XI0_13/d__5_ xsel_13_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_4 XI11_7/XI0/XI0_13/d__4_ xsel_13_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_3 XI11_7/XI0/XI0_13/d__3_ xsel_13_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_2 XI11_7/XI0/XI0_13/d__2_ xsel_13_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_1 XI11_7/XI0/XI0_13/d__1_ xsel_13_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_13/MN1_0 XI11_7/XI0/XI0_13/d__0_ xsel_13_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_15 XI11_7/net21_0_ xsel_12_ XI11_7/XI0/XI0_12/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_14 XI11_7/net21_1_ xsel_12_ XI11_7/XI0/XI0_12/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_13 XI11_7/net21_2_ xsel_12_ XI11_7/XI0/XI0_12/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_12 XI11_7/net21_3_ xsel_12_ XI11_7/XI0/XI0_12/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_11 XI11_7/net21_4_ xsel_12_ XI11_7/XI0/XI0_12/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_10 XI11_7/net21_5_ xsel_12_ XI11_7/XI0/XI0_12/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_9 XI11_7/net21_6_ xsel_12_ XI11_7/XI0/XI0_12/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_8 XI11_7/net21_7_ xsel_12_ XI11_7/XI0/XI0_12/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_7 XI11_7/net21_8_ xsel_12_ XI11_7/XI0/XI0_12/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_6 XI11_7/net21_9_ xsel_12_ XI11_7/XI0/XI0_12/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_5 XI11_7/net21_10_ xsel_12_ XI11_7/XI0/XI0_12/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_4 XI11_7/net21_11_ xsel_12_ XI11_7/XI0/XI0_12/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_3 XI11_7/net21_12_ xsel_12_ XI11_7/XI0/XI0_12/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_2 XI11_7/net21_13_ xsel_12_ XI11_7/XI0/XI0_12/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_1 XI11_7/net21_14_ xsel_12_ XI11_7/XI0/XI0_12/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN0_0 XI11_7/net21_15_ xsel_12_ XI11_7/XI0/XI0_12/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_15 XI11_7/XI0/XI0_12/d__15_ xsel_12_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_14 XI11_7/XI0/XI0_12/d__14_ xsel_12_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_13 XI11_7/XI0/XI0_12/d__13_ xsel_12_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_12 XI11_7/XI0/XI0_12/d__12_ xsel_12_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_11 XI11_7/XI0/XI0_12/d__11_ xsel_12_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_10 XI11_7/XI0/XI0_12/d__10_ xsel_12_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_9 XI11_7/XI0/XI0_12/d__9_ xsel_12_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_8 XI11_7/XI0/XI0_12/d__8_ xsel_12_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_7 XI11_7/XI0/XI0_12/d__7_ xsel_12_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_6 XI11_7/XI0/XI0_12/d__6_ xsel_12_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_5 XI11_7/XI0/XI0_12/d__5_ xsel_12_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_4 XI11_7/XI0/XI0_12/d__4_ xsel_12_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_3 XI11_7/XI0/XI0_12/d__3_ xsel_12_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_2 XI11_7/XI0/XI0_12/d__2_ xsel_12_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_1 XI11_7/XI0/XI0_12/d__1_ xsel_12_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_12/MN1_0 XI11_7/XI0/XI0_12/d__0_ xsel_12_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_15 XI11_7/net21_0_ xsel_11_ XI11_7/XI0/XI0_11/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_14 XI11_7/net21_1_ xsel_11_ XI11_7/XI0/XI0_11/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_13 XI11_7/net21_2_ xsel_11_ XI11_7/XI0/XI0_11/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_12 XI11_7/net21_3_ xsel_11_ XI11_7/XI0/XI0_11/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_11 XI11_7/net21_4_ xsel_11_ XI11_7/XI0/XI0_11/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_10 XI11_7/net21_5_ xsel_11_ XI11_7/XI0/XI0_11/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_9 XI11_7/net21_6_ xsel_11_ XI11_7/XI0/XI0_11/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_8 XI11_7/net21_7_ xsel_11_ XI11_7/XI0/XI0_11/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_7 XI11_7/net21_8_ xsel_11_ XI11_7/XI0/XI0_11/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_6 XI11_7/net21_9_ xsel_11_ XI11_7/XI0/XI0_11/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_5 XI11_7/net21_10_ xsel_11_ XI11_7/XI0/XI0_11/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_4 XI11_7/net21_11_ xsel_11_ XI11_7/XI0/XI0_11/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_3 XI11_7/net21_12_ xsel_11_ XI11_7/XI0/XI0_11/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_2 XI11_7/net21_13_ xsel_11_ XI11_7/XI0/XI0_11/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_1 XI11_7/net21_14_ xsel_11_ XI11_7/XI0/XI0_11/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN0_0 XI11_7/net21_15_ xsel_11_ XI11_7/XI0/XI0_11/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_15 XI11_7/XI0/XI0_11/d__15_ xsel_11_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_14 XI11_7/XI0/XI0_11/d__14_ xsel_11_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_13 XI11_7/XI0/XI0_11/d__13_ xsel_11_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_12 XI11_7/XI0/XI0_11/d__12_ xsel_11_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_11 XI11_7/XI0/XI0_11/d__11_ xsel_11_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_10 XI11_7/XI0/XI0_11/d__10_ xsel_11_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_9 XI11_7/XI0/XI0_11/d__9_ xsel_11_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_8 XI11_7/XI0/XI0_11/d__8_ xsel_11_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_7 XI11_7/XI0/XI0_11/d__7_ xsel_11_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_6 XI11_7/XI0/XI0_11/d__6_ xsel_11_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_5 XI11_7/XI0/XI0_11/d__5_ xsel_11_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_4 XI11_7/XI0/XI0_11/d__4_ xsel_11_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_3 XI11_7/XI0/XI0_11/d__3_ xsel_11_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_2 XI11_7/XI0/XI0_11/d__2_ xsel_11_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_1 XI11_7/XI0/XI0_11/d__1_ xsel_11_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_11/MN1_0 XI11_7/XI0/XI0_11/d__0_ xsel_11_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_15 XI11_7/net21_0_ xsel_10_ XI11_7/XI0/XI0_10/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_14 XI11_7/net21_1_ xsel_10_ XI11_7/XI0/XI0_10/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_13 XI11_7/net21_2_ xsel_10_ XI11_7/XI0/XI0_10/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_12 XI11_7/net21_3_ xsel_10_ XI11_7/XI0/XI0_10/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_11 XI11_7/net21_4_ xsel_10_ XI11_7/XI0/XI0_10/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_10 XI11_7/net21_5_ xsel_10_ XI11_7/XI0/XI0_10/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_9 XI11_7/net21_6_ xsel_10_ XI11_7/XI0/XI0_10/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_8 XI11_7/net21_7_ xsel_10_ XI11_7/XI0/XI0_10/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_7 XI11_7/net21_8_ xsel_10_ XI11_7/XI0/XI0_10/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_6 XI11_7/net21_9_ xsel_10_ XI11_7/XI0/XI0_10/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_5 XI11_7/net21_10_ xsel_10_ XI11_7/XI0/XI0_10/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_4 XI11_7/net21_11_ xsel_10_ XI11_7/XI0/XI0_10/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_3 XI11_7/net21_12_ xsel_10_ XI11_7/XI0/XI0_10/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_2 XI11_7/net21_13_ xsel_10_ XI11_7/XI0/XI0_10/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_1 XI11_7/net21_14_ xsel_10_ XI11_7/XI0/XI0_10/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN0_0 XI11_7/net21_15_ xsel_10_ XI11_7/XI0/XI0_10/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_15 XI11_7/XI0/XI0_10/d__15_ xsel_10_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_14 XI11_7/XI0/XI0_10/d__14_ xsel_10_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_13 XI11_7/XI0/XI0_10/d__13_ xsel_10_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_12 XI11_7/XI0/XI0_10/d__12_ xsel_10_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_11 XI11_7/XI0/XI0_10/d__11_ xsel_10_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_10 XI11_7/XI0/XI0_10/d__10_ xsel_10_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_9 XI11_7/XI0/XI0_10/d__9_ xsel_10_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_8 XI11_7/XI0/XI0_10/d__8_ xsel_10_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_7 XI11_7/XI0/XI0_10/d__7_ xsel_10_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_6 XI11_7/XI0/XI0_10/d__6_ xsel_10_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_5 XI11_7/XI0/XI0_10/d__5_ xsel_10_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_4 XI11_7/XI0/XI0_10/d__4_ xsel_10_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_3 XI11_7/XI0/XI0_10/d__3_ xsel_10_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_2 XI11_7/XI0/XI0_10/d__2_ xsel_10_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_1 XI11_7/XI0/XI0_10/d__1_ xsel_10_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_10/MN1_0 XI11_7/XI0/XI0_10/d__0_ xsel_10_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_15 XI11_7/net21_0_ xsel_9_ XI11_7/XI0/XI0_9/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_14 XI11_7/net21_1_ xsel_9_ XI11_7/XI0/XI0_9/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_13 XI11_7/net21_2_ xsel_9_ XI11_7/XI0/XI0_9/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_12 XI11_7/net21_3_ xsel_9_ XI11_7/XI0/XI0_9/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_11 XI11_7/net21_4_ xsel_9_ XI11_7/XI0/XI0_9/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_10 XI11_7/net21_5_ xsel_9_ XI11_7/XI0/XI0_9/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_9 XI11_7/net21_6_ xsel_9_ XI11_7/XI0/XI0_9/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_8 XI11_7/net21_7_ xsel_9_ XI11_7/XI0/XI0_9/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_7 XI11_7/net21_8_ xsel_9_ XI11_7/XI0/XI0_9/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_6 XI11_7/net21_9_ xsel_9_ XI11_7/XI0/XI0_9/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_5 XI11_7/net21_10_ xsel_9_ XI11_7/XI0/XI0_9/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_4 XI11_7/net21_11_ xsel_9_ XI11_7/XI0/XI0_9/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_3 XI11_7/net21_12_ xsel_9_ XI11_7/XI0/XI0_9/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_2 XI11_7/net21_13_ xsel_9_ XI11_7/XI0/XI0_9/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_1 XI11_7/net21_14_ xsel_9_ XI11_7/XI0/XI0_9/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN0_0 XI11_7/net21_15_ xsel_9_ XI11_7/XI0/XI0_9/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_15 XI11_7/XI0/XI0_9/d__15_ xsel_9_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_14 XI11_7/XI0/XI0_9/d__14_ xsel_9_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_13 XI11_7/XI0/XI0_9/d__13_ xsel_9_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_12 XI11_7/XI0/XI0_9/d__12_ xsel_9_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_11 XI11_7/XI0/XI0_9/d__11_ xsel_9_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_10 XI11_7/XI0/XI0_9/d__10_ xsel_9_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_9 XI11_7/XI0/XI0_9/d__9_ xsel_9_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_8 XI11_7/XI0/XI0_9/d__8_ xsel_9_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_7 XI11_7/XI0/XI0_9/d__7_ xsel_9_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_6 XI11_7/XI0/XI0_9/d__6_ xsel_9_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_5 XI11_7/XI0/XI0_9/d__5_ xsel_9_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_4 XI11_7/XI0/XI0_9/d__4_ xsel_9_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_3 XI11_7/XI0/XI0_9/d__3_ xsel_9_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_2 XI11_7/XI0/XI0_9/d__2_ xsel_9_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_1 XI11_7/XI0/XI0_9/d__1_ xsel_9_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_9/MN1_0 XI11_7/XI0/XI0_9/d__0_ xsel_9_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_15 XI11_7/net21_0_ xsel_8_ XI11_7/XI0/XI0_8/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_14 XI11_7/net21_1_ xsel_8_ XI11_7/XI0/XI0_8/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_13 XI11_7/net21_2_ xsel_8_ XI11_7/XI0/XI0_8/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_12 XI11_7/net21_3_ xsel_8_ XI11_7/XI0/XI0_8/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_11 XI11_7/net21_4_ xsel_8_ XI11_7/XI0/XI0_8/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_10 XI11_7/net21_5_ xsel_8_ XI11_7/XI0/XI0_8/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_9 XI11_7/net21_6_ xsel_8_ XI11_7/XI0/XI0_8/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_8 XI11_7/net21_7_ xsel_8_ XI11_7/XI0/XI0_8/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_7 XI11_7/net21_8_ xsel_8_ XI11_7/XI0/XI0_8/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_6 XI11_7/net21_9_ xsel_8_ XI11_7/XI0/XI0_8/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_5 XI11_7/net21_10_ xsel_8_ XI11_7/XI0/XI0_8/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_4 XI11_7/net21_11_ xsel_8_ XI11_7/XI0/XI0_8/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_3 XI11_7/net21_12_ xsel_8_ XI11_7/XI0/XI0_8/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_2 XI11_7/net21_13_ xsel_8_ XI11_7/XI0/XI0_8/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_1 XI11_7/net21_14_ xsel_8_ XI11_7/XI0/XI0_8/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN0_0 XI11_7/net21_15_ xsel_8_ XI11_7/XI0/XI0_8/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_15 XI11_7/XI0/XI0_8/d__15_ xsel_8_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_14 XI11_7/XI0/XI0_8/d__14_ xsel_8_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_13 XI11_7/XI0/XI0_8/d__13_ xsel_8_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_12 XI11_7/XI0/XI0_8/d__12_ xsel_8_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_11 XI11_7/XI0/XI0_8/d__11_ xsel_8_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_10 XI11_7/XI0/XI0_8/d__10_ xsel_8_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_9 XI11_7/XI0/XI0_8/d__9_ xsel_8_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_8 XI11_7/XI0/XI0_8/d__8_ xsel_8_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_7 XI11_7/XI0/XI0_8/d__7_ xsel_8_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_6 XI11_7/XI0/XI0_8/d__6_ xsel_8_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_5 XI11_7/XI0/XI0_8/d__5_ xsel_8_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_4 XI11_7/XI0/XI0_8/d__4_ xsel_8_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_3 XI11_7/XI0/XI0_8/d__3_ xsel_8_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_2 XI11_7/XI0/XI0_8/d__2_ xsel_8_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_1 XI11_7/XI0/XI0_8/d__1_ xsel_8_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_8/MN1_0 XI11_7/XI0/XI0_8/d__0_ xsel_8_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_15 XI11_7/net21_0_ xsel_7_ XI11_7/XI0/XI0_7/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_14 XI11_7/net21_1_ xsel_7_ XI11_7/XI0/XI0_7/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_13 XI11_7/net21_2_ xsel_7_ XI11_7/XI0/XI0_7/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_12 XI11_7/net21_3_ xsel_7_ XI11_7/XI0/XI0_7/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_11 XI11_7/net21_4_ xsel_7_ XI11_7/XI0/XI0_7/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_10 XI11_7/net21_5_ xsel_7_ XI11_7/XI0/XI0_7/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_9 XI11_7/net21_6_ xsel_7_ XI11_7/XI0/XI0_7/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_8 XI11_7/net21_7_ xsel_7_ XI11_7/XI0/XI0_7/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_7 XI11_7/net21_8_ xsel_7_ XI11_7/XI0/XI0_7/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_6 XI11_7/net21_9_ xsel_7_ XI11_7/XI0/XI0_7/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_5 XI11_7/net21_10_ xsel_7_ XI11_7/XI0/XI0_7/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_4 XI11_7/net21_11_ xsel_7_ XI11_7/XI0/XI0_7/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_3 XI11_7/net21_12_ xsel_7_ XI11_7/XI0/XI0_7/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_2 XI11_7/net21_13_ xsel_7_ XI11_7/XI0/XI0_7/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_1 XI11_7/net21_14_ xsel_7_ XI11_7/XI0/XI0_7/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN0_0 XI11_7/net21_15_ xsel_7_ XI11_7/XI0/XI0_7/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_15 XI11_7/XI0/XI0_7/d__15_ xsel_7_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_14 XI11_7/XI0/XI0_7/d__14_ xsel_7_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_13 XI11_7/XI0/XI0_7/d__13_ xsel_7_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_12 XI11_7/XI0/XI0_7/d__12_ xsel_7_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_11 XI11_7/XI0/XI0_7/d__11_ xsel_7_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_10 XI11_7/XI0/XI0_7/d__10_ xsel_7_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_9 XI11_7/XI0/XI0_7/d__9_ xsel_7_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_8 XI11_7/XI0/XI0_7/d__8_ xsel_7_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_7 XI11_7/XI0/XI0_7/d__7_ xsel_7_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_6 XI11_7/XI0/XI0_7/d__6_ xsel_7_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_5 XI11_7/XI0/XI0_7/d__5_ xsel_7_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_4 XI11_7/XI0/XI0_7/d__4_ xsel_7_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_3 XI11_7/XI0/XI0_7/d__3_ xsel_7_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_2 XI11_7/XI0/XI0_7/d__2_ xsel_7_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_1 XI11_7/XI0/XI0_7/d__1_ xsel_7_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_7/MN1_0 XI11_7/XI0/XI0_7/d__0_ xsel_7_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_15 XI11_7/net21_0_ xsel_6_ XI11_7/XI0/XI0_6/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_14 XI11_7/net21_1_ xsel_6_ XI11_7/XI0/XI0_6/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_13 XI11_7/net21_2_ xsel_6_ XI11_7/XI0/XI0_6/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_12 XI11_7/net21_3_ xsel_6_ XI11_7/XI0/XI0_6/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_11 XI11_7/net21_4_ xsel_6_ XI11_7/XI0/XI0_6/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_10 XI11_7/net21_5_ xsel_6_ XI11_7/XI0/XI0_6/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_9 XI11_7/net21_6_ xsel_6_ XI11_7/XI0/XI0_6/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_8 XI11_7/net21_7_ xsel_6_ XI11_7/XI0/XI0_6/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_7 XI11_7/net21_8_ xsel_6_ XI11_7/XI0/XI0_6/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_6 XI11_7/net21_9_ xsel_6_ XI11_7/XI0/XI0_6/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_5 XI11_7/net21_10_ xsel_6_ XI11_7/XI0/XI0_6/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_4 XI11_7/net21_11_ xsel_6_ XI11_7/XI0/XI0_6/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_3 XI11_7/net21_12_ xsel_6_ XI11_7/XI0/XI0_6/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_2 XI11_7/net21_13_ xsel_6_ XI11_7/XI0/XI0_6/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_1 XI11_7/net21_14_ xsel_6_ XI11_7/XI0/XI0_6/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN0_0 XI11_7/net21_15_ xsel_6_ XI11_7/XI0/XI0_6/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_15 XI11_7/XI0/XI0_6/d__15_ xsel_6_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_14 XI11_7/XI0/XI0_6/d__14_ xsel_6_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_13 XI11_7/XI0/XI0_6/d__13_ xsel_6_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_12 XI11_7/XI0/XI0_6/d__12_ xsel_6_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_11 XI11_7/XI0/XI0_6/d__11_ xsel_6_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_10 XI11_7/XI0/XI0_6/d__10_ xsel_6_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_9 XI11_7/XI0/XI0_6/d__9_ xsel_6_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_8 XI11_7/XI0/XI0_6/d__8_ xsel_6_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_7 XI11_7/XI0/XI0_6/d__7_ xsel_6_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_6 XI11_7/XI0/XI0_6/d__6_ xsel_6_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_5 XI11_7/XI0/XI0_6/d__5_ xsel_6_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_4 XI11_7/XI0/XI0_6/d__4_ xsel_6_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_3 XI11_7/XI0/XI0_6/d__3_ xsel_6_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_2 XI11_7/XI0/XI0_6/d__2_ xsel_6_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_1 XI11_7/XI0/XI0_6/d__1_ xsel_6_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_6/MN1_0 XI11_7/XI0/XI0_6/d__0_ xsel_6_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_15 XI11_7/net21_0_ xsel_5_ XI11_7/XI0/XI0_5/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_14 XI11_7/net21_1_ xsel_5_ XI11_7/XI0/XI0_5/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_13 XI11_7/net21_2_ xsel_5_ XI11_7/XI0/XI0_5/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_12 XI11_7/net21_3_ xsel_5_ XI11_7/XI0/XI0_5/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_11 XI11_7/net21_4_ xsel_5_ XI11_7/XI0/XI0_5/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_10 XI11_7/net21_5_ xsel_5_ XI11_7/XI0/XI0_5/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_9 XI11_7/net21_6_ xsel_5_ XI11_7/XI0/XI0_5/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_8 XI11_7/net21_7_ xsel_5_ XI11_7/XI0/XI0_5/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_7 XI11_7/net21_8_ xsel_5_ XI11_7/XI0/XI0_5/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_6 XI11_7/net21_9_ xsel_5_ XI11_7/XI0/XI0_5/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_5 XI11_7/net21_10_ xsel_5_ XI11_7/XI0/XI0_5/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_4 XI11_7/net21_11_ xsel_5_ XI11_7/XI0/XI0_5/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_3 XI11_7/net21_12_ xsel_5_ XI11_7/XI0/XI0_5/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_2 XI11_7/net21_13_ xsel_5_ XI11_7/XI0/XI0_5/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_1 XI11_7/net21_14_ xsel_5_ XI11_7/XI0/XI0_5/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN0_0 XI11_7/net21_15_ xsel_5_ XI11_7/XI0/XI0_5/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_15 XI11_7/XI0/XI0_5/d__15_ xsel_5_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_14 XI11_7/XI0/XI0_5/d__14_ xsel_5_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_13 XI11_7/XI0/XI0_5/d__13_ xsel_5_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_12 XI11_7/XI0/XI0_5/d__12_ xsel_5_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_11 XI11_7/XI0/XI0_5/d__11_ xsel_5_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_10 XI11_7/XI0/XI0_5/d__10_ xsel_5_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_9 XI11_7/XI0/XI0_5/d__9_ xsel_5_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_8 XI11_7/XI0/XI0_5/d__8_ xsel_5_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_7 XI11_7/XI0/XI0_5/d__7_ xsel_5_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_6 XI11_7/XI0/XI0_5/d__6_ xsel_5_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_5 XI11_7/XI0/XI0_5/d__5_ xsel_5_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_4 XI11_7/XI0/XI0_5/d__4_ xsel_5_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_3 XI11_7/XI0/XI0_5/d__3_ xsel_5_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_2 XI11_7/XI0/XI0_5/d__2_ xsel_5_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_1 XI11_7/XI0/XI0_5/d__1_ xsel_5_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_5/MN1_0 XI11_7/XI0/XI0_5/d__0_ xsel_5_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_15 XI11_7/net21_0_ xsel_4_ XI11_7/XI0/XI0_4/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_14 XI11_7/net21_1_ xsel_4_ XI11_7/XI0/XI0_4/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_13 XI11_7/net21_2_ xsel_4_ XI11_7/XI0/XI0_4/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_12 XI11_7/net21_3_ xsel_4_ XI11_7/XI0/XI0_4/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_11 XI11_7/net21_4_ xsel_4_ XI11_7/XI0/XI0_4/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_10 XI11_7/net21_5_ xsel_4_ XI11_7/XI0/XI0_4/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_9 XI11_7/net21_6_ xsel_4_ XI11_7/XI0/XI0_4/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_8 XI11_7/net21_7_ xsel_4_ XI11_7/XI0/XI0_4/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_7 XI11_7/net21_8_ xsel_4_ XI11_7/XI0/XI0_4/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_6 XI11_7/net21_9_ xsel_4_ XI11_7/XI0/XI0_4/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_5 XI11_7/net21_10_ xsel_4_ XI11_7/XI0/XI0_4/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_4 XI11_7/net21_11_ xsel_4_ XI11_7/XI0/XI0_4/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_3 XI11_7/net21_12_ xsel_4_ XI11_7/XI0/XI0_4/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_2 XI11_7/net21_13_ xsel_4_ XI11_7/XI0/XI0_4/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_1 XI11_7/net21_14_ xsel_4_ XI11_7/XI0/XI0_4/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN0_0 XI11_7/net21_15_ xsel_4_ XI11_7/XI0/XI0_4/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_15 XI11_7/XI0/XI0_4/d__15_ xsel_4_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_14 XI11_7/XI0/XI0_4/d__14_ xsel_4_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_13 XI11_7/XI0/XI0_4/d__13_ xsel_4_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_12 XI11_7/XI0/XI0_4/d__12_ xsel_4_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_11 XI11_7/XI0/XI0_4/d__11_ xsel_4_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_10 XI11_7/XI0/XI0_4/d__10_ xsel_4_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_9 XI11_7/XI0/XI0_4/d__9_ xsel_4_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_8 XI11_7/XI0/XI0_4/d__8_ xsel_4_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_7 XI11_7/XI0/XI0_4/d__7_ xsel_4_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_6 XI11_7/XI0/XI0_4/d__6_ xsel_4_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_5 XI11_7/XI0/XI0_4/d__5_ xsel_4_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_4 XI11_7/XI0/XI0_4/d__4_ xsel_4_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_3 XI11_7/XI0/XI0_4/d__3_ xsel_4_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_2 XI11_7/XI0/XI0_4/d__2_ xsel_4_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_1 XI11_7/XI0/XI0_4/d__1_ xsel_4_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_4/MN1_0 XI11_7/XI0/XI0_4/d__0_ xsel_4_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_15 XI11_7/net21_0_ xsel_3_ XI11_7/XI0/XI0_3/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_14 XI11_7/net21_1_ xsel_3_ XI11_7/XI0/XI0_3/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_13 XI11_7/net21_2_ xsel_3_ XI11_7/XI0/XI0_3/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_12 XI11_7/net21_3_ xsel_3_ XI11_7/XI0/XI0_3/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_11 XI11_7/net21_4_ xsel_3_ XI11_7/XI0/XI0_3/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_10 XI11_7/net21_5_ xsel_3_ XI11_7/XI0/XI0_3/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_9 XI11_7/net21_6_ xsel_3_ XI11_7/XI0/XI0_3/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_8 XI11_7/net21_7_ xsel_3_ XI11_7/XI0/XI0_3/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_7 XI11_7/net21_8_ xsel_3_ XI11_7/XI0/XI0_3/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_6 XI11_7/net21_9_ xsel_3_ XI11_7/XI0/XI0_3/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_5 XI11_7/net21_10_ xsel_3_ XI11_7/XI0/XI0_3/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_4 XI11_7/net21_11_ xsel_3_ XI11_7/XI0/XI0_3/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_3 XI11_7/net21_12_ xsel_3_ XI11_7/XI0/XI0_3/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_2 XI11_7/net21_13_ xsel_3_ XI11_7/XI0/XI0_3/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_1 XI11_7/net21_14_ xsel_3_ XI11_7/XI0/XI0_3/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN0_0 XI11_7/net21_15_ xsel_3_ XI11_7/XI0/XI0_3/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_15 XI11_7/XI0/XI0_3/d__15_ xsel_3_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_14 XI11_7/XI0/XI0_3/d__14_ xsel_3_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_13 XI11_7/XI0/XI0_3/d__13_ xsel_3_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_12 XI11_7/XI0/XI0_3/d__12_ xsel_3_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_11 XI11_7/XI0/XI0_3/d__11_ xsel_3_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_10 XI11_7/XI0/XI0_3/d__10_ xsel_3_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_9 XI11_7/XI0/XI0_3/d__9_ xsel_3_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_8 XI11_7/XI0/XI0_3/d__8_ xsel_3_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_7 XI11_7/XI0/XI0_3/d__7_ xsel_3_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_6 XI11_7/XI0/XI0_3/d__6_ xsel_3_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_5 XI11_7/XI0/XI0_3/d__5_ xsel_3_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_4 XI11_7/XI0/XI0_3/d__4_ xsel_3_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_3 XI11_7/XI0/XI0_3/d__3_ xsel_3_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_2 XI11_7/XI0/XI0_3/d__2_ xsel_3_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_1 XI11_7/XI0/XI0_3/d__1_ xsel_3_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_3/MN1_0 XI11_7/XI0/XI0_3/d__0_ xsel_3_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_15 XI11_7/net21_0_ xsel_2_ XI11_7/XI0/XI0_2/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_14 XI11_7/net21_1_ xsel_2_ XI11_7/XI0/XI0_2/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_13 XI11_7/net21_2_ xsel_2_ XI11_7/XI0/XI0_2/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_12 XI11_7/net21_3_ xsel_2_ XI11_7/XI0/XI0_2/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_11 XI11_7/net21_4_ xsel_2_ XI11_7/XI0/XI0_2/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_10 XI11_7/net21_5_ xsel_2_ XI11_7/XI0/XI0_2/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_9 XI11_7/net21_6_ xsel_2_ XI11_7/XI0/XI0_2/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_8 XI11_7/net21_7_ xsel_2_ XI11_7/XI0/XI0_2/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_7 XI11_7/net21_8_ xsel_2_ XI11_7/XI0/XI0_2/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_6 XI11_7/net21_9_ xsel_2_ XI11_7/XI0/XI0_2/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_5 XI11_7/net21_10_ xsel_2_ XI11_7/XI0/XI0_2/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_4 XI11_7/net21_11_ xsel_2_ XI11_7/XI0/XI0_2/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_3 XI11_7/net21_12_ xsel_2_ XI11_7/XI0/XI0_2/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_2 XI11_7/net21_13_ xsel_2_ XI11_7/XI0/XI0_2/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_1 XI11_7/net21_14_ xsel_2_ XI11_7/XI0/XI0_2/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN0_0 XI11_7/net21_15_ xsel_2_ XI11_7/XI0/XI0_2/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_15 XI11_7/XI0/XI0_2/d__15_ xsel_2_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_14 XI11_7/XI0/XI0_2/d__14_ xsel_2_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_13 XI11_7/XI0/XI0_2/d__13_ xsel_2_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_12 XI11_7/XI0/XI0_2/d__12_ xsel_2_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_11 XI11_7/XI0/XI0_2/d__11_ xsel_2_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_10 XI11_7/XI0/XI0_2/d__10_ xsel_2_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_9 XI11_7/XI0/XI0_2/d__9_ xsel_2_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_8 XI11_7/XI0/XI0_2/d__8_ xsel_2_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_7 XI11_7/XI0/XI0_2/d__7_ xsel_2_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_6 XI11_7/XI0/XI0_2/d__6_ xsel_2_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_5 XI11_7/XI0/XI0_2/d__5_ xsel_2_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_4 XI11_7/XI0/XI0_2/d__4_ xsel_2_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_3 XI11_7/XI0/XI0_2/d__3_ xsel_2_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_2 XI11_7/XI0/XI0_2/d__2_ xsel_2_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_1 XI11_7/XI0/XI0_2/d__1_ xsel_2_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_2/MN1_0 XI11_7/XI0/XI0_2/d__0_ xsel_2_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_15 XI11_7/net21_0_ xsel_1_ XI11_7/XI0/XI0_1/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_14 XI11_7/net21_1_ xsel_1_ XI11_7/XI0/XI0_1/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_13 XI11_7/net21_2_ xsel_1_ XI11_7/XI0/XI0_1/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_12 XI11_7/net21_3_ xsel_1_ XI11_7/XI0/XI0_1/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_11 XI11_7/net21_4_ xsel_1_ XI11_7/XI0/XI0_1/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_10 XI11_7/net21_5_ xsel_1_ XI11_7/XI0/XI0_1/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_9 XI11_7/net21_6_ xsel_1_ XI11_7/XI0/XI0_1/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_8 XI11_7/net21_7_ xsel_1_ XI11_7/XI0/XI0_1/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_7 XI11_7/net21_8_ xsel_1_ XI11_7/XI0/XI0_1/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_6 XI11_7/net21_9_ xsel_1_ XI11_7/XI0/XI0_1/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_5 XI11_7/net21_10_ xsel_1_ XI11_7/XI0/XI0_1/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_4 XI11_7/net21_11_ xsel_1_ XI11_7/XI0/XI0_1/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_3 XI11_7/net21_12_ xsel_1_ XI11_7/XI0/XI0_1/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_2 XI11_7/net21_13_ xsel_1_ XI11_7/XI0/XI0_1/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_1 XI11_7/net21_14_ xsel_1_ XI11_7/XI0/XI0_1/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN0_0 XI11_7/net21_15_ xsel_1_ XI11_7/XI0/XI0_1/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_15 XI11_7/XI0/XI0_1/d__15_ xsel_1_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_14 XI11_7/XI0/XI0_1/d__14_ xsel_1_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_13 XI11_7/XI0/XI0_1/d__13_ xsel_1_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_12 XI11_7/XI0/XI0_1/d__12_ xsel_1_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_11 XI11_7/XI0/XI0_1/d__11_ xsel_1_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_10 XI11_7/XI0/XI0_1/d__10_ xsel_1_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_9 XI11_7/XI0/XI0_1/d__9_ xsel_1_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_8 XI11_7/XI0/XI0_1/d__8_ xsel_1_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_7 XI11_7/XI0/XI0_1/d__7_ xsel_1_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_6 XI11_7/XI0/XI0_1/d__6_ xsel_1_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_5 XI11_7/XI0/XI0_1/d__5_ xsel_1_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_4 XI11_7/XI0/XI0_1/d__4_ xsel_1_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_3 XI11_7/XI0/XI0_1/d__3_ xsel_1_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_2 XI11_7/XI0/XI0_1/d__2_ xsel_1_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_1 XI11_7/XI0/XI0_1/d__1_ xsel_1_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_1/MN1_0 XI11_7/XI0/XI0_1/d__0_ xsel_1_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_15 XI11_7/net21_0_ xsel_0_ XI11_7/XI0/XI0_0/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_14 XI11_7/net21_1_ xsel_0_ XI11_7/XI0/XI0_0/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_13 XI11_7/net21_2_ xsel_0_ XI11_7/XI0/XI0_0/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_12 XI11_7/net21_3_ xsel_0_ XI11_7/XI0/XI0_0/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_11 XI11_7/net21_4_ xsel_0_ XI11_7/XI0/XI0_0/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_10 XI11_7/net21_5_ xsel_0_ XI11_7/XI0/XI0_0/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_9 XI11_7/net21_6_ xsel_0_ XI11_7/XI0/XI0_0/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_8 XI11_7/net21_7_ xsel_0_ XI11_7/XI0/XI0_0/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_7 XI11_7/net21_8_ xsel_0_ XI11_7/XI0/XI0_0/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_6 XI11_7/net21_9_ xsel_0_ XI11_7/XI0/XI0_0/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_5 XI11_7/net21_10_ xsel_0_ XI11_7/XI0/XI0_0/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_4 XI11_7/net21_11_ xsel_0_ XI11_7/XI0/XI0_0/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_3 XI11_7/net21_12_ xsel_0_ XI11_7/XI0/XI0_0/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_2 XI11_7/net21_13_ xsel_0_ XI11_7/XI0/XI0_0/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_1 XI11_7/net21_14_ xsel_0_ XI11_7/XI0/XI0_0/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN0_0 XI11_7/net21_15_ xsel_0_ XI11_7/XI0/XI0_0/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_15 XI11_7/XI0/XI0_0/d__15_ xsel_0_ XI11_7/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_14 XI11_7/XI0/XI0_0/d__14_ xsel_0_ XI11_7/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_13 XI11_7/XI0/XI0_0/d__13_ xsel_0_ XI11_7/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_12 XI11_7/XI0/XI0_0/d__12_ xsel_0_ XI11_7/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_11 XI11_7/XI0/XI0_0/d__11_ xsel_0_ XI11_7/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_10 XI11_7/XI0/XI0_0/d__10_ xsel_0_ XI11_7/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_9 XI11_7/XI0/XI0_0/d__9_ xsel_0_ XI11_7/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_8 XI11_7/XI0/XI0_0/d__8_ xsel_0_ XI11_7/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_7 XI11_7/XI0/XI0_0/d__7_ xsel_0_ XI11_7/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_6 XI11_7/XI0/XI0_0/d__6_ xsel_0_ XI11_7/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_5 XI11_7/XI0/XI0_0/d__5_ xsel_0_ XI11_7/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_4 XI11_7/XI0/XI0_0/d__4_ xsel_0_ XI11_7/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_3 XI11_7/XI0/XI0_0/d__3_ xsel_0_ XI11_7/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_2 XI11_7/XI0/XI0_0/d__2_ xsel_0_ XI11_7/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_1 XI11_7/XI0/XI0_0/d__1_ xsel_0_ XI11_7/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_7/XI0/XI0_0/MN1_0 XI11_7/XI0/XI0_0/d__0_ xsel_0_ XI11_7/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI2/MN0_15 XI11_6/net21_0_ ysel_15_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_14 XI11_6/net21_1_ ysel_14_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_13 XI11_6/net21_2_ ysel_13_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_12 XI11_6/net21_3_ ysel_12_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_11 XI11_6/net21_4_ ysel_11_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_10 XI11_6/net21_5_ ysel_10_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_9 XI11_6/net21_6_ ysel_9_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_8 XI11_6/net21_7_ ysel_8_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_7 XI11_6/net21_8_ ysel_7_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_6 XI11_6/net21_9_ ysel_6_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_5 XI11_6/net21_10_ ysel_5_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_4 XI11_6/net21_11_ ysel_4_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_3 XI11_6/net21_12_ ysel_3_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_2 XI11_6/net21_13_ ysel_2_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_1 XI11_6/net21_14_ ysel_1_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN0_0 XI11_6/net21_15_ ysel_0_ XI11_6/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_15 XI11_6/net20_0_ ysel_15_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_14 XI11_6/net20_1_ ysel_14_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_13 XI11_6/net20_2_ ysel_13_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_12 XI11_6/net20_3_ ysel_12_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_11 XI11_6/net20_4_ ysel_11_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_10 XI11_6/net20_5_ ysel_10_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_9 XI11_6/net20_6_ ysel_9_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_8 XI11_6/net20_7_ ysel_8_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_7 XI11_6/net20_8_ ysel_7_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_6 XI11_6/net20_9_ ysel_6_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_5 XI11_6/net20_10_ ysel_5_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_4 XI11_6/net20_11_ ysel_4_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_3 XI11_6/net20_12_ ysel_3_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_2 XI11_6/net20_13_ ysel_2_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_1 XI11_6/net20_14_ ysel_1_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI2/MN1_0 XI11_6/net20_15_ ysel_0_ XI11_6/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_6/XI4/MN8 vdd XI11_6/XI4/net8 XI11_6/net12 vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_6/XI4/MP0 XI11_6/net9 XI11_6/XI4/net23 vdd vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_6/XI4/MP4 XI11_6/net12 XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI4/MP1 XI11_6/net9 XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI4/MP5 XI11_6/net12 XI11_6/preck XI11_6/net9 vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI4/MN7 vdd XI11_6/XI4/net090 DOUT_6_ vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_6/XI4/MP3 gnd XI11_6/XI4/net089 XI11_6/net12 gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_6/XI4/MN5 XI11_6/net9 XI11_6/XI4/net0103 gnd gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_6/XI4/MN4 XI11_6/XI4/data_out_ XI11_6/XI4/net32 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_6/XI4/MN0 XI11_6/XI4/data_out XI11_6/XI4/net52 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_6/XI4/MN9 gnd XI11_6/XI4/net0112 DOUT_6_ gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_6/XI1_15/MP2 XI11_6/net20_0_ XI11_6/preck XI11_6/net21_0_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_15/MP1 XI11_6/net20_0_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_15/MP0 XI11_6/net21_0_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_14/MP2 XI11_6/net20_1_ XI11_6/preck XI11_6/net21_1_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_14/MP1 XI11_6/net20_1_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_14/MP0 XI11_6/net21_1_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_13/MP2 XI11_6/net20_2_ XI11_6/preck XI11_6/net21_2_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_13/MP1 XI11_6/net20_2_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_13/MP0 XI11_6/net21_2_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_12/MP2 XI11_6/net20_3_ XI11_6/preck XI11_6/net21_3_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_12/MP1 XI11_6/net20_3_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_12/MP0 XI11_6/net21_3_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_11/MP2 XI11_6/net20_4_ XI11_6/preck XI11_6/net21_4_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_11/MP1 XI11_6/net20_4_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_11/MP0 XI11_6/net21_4_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_10/MP2 XI11_6/net20_5_ XI11_6/preck XI11_6/net21_5_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_10/MP1 XI11_6/net20_5_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_10/MP0 XI11_6/net21_5_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_9/MP2 XI11_6/net20_6_ XI11_6/preck XI11_6/net21_6_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_9/MP1 XI11_6/net20_6_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_9/MP0 XI11_6/net21_6_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_8/MP2 XI11_6/net20_7_ XI11_6/preck XI11_6/net21_7_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_8/MP1 XI11_6/net20_7_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_8/MP0 XI11_6/net21_7_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_7/MP2 XI11_6/net20_8_ XI11_6/preck XI11_6/net21_8_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_7/MP1 XI11_6/net20_8_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_7/MP0 XI11_6/net21_8_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_6/MP2 XI11_6/net20_9_ XI11_6/preck XI11_6/net21_9_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_6/MP1 XI11_6/net20_9_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_6/MP0 XI11_6/net21_9_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_5/MP2 XI11_6/net20_10_ XI11_6/preck XI11_6/net21_10_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_5/MP1 XI11_6/net20_10_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_5/MP0 XI11_6/net21_10_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_4/MP2 XI11_6/net20_11_ XI11_6/preck XI11_6/net21_11_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_4/MP1 XI11_6/net20_11_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_4/MP0 XI11_6/net21_11_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_3/MP2 XI11_6/net20_12_ XI11_6/preck XI11_6/net21_12_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_3/MP1 XI11_6/net20_12_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_3/MP0 XI11_6/net21_12_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_2/MP2 XI11_6/net20_13_ XI11_6/preck XI11_6/net21_13_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_2/MP1 XI11_6/net20_13_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_2/MP0 XI11_6/net21_13_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_1/MP2 XI11_6/net20_14_ XI11_6/preck XI11_6/net21_14_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_1/MP1 XI11_6/net20_14_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_1/MP0 XI11_6/net21_14_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_0/MP2 XI11_6/net20_15_ XI11_6/preck XI11_6/net21_15_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_6/XI1_0/MP1 XI11_6/net20_15_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI1_0/MP0 XI11_6/net21_15_ XI11_6/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_6/XI0/MN0_15 gnd gnd XI11_6/net21_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_14 gnd gnd XI11_6/net21_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_13 gnd gnd XI11_6/net21_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_12 gnd gnd XI11_6/net21_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_11 gnd gnd XI11_6/net21_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_10 gnd gnd XI11_6/net21_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_9 gnd gnd XI11_6/net21_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_8 gnd gnd XI11_6/net21_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_7 gnd gnd XI11_6/net21_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_6 gnd gnd XI11_6/net21_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_5 gnd gnd XI11_6/net21_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_4 gnd gnd XI11_6/net21_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_3 gnd gnd XI11_6/net21_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_2 gnd gnd XI11_6/net21_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_1 gnd gnd XI11_6/net21_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN0_0 gnd gnd XI11_6/net21_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_15 gnd gnd XI11_6/net20_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_14 gnd gnd XI11_6/net20_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_13 gnd gnd XI11_6/net20_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_12 gnd gnd XI11_6/net20_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_11 gnd gnd XI11_6/net20_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_10 gnd gnd XI11_6/net20_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_9 gnd gnd XI11_6/net20_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_8 gnd gnd XI11_6/net20_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_7 gnd gnd XI11_6/net20_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_6 gnd gnd XI11_6/net20_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_5 gnd gnd XI11_6/net20_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_4 gnd gnd XI11_6/net20_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_3 gnd gnd XI11_6/net20_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_2 gnd gnd XI11_6/net20_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_1 gnd gnd XI11_6/net20_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/MN1_0 gnd gnd XI11_6/net20_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_15 XI11_6/net21_0_ xsel_63_ XI11_6/XI0/XI0_63/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_14 XI11_6/net21_1_ xsel_63_ XI11_6/XI0/XI0_63/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_13 XI11_6/net21_2_ xsel_63_ XI11_6/XI0/XI0_63/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_12 XI11_6/net21_3_ xsel_63_ XI11_6/XI0/XI0_63/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_11 XI11_6/net21_4_ xsel_63_ XI11_6/XI0/XI0_63/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_10 XI11_6/net21_5_ xsel_63_ XI11_6/XI0/XI0_63/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_9 XI11_6/net21_6_ xsel_63_ XI11_6/XI0/XI0_63/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_8 XI11_6/net21_7_ xsel_63_ XI11_6/XI0/XI0_63/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_7 XI11_6/net21_8_ xsel_63_ XI11_6/XI0/XI0_63/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_6 XI11_6/net21_9_ xsel_63_ XI11_6/XI0/XI0_63/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_5 XI11_6/net21_10_ xsel_63_ XI11_6/XI0/XI0_63/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_4 XI11_6/net21_11_ xsel_63_ XI11_6/XI0/XI0_63/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_3 XI11_6/net21_12_ xsel_63_ XI11_6/XI0/XI0_63/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_2 XI11_6/net21_13_ xsel_63_ XI11_6/XI0/XI0_63/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_1 XI11_6/net21_14_ xsel_63_ XI11_6/XI0/XI0_63/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN0_0 XI11_6/net21_15_ xsel_63_ XI11_6/XI0/XI0_63/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_15 XI11_6/XI0/XI0_63/d__15_ xsel_63_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_14 XI11_6/XI0/XI0_63/d__14_ xsel_63_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_13 XI11_6/XI0/XI0_63/d__13_ xsel_63_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_12 XI11_6/XI0/XI0_63/d__12_ xsel_63_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_11 XI11_6/XI0/XI0_63/d__11_ xsel_63_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_10 XI11_6/XI0/XI0_63/d__10_ xsel_63_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_9 XI11_6/XI0/XI0_63/d__9_ xsel_63_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_8 XI11_6/XI0/XI0_63/d__8_ xsel_63_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_7 XI11_6/XI0/XI0_63/d__7_ xsel_63_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_6 XI11_6/XI0/XI0_63/d__6_ xsel_63_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_5 XI11_6/XI0/XI0_63/d__5_ xsel_63_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_4 XI11_6/XI0/XI0_63/d__4_ xsel_63_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_3 XI11_6/XI0/XI0_63/d__3_ xsel_63_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_2 XI11_6/XI0/XI0_63/d__2_ xsel_63_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_1 XI11_6/XI0/XI0_63/d__1_ xsel_63_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_63/MN1_0 XI11_6/XI0/XI0_63/d__0_ xsel_63_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_15 XI11_6/net21_0_ xsel_62_ XI11_6/XI0/XI0_62/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_14 XI11_6/net21_1_ xsel_62_ XI11_6/XI0/XI0_62/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_13 XI11_6/net21_2_ xsel_62_ XI11_6/XI0/XI0_62/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_12 XI11_6/net21_3_ xsel_62_ XI11_6/XI0/XI0_62/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_11 XI11_6/net21_4_ xsel_62_ XI11_6/XI0/XI0_62/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_10 XI11_6/net21_5_ xsel_62_ XI11_6/XI0/XI0_62/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_9 XI11_6/net21_6_ xsel_62_ XI11_6/XI0/XI0_62/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_8 XI11_6/net21_7_ xsel_62_ XI11_6/XI0/XI0_62/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_7 XI11_6/net21_8_ xsel_62_ XI11_6/XI0/XI0_62/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_6 XI11_6/net21_9_ xsel_62_ XI11_6/XI0/XI0_62/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_5 XI11_6/net21_10_ xsel_62_ XI11_6/XI0/XI0_62/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_4 XI11_6/net21_11_ xsel_62_ XI11_6/XI0/XI0_62/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_3 XI11_6/net21_12_ xsel_62_ XI11_6/XI0/XI0_62/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_2 XI11_6/net21_13_ xsel_62_ XI11_6/XI0/XI0_62/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_1 XI11_6/net21_14_ xsel_62_ XI11_6/XI0/XI0_62/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN0_0 XI11_6/net21_15_ xsel_62_ XI11_6/XI0/XI0_62/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_15 XI11_6/XI0/XI0_62/d__15_ xsel_62_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_14 XI11_6/XI0/XI0_62/d__14_ xsel_62_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_13 XI11_6/XI0/XI0_62/d__13_ xsel_62_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_12 XI11_6/XI0/XI0_62/d__12_ xsel_62_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_11 XI11_6/XI0/XI0_62/d__11_ xsel_62_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_10 XI11_6/XI0/XI0_62/d__10_ xsel_62_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_9 XI11_6/XI0/XI0_62/d__9_ xsel_62_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_8 XI11_6/XI0/XI0_62/d__8_ xsel_62_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_7 XI11_6/XI0/XI0_62/d__7_ xsel_62_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_6 XI11_6/XI0/XI0_62/d__6_ xsel_62_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_5 XI11_6/XI0/XI0_62/d__5_ xsel_62_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_4 XI11_6/XI0/XI0_62/d__4_ xsel_62_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_3 XI11_6/XI0/XI0_62/d__3_ xsel_62_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_2 XI11_6/XI0/XI0_62/d__2_ xsel_62_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_1 XI11_6/XI0/XI0_62/d__1_ xsel_62_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_62/MN1_0 XI11_6/XI0/XI0_62/d__0_ xsel_62_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_15 XI11_6/net21_0_ xsel_61_ XI11_6/XI0/XI0_61/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_14 XI11_6/net21_1_ xsel_61_ XI11_6/XI0/XI0_61/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_13 XI11_6/net21_2_ xsel_61_ XI11_6/XI0/XI0_61/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_12 XI11_6/net21_3_ xsel_61_ XI11_6/XI0/XI0_61/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_11 XI11_6/net21_4_ xsel_61_ XI11_6/XI0/XI0_61/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_10 XI11_6/net21_5_ xsel_61_ XI11_6/XI0/XI0_61/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_9 XI11_6/net21_6_ xsel_61_ XI11_6/XI0/XI0_61/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_8 XI11_6/net21_7_ xsel_61_ XI11_6/XI0/XI0_61/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_7 XI11_6/net21_8_ xsel_61_ XI11_6/XI0/XI0_61/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_6 XI11_6/net21_9_ xsel_61_ XI11_6/XI0/XI0_61/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_5 XI11_6/net21_10_ xsel_61_ XI11_6/XI0/XI0_61/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_4 XI11_6/net21_11_ xsel_61_ XI11_6/XI0/XI0_61/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_3 XI11_6/net21_12_ xsel_61_ XI11_6/XI0/XI0_61/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_2 XI11_6/net21_13_ xsel_61_ XI11_6/XI0/XI0_61/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_1 XI11_6/net21_14_ xsel_61_ XI11_6/XI0/XI0_61/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN0_0 XI11_6/net21_15_ xsel_61_ XI11_6/XI0/XI0_61/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_15 XI11_6/XI0/XI0_61/d__15_ xsel_61_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_14 XI11_6/XI0/XI0_61/d__14_ xsel_61_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_13 XI11_6/XI0/XI0_61/d__13_ xsel_61_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_12 XI11_6/XI0/XI0_61/d__12_ xsel_61_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_11 XI11_6/XI0/XI0_61/d__11_ xsel_61_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_10 XI11_6/XI0/XI0_61/d__10_ xsel_61_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_9 XI11_6/XI0/XI0_61/d__9_ xsel_61_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_8 XI11_6/XI0/XI0_61/d__8_ xsel_61_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_7 XI11_6/XI0/XI0_61/d__7_ xsel_61_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_6 XI11_6/XI0/XI0_61/d__6_ xsel_61_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_5 XI11_6/XI0/XI0_61/d__5_ xsel_61_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_4 XI11_6/XI0/XI0_61/d__4_ xsel_61_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_3 XI11_6/XI0/XI0_61/d__3_ xsel_61_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_2 XI11_6/XI0/XI0_61/d__2_ xsel_61_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_1 XI11_6/XI0/XI0_61/d__1_ xsel_61_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_61/MN1_0 XI11_6/XI0/XI0_61/d__0_ xsel_61_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_15 XI11_6/net21_0_ xsel_60_ XI11_6/XI0/XI0_60/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_14 XI11_6/net21_1_ xsel_60_ XI11_6/XI0/XI0_60/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_13 XI11_6/net21_2_ xsel_60_ XI11_6/XI0/XI0_60/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_12 XI11_6/net21_3_ xsel_60_ XI11_6/XI0/XI0_60/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_11 XI11_6/net21_4_ xsel_60_ XI11_6/XI0/XI0_60/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_10 XI11_6/net21_5_ xsel_60_ XI11_6/XI0/XI0_60/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_9 XI11_6/net21_6_ xsel_60_ XI11_6/XI0/XI0_60/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_8 XI11_6/net21_7_ xsel_60_ XI11_6/XI0/XI0_60/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_7 XI11_6/net21_8_ xsel_60_ XI11_6/XI0/XI0_60/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_6 XI11_6/net21_9_ xsel_60_ XI11_6/XI0/XI0_60/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_5 XI11_6/net21_10_ xsel_60_ XI11_6/XI0/XI0_60/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_4 XI11_6/net21_11_ xsel_60_ XI11_6/XI0/XI0_60/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_3 XI11_6/net21_12_ xsel_60_ XI11_6/XI0/XI0_60/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_2 XI11_6/net21_13_ xsel_60_ XI11_6/XI0/XI0_60/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_1 XI11_6/net21_14_ xsel_60_ XI11_6/XI0/XI0_60/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN0_0 XI11_6/net21_15_ xsel_60_ XI11_6/XI0/XI0_60/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_15 XI11_6/XI0/XI0_60/d__15_ xsel_60_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_14 XI11_6/XI0/XI0_60/d__14_ xsel_60_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_13 XI11_6/XI0/XI0_60/d__13_ xsel_60_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_12 XI11_6/XI0/XI0_60/d__12_ xsel_60_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_11 XI11_6/XI0/XI0_60/d__11_ xsel_60_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_10 XI11_6/XI0/XI0_60/d__10_ xsel_60_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_9 XI11_6/XI0/XI0_60/d__9_ xsel_60_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_8 XI11_6/XI0/XI0_60/d__8_ xsel_60_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_7 XI11_6/XI0/XI0_60/d__7_ xsel_60_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_6 XI11_6/XI0/XI0_60/d__6_ xsel_60_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_5 XI11_6/XI0/XI0_60/d__5_ xsel_60_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_4 XI11_6/XI0/XI0_60/d__4_ xsel_60_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_3 XI11_6/XI0/XI0_60/d__3_ xsel_60_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_2 XI11_6/XI0/XI0_60/d__2_ xsel_60_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_1 XI11_6/XI0/XI0_60/d__1_ xsel_60_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_60/MN1_0 XI11_6/XI0/XI0_60/d__0_ xsel_60_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_15 XI11_6/net21_0_ xsel_59_ XI11_6/XI0/XI0_59/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_14 XI11_6/net21_1_ xsel_59_ XI11_6/XI0/XI0_59/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_13 XI11_6/net21_2_ xsel_59_ XI11_6/XI0/XI0_59/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_12 XI11_6/net21_3_ xsel_59_ XI11_6/XI0/XI0_59/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_11 XI11_6/net21_4_ xsel_59_ XI11_6/XI0/XI0_59/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_10 XI11_6/net21_5_ xsel_59_ XI11_6/XI0/XI0_59/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_9 XI11_6/net21_6_ xsel_59_ XI11_6/XI0/XI0_59/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_8 XI11_6/net21_7_ xsel_59_ XI11_6/XI0/XI0_59/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_7 XI11_6/net21_8_ xsel_59_ XI11_6/XI0/XI0_59/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_6 XI11_6/net21_9_ xsel_59_ XI11_6/XI0/XI0_59/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_5 XI11_6/net21_10_ xsel_59_ XI11_6/XI0/XI0_59/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_4 XI11_6/net21_11_ xsel_59_ XI11_6/XI0/XI0_59/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_3 XI11_6/net21_12_ xsel_59_ XI11_6/XI0/XI0_59/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_2 XI11_6/net21_13_ xsel_59_ XI11_6/XI0/XI0_59/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_1 XI11_6/net21_14_ xsel_59_ XI11_6/XI0/XI0_59/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN0_0 XI11_6/net21_15_ xsel_59_ XI11_6/XI0/XI0_59/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_15 XI11_6/XI0/XI0_59/d__15_ xsel_59_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_14 XI11_6/XI0/XI0_59/d__14_ xsel_59_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_13 XI11_6/XI0/XI0_59/d__13_ xsel_59_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_12 XI11_6/XI0/XI0_59/d__12_ xsel_59_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_11 XI11_6/XI0/XI0_59/d__11_ xsel_59_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_10 XI11_6/XI0/XI0_59/d__10_ xsel_59_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_9 XI11_6/XI0/XI0_59/d__9_ xsel_59_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_8 XI11_6/XI0/XI0_59/d__8_ xsel_59_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_7 XI11_6/XI0/XI0_59/d__7_ xsel_59_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_6 XI11_6/XI0/XI0_59/d__6_ xsel_59_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_5 XI11_6/XI0/XI0_59/d__5_ xsel_59_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_4 XI11_6/XI0/XI0_59/d__4_ xsel_59_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_3 XI11_6/XI0/XI0_59/d__3_ xsel_59_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_2 XI11_6/XI0/XI0_59/d__2_ xsel_59_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_1 XI11_6/XI0/XI0_59/d__1_ xsel_59_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_59/MN1_0 XI11_6/XI0/XI0_59/d__0_ xsel_59_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_15 XI11_6/net21_0_ xsel_58_ XI11_6/XI0/XI0_58/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_14 XI11_6/net21_1_ xsel_58_ XI11_6/XI0/XI0_58/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_13 XI11_6/net21_2_ xsel_58_ XI11_6/XI0/XI0_58/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_12 XI11_6/net21_3_ xsel_58_ XI11_6/XI0/XI0_58/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_11 XI11_6/net21_4_ xsel_58_ XI11_6/XI0/XI0_58/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_10 XI11_6/net21_5_ xsel_58_ XI11_6/XI0/XI0_58/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_9 XI11_6/net21_6_ xsel_58_ XI11_6/XI0/XI0_58/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_8 XI11_6/net21_7_ xsel_58_ XI11_6/XI0/XI0_58/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_7 XI11_6/net21_8_ xsel_58_ XI11_6/XI0/XI0_58/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_6 XI11_6/net21_9_ xsel_58_ XI11_6/XI0/XI0_58/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_5 XI11_6/net21_10_ xsel_58_ XI11_6/XI0/XI0_58/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_4 XI11_6/net21_11_ xsel_58_ XI11_6/XI0/XI0_58/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_3 XI11_6/net21_12_ xsel_58_ XI11_6/XI0/XI0_58/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_2 XI11_6/net21_13_ xsel_58_ XI11_6/XI0/XI0_58/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_1 XI11_6/net21_14_ xsel_58_ XI11_6/XI0/XI0_58/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN0_0 XI11_6/net21_15_ xsel_58_ XI11_6/XI0/XI0_58/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_15 XI11_6/XI0/XI0_58/d__15_ xsel_58_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_14 XI11_6/XI0/XI0_58/d__14_ xsel_58_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_13 XI11_6/XI0/XI0_58/d__13_ xsel_58_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_12 XI11_6/XI0/XI0_58/d__12_ xsel_58_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_11 XI11_6/XI0/XI0_58/d__11_ xsel_58_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_10 XI11_6/XI0/XI0_58/d__10_ xsel_58_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_9 XI11_6/XI0/XI0_58/d__9_ xsel_58_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_8 XI11_6/XI0/XI0_58/d__8_ xsel_58_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_7 XI11_6/XI0/XI0_58/d__7_ xsel_58_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_6 XI11_6/XI0/XI0_58/d__6_ xsel_58_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_5 XI11_6/XI0/XI0_58/d__5_ xsel_58_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_4 XI11_6/XI0/XI0_58/d__4_ xsel_58_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_3 XI11_6/XI0/XI0_58/d__3_ xsel_58_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_2 XI11_6/XI0/XI0_58/d__2_ xsel_58_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_1 XI11_6/XI0/XI0_58/d__1_ xsel_58_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_58/MN1_0 XI11_6/XI0/XI0_58/d__0_ xsel_58_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_15 XI11_6/net21_0_ xsel_57_ XI11_6/XI0/XI0_57/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_14 XI11_6/net21_1_ xsel_57_ XI11_6/XI0/XI0_57/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_13 XI11_6/net21_2_ xsel_57_ XI11_6/XI0/XI0_57/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_12 XI11_6/net21_3_ xsel_57_ XI11_6/XI0/XI0_57/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_11 XI11_6/net21_4_ xsel_57_ XI11_6/XI0/XI0_57/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_10 XI11_6/net21_5_ xsel_57_ XI11_6/XI0/XI0_57/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_9 XI11_6/net21_6_ xsel_57_ XI11_6/XI0/XI0_57/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_8 XI11_6/net21_7_ xsel_57_ XI11_6/XI0/XI0_57/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_7 XI11_6/net21_8_ xsel_57_ XI11_6/XI0/XI0_57/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_6 XI11_6/net21_9_ xsel_57_ XI11_6/XI0/XI0_57/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_5 XI11_6/net21_10_ xsel_57_ XI11_6/XI0/XI0_57/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_4 XI11_6/net21_11_ xsel_57_ XI11_6/XI0/XI0_57/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_3 XI11_6/net21_12_ xsel_57_ XI11_6/XI0/XI0_57/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_2 XI11_6/net21_13_ xsel_57_ XI11_6/XI0/XI0_57/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_1 XI11_6/net21_14_ xsel_57_ XI11_6/XI0/XI0_57/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN0_0 XI11_6/net21_15_ xsel_57_ XI11_6/XI0/XI0_57/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_15 XI11_6/XI0/XI0_57/d__15_ xsel_57_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_14 XI11_6/XI0/XI0_57/d__14_ xsel_57_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_13 XI11_6/XI0/XI0_57/d__13_ xsel_57_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_12 XI11_6/XI0/XI0_57/d__12_ xsel_57_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_11 XI11_6/XI0/XI0_57/d__11_ xsel_57_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_10 XI11_6/XI0/XI0_57/d__10_ xsel_57_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_9 XI11_6/XI0/XI0_57/d__9_ xsel_57_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_8 XI11_6/XI0/XI0_57/d__8_ xsel_57_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_7 XI11_6/XI0/XI0_57/d__7_ xsel_57_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_6 XI11_6/XI0/XI0_57/d__6_ xsel_57_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_5 XI11_6/XI0/XI0_57/d__5_ xsel_57_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_4 XI11_6/XI0/XI0_57/d__4_ xsel_57_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_3 XI11_6/XI0/XI0_57/d__3_ xsel_57_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_2 XI11_6/XI0/XI0_57/d__2_ xsel_57_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_1 XI11_6/XI0/XI0_57/d__1_ xsel_57_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_57/MN1_0 XI11_6/XI0/XI0_57/d__0_ xsel_57_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_15 XI11_6/net21_0_ xsel_56_ XI11_6/XI0/XI0_56/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_14 XI11_6/net21_1_ xsel_56_ XI11_6/XI0/XI0_56/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_13 XI11_6/net21_2_ xsel_56_ XI11_6/XI0/XI0_56/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_12 XI11_6/net21_3_ xsel_56_ XI11_6/XI0/XI0_56/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_11 XI11_6/net21_4_ xsel_56_ XI11_6/XI0/XI0_56/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_10 XI11_6/net21_5_ xsel_56_ XI11_6/XI0/XI0_56/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_9 XI11_6/net21_6_ xsel_56_ XI11_6/XI0/XI0_56/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_8 XI11_6/net21_7_ xsel_56_ XI11_6/XI0/XI0_56/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_7 XI11_6/net21_8_ xsel_56_ XI11_6/XI0/XI0_56/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_6 XI11_6/net21_9_ xsel_56_ XI11_6/XI0/XI0_56/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_5 XI11_6/net21_10_ xsel_56_ XI11_6/XI0/XI0_56/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_4 XI11_6/net21_11_ xsel_56_ XI11_6/XI0/XI0_56/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_3 XI11_6/net21_12_ xsel_56_ XI11_6/XI0/XI0_56/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_2 XI11_6/net21_13_ xsel_56_ XI11_6/XI0/XI0_56/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_1 XI11_6/net21_14_ xsel_56_ XI11_6/XI0/XI0_56/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN0_0 XI11_6/net21_15_ xsel_56_ XI11_6/XI0/XI0_56/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_15 XI11_6/XI0/XI0_56/d__15_ xsel_56_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_14 XI11_6/XI0/XI0_56/d__14_ xsel_56_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_13 XI11_6/XI0/XI0_56/d__13_ xsel_56_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_12 XI11_6/XI0/XI0_56/d__12_ xsel_56_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_11 XI11_6/XI0/XI0_56/d__11_ xsel_56_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_10 XI11_6/XI0/XI0_56/d__10_ xsel_56_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_9 XI11_6/XI0/XI0_56/d__9_ xsel_56_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_8 XI11_6/XI0/XI0_56/d__8_ xsel_56_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_7 XI11_6/XI0/XI0_56/d__7_ xsel_56_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_6 XI11_6/XI0/XI0_56/d__6_ xsel_56_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_5 XI11_6/XI0/XI0_56/d__5_ xsel_56_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_4 XI11_6/XI0/XI0_56/d__4_ xsel_56_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_3 XI11_6/XI0/XI0_56/d__3_ xsel_56_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_2 XI11_6/XI0/XI0_56/d__2_ xsel_56_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_1 XI11_6/XI0/XI0_56/d__1_ xsel_56_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_56/MN1_0 XI11_6/XI0/XI0_56/d__0_ xsel_56_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_15 XI11_6/net21_0_ xsel_55_ XI11_6/XI0/XI0_55/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_14 XI11_6/net21_1_ xsel_55_ XI11_6/XI0/XI0_55/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_13 XI11_6/net21_2_ xsel_55_ XI11_6/XI0/XI0_55/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_12 XI11_6/net21_3_ xsel_55_ XI11_6/XI0/XI0_55/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_11 XI11_6/net21_4_ xsel_55_ XI11_6/XI0/XI0_55/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_10 XI11_6/net21_5_ xsel_55_ XI11_6/XI0/XI0_55/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_9 XI11_6/net21_6_ xsel_55_ XI11_6/XI0/XI0_55/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_8 XI11_6/net21_7_ xsel_55_ XI11_6/XI0/XI0_55/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_7 XI11_6/net21_8_ xsel_55_ XI11_6/XI0/XI0_55/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_6 XI11_6/net21_9_ xsel_55_ XI11_6/XI0/XI0_55/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_5 XI11_6/net21_10_ xsel_55_ XI11_6/XI0/XI0_55/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_4 XI11_6/net21_11_ xsel_55_ XI11_6/XI0/XI0_55/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_3 XI11_6/net21_12_ xsel_55_ XI11_6/XI0/XI0_55/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_2 XI11_6/net21_13_ xsel_55_ XI11_6/XI0/XI0_55/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_1 XI11_6/net21_14_ xsel_55_ XI11_6/XI0/XI0_55/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN0_0 XI11_6/net21_15_ xsel_55_ XI11_6/XI0/XI0_55/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_15 XI11_6/XI0/XI0_55/d__15_ xsel_55_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_14 XI11_6/XI0/XI0_55/d__14_ xsel_55_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_13 XI11_6/XI0/XI0_55/d__13_ xsel_55_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_12 XI11_6/XI0/XI0_55/d__12_ xsel_55_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_11 XI11_6/XI0/XI0_55/d__11_ xsel_55_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_10 XI11_6/XI0/XI0_55/d__10_ xsel_55_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_9 XI11_6/XI0/XI0_55/d__9_ xsel_55_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_8 XI11_6/XI0/XI0_55/d__8_ xsel_55_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_7 XI11_6/XI0/XI0_55/d__7_ xsel_55_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_6 XI11_6/XI0/XI0_55/d__6_ xsel_55_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_5 XI11_6/XI0/XI0_55/d__5_ xsel_55_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_4 XI11_6/XI0/XI0_55/d__4_ xsel_55_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_3 XI11_6/XI0/XI0_55/d__3_ xsel_55_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_2 XI11_6/XI0/XI0_55/d__2_ xsel_55_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_1 XI11_6/XI0/XI0_55/d__1_ xsel_55_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_55/MN1_0 XI11_6/XI0/XI0_55/d__0_ xsel_55_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_15 XI11_6/net21_0_ xsel_54_ XI11_6/XI0/XI0_54/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_14 XI11_6/net21_1_ xsel_54_ XI11_6/XI0/XI0_54/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_13 XI11_6/net21_2_ xsel_54_ XI11_6/XI0/XI0_54/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_12 XI11_6/net21_3_ xsel_54_ XI11_6/XI0/XI0_54/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_11 XI11_6/net21_4_ xsel_54_ XI11_6/XI0/XI0_54/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_10 XI11_6/net21_5_ xsel_54_ XI11_6/XI0/XI0_54/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_9 XI11_6/net21_6_ xsel_54_ XI11_6/XI0/XI0_54/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_8 XI11_6/net21_7_ xsel_54_ XI11_6/XI0/XI0_54/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_7 XI11_6/net21_8_ xsel_54_ XI11_6/XI0/XI0_54/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_6 XI11_6/net21_9_ xsel_54_ XI11_6/XI0/XI0_54/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_5 XI11_6/net21_10_ xsel_54_ XI11_6/XI0/XI0_54/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_4 XI11_6/net21_11_ xsel_54_ XI11_6/XI0/XI0_54/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_3 XI11_6/net21_12_ xsel_54_ XI11_6/XI0/XI0_54/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_2 XI11_6/net21_13_ xsel_54_ XI11_6/XI0/XI0_54/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_1 XI11_6/net21_14_ xsel_54_ XI11_6/XI0/XI0_54/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN0_0 XI11_6/net21_15_ xsel_54_ XI11_6/XI0/XI0_54/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_15 XI11_6/XI0/XI0_54/d__15_ xsel_54_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_14 XI11_6/XI0/XI0_54/d__14_ xsel_54_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_13 XI11_6/XI0/XI0_54/d__13_ xsel_54_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_12 XI11_6/XI0/XI0_54/d__12_ xsel_54_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_11 XI11_6/XI0/XI0_54/d__11_ xsel_54_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_10 XI11_6/XI0/XI0_54/d__10_ xsel_54_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_9 XI11_6/XI0/XI0_54/d__9_ xsel_54_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_8 XI11_6/XI0/XI0_54/d__8_ xsel_54_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_7 XI11_6/XI0/XI0_54/d__7_ xsel_54_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_6 XI11_6/XI0/XI0_54/d__6_ xsel_54_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_5 XI11_6/XI0/XI0_54/d__5_ xsel_54_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_4 XI11_6/XI0/XI0_54/d__4_ xsel_54_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_3 XI11_6/XI0/XI0_54/d__3_ xsel_54_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_2 XI11_6/XI0/XI0_54/d__2_ xsel_54_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_1 XI11_6/XI0/XI0_54/d__1_ xsel_54_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_54/MN1_0 XI11_6/XI0/XI0_54/d__0_ xsel_54_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_15 XI11_6/net21_0_ xsel_53_ XI11_6/XI0/XI0_53/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_14 XI11_6/net21_1_ xsel_53_ XI11_6/XI0/XI0_53/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_13 XI11_6/net21_2_ xsel_53_ XI11_6/XI0/XI0_53/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_12 XI11_6/net21_3_ xsel_53_ XI11_6/XI0/XI0_53/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_11 XI11_6/net21_4_ xsel_53_ XI11_6/XI0/XI0_53/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_10 XI11_6/net21_5_ xsel_53_ XI11_6/XI0/XI0_53/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_9 XI11_6/net21_6_ xsel_53_ XI11_6/XI0/XI0_53/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_8 XI11_6/net21_7_ xsel_53_ XI11_6/XI0/XI0_53/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_7 XI11_6/net21_8_ xsel_53_ XI11_6/XI0/XI0_53/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_6 XI11_6/net21_9_ xsel_53_ XI11_6/XI0/XI0_53/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_5 XI11_6/net21_10_ xsel_53_ XI11_6/XI0/XI0_53/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_4 XI11_6/net21_11_ xsel_53_ XI11_6/XI0/XI0_53/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_3 XI11_6/net21_12_ xsel_53_ XI11_6/XI0/XI0_53/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_2 XI11_6/net21_13_ xsel_53_ XI11_6/XI0/XI0_53/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_1 XI11_6/net21_14_ xsel_53_ XI11_6/XI0/XI0_53/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN0_0 XI11_6/net21_15_ xsel_53_ XI11_6/XI0/XI0_53/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_15 XI11_6/XI0/XI0_53/d__15_ xsel_53_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_14 XI11_6/XI0/XI0_53/d__14_ xsel_53_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_13 XI11_6/XI0/XI0_53/d__13_ xsel_53_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_12 XI11_6/XI0/XI0_53/d__12_ xsel_53_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_11 XI11_6/XI0/XI0_53/d__11_ xsel_53_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_10 XI11_6/XI0/XI0_53/d__10_ xsel_53_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_9 XI11_6/XI0/XI0_53/d__9_ xsel_53_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_8 XI11_6/XI0/XI0_53/d__8_ xsel_53_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_7 XI11_6/XI0/XI0_53/d__7_ xsel_53_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_6 XI11_6/XI0/XI0_53/d__6_ xsel_53_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_5 XI11_6/XI0/XI0_53/d__5_ xsel_53_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_4 XI11_6/XI0/XI0_53/d__4_ xsel_53_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_3 XI11_6/XI0/XI0_53/d__3_ xsel_53_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_2 XI11_6/XI0/XI0_53/d__2_ xsel_53_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_1 XI11_6/XI0/XI0_53/d__1_ xsel_53_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_53/MN1_0 XI11_6/XI0/XI0_53/d__0_ xsel_53_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_15 XI11_6/net21_0_ xsel_52_ XI11_6/XI0/XI0_52/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_14 XI11_6/net21_1_ xsel_52_ XI11_6/XI0/XI0_52/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_13 XI11_6/net21_2_ xsel_52_ XI11_6/XI0/XI0_52/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_12 XI11_6/net21_3_ xsel_52_ XI11_6/XI0/XI0_52/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_11 XI11_6/net21_4_ xsel_52_ XI11_6/XI0/XI0_52/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_10 XI11_6/net21_5_ xsel_52_ XI11_6/XI0/XI0_52/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_9 XI11_6/net21_6_ xsel_52_ XI11_6/XI0/XI0_52/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_8 XI11_6/net21_7_ xsel_52_ XI11_6/XI0/XI0_52/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_7 XI11_6/net21_8_ xsel_52_ XI11_6/XI0/XI0_52/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_6 XI11_6/net21_9_ xsel_52_ XI11_6/XI0/XI0_52/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_5 XI11_6/net21_10_ xsel_52_ XI11_6/XI0/XI0_52/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_4 XI11_6/net21_11_ xsel_52_ XI11_6/XI0/XI0_52/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_3 XI11_6/net21_12_ xsel_52_ XI11_6/XI0/XI0_52/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_2 XI11_6/net21_13_ xsel_52_ XI11_6/XI0/XI0_52/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_1 XI11_6/net21_14_ xsel_52_ XI11_6/XI0/XI0_52/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN0_0 XI11_6/net21_15_ xsel_52_ XI11_6/XI0/XI0_52/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_15 XI11_6/XI0/XI0_52/d__15_ xsel_52_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_14 XI11_6/XI0/XI0_52/d__14_ xsel_52_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_13 XI11_6/XI0/XI0_52/d__13_ xsel_52_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_12 XI11_6/XI0/XI0_52/d__12_ xsel_52_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_11 XI11_6/XI0/XI0_52/d__11_ xsel_52_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_10 XI11_6/XI0/XI0_52/d__10_ xsel_52_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_9 XI11_6/XI0/XI0_52/d__9_ xsel_52_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_8 XI11_6/XI0/XI0_52/d__8_ xsel_52_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_7 XI11_6/XI0/XI0_52/d__7_ xsel_52_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_6 XI11_6/XI0/XI0_52/d__6_ xsel_52_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_5 XI11_6/XI0/XI0_52/d__5_ xsel_52_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_4 XI11_6/XI0/XI0_52/d__4_ xsel_52_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_3 XI11_6/XI0/XI0_52/d__3_ xsel_52_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_2 XI11_6/XI0/XI0_52/d__2_ xsel_52_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_1 XI11_6/XI0/XI0_52/d__1_ xsel_52_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_52/MN1_0 XI11_6/XI0/XI0_52/d__0_ xsel_52_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_15 XI11_6/net21_0_ xsel_51_ XI11_6/XI0/XI0_51/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_14 XI11_6/net21_1_ xsel_51_ XI11_6/XI0/XI0_51/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_13 XI11_6/net21_2_ xsel_51_ XI11_6/XI0/XI0_51/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_12 XI11_6/net21_3_ xsel_51_ XI11_6/XI0/XI0_51/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_11 XI11_6/net21_4_ xsel_51_ XI11_6/XI0/XI0_51/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_10 XI11_6/net21_5_ xsel_51_ XI11_6/XI0/XI0_51/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_9 XI11_6/net21_6_ xsel_51_ XI11_6/XI0/XI0_51/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_8 XI11_6/net21_7_ xsel_51_ XI11_6/XI0/XI0_51/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_7 XI11_6/net21_8_ xsel_51_ XI11_6/XI0/XI0_51/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_6 XI11_6/net21_9_ xsel_51_ XI11_6/XI0/XI0_51/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_5 XI11_6/net21_10_ xsel_51_ XI11_6/XI0/XI0_51/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_4 XI11_6/net21_11_ xsel_51_ XI11_6/XI0/XI0_51/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_3 XI11_6/net21_12_ xsel_51_ XI11_6/XI0/XI0_51/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_2 XI11_6/net21_13_ xsel_51_ XI11_6/XI0/XI0_51/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_1 XI11_6/net21_14_ xsel_51_ XI11_6/XI0/XI0_51/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN0_0 XI11_6/net21_15_ xsel_51_ XI11_6/XI0/XI0_51/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_15 XI11_6/XI0/XI0_51/d__15_ xsel_51_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_14 XI11_6/XI0/XI0_51/d__14_ xsel_51_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_13 XI11_6/XI0/XI0_51/d__13_ xsel_51_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_12 XI11_6/XI0/XI0_51/d__12_ xsel_51_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_11 XI11_6/XI0/XI0_51/d__11_ xsel_51_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_10 XI11_6/XI0/XI0_51/d__10_ xsel_51_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_9 XI11_6/XI0/XI0_51/d__9_ xsel_51_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_8 XI11_6/XI0/XI0_51/d__8_ xsel_51_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_7 XI11_6/XI0/XI0_51/d__7_ xsel_51_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_6 XI11_6/XI0/XI0_51/d__6_ xsel_51_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_5 XI11_6/XI0/XI0_51/d__5_ xsel_51_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_4 XI11_6/XI0/XI0_51/d__4_ xsel_51_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_3 XI11_6/XI0/XI0_51/d__3_ xsel_51_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_2 XI11_6/XI0/XI0_51/d__2_ xsel_51_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_1 XI11_6/XI0/XI0_51/d__1_ xsel_51_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_51/MN1_0 XI11_6/XI0/XI0_51/d__0_ xsel_51_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_15 XI11_6/net21_0_ xsel_50_ XI11_6/XI0/XI0_50/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_14 XI11_6/net21_1_ xsel_50_ XI11_6/XI0/XI0_50/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_13 XI11_6/net21_2_ xsel_50_ XI11_6/XI0/XI0_50/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_12 XI11_6/net21_3_ xsel_50_ XI11_6/XI0/XI0_50/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_11 XI11_6/net21_4_ xsel_50_ XI11_6/XI0/XI0_50/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_10 XI11_6/net21_5_ xsel_50_ XI11_6/XI0/XI0_50/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_9 XI11_6/net21_6_ xsel_50_ XI11_6/XI0/XI0_50/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_8 XI11_6/net21_7_ xsel_50_ XI11_6/XI0/XI0_50/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_7 XI11_6/net21_8_ xsel_50_ XI11_6/XI0/XI0_50/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_6 XI11_6/net21_9_ xsel_50_ XI11_6/XI0/XI0_50/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_5 XI11_6/net21_10_ xsel_50_ XI11_6/XI0/XI0_50/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_4 XI11_6/net21_11_ xsel_50_ XI11_6/XI0/XI0_50/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_3 XI11_6/net21_12_ xsel_50_ XI11_6/XI0/XI0_50/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_2 XI11_6/net21_13_ xsel_50_ XI11_6/XI0/XI0_50/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_1 XI11_6/net21_14_ xsel_50_ XI11_6/XI0/XI0_50/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN0_0 XI11_6/net21_15_ xsel_50_ XI11_6/XI0/XI0_50/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_15 XI11_6/XI0/XI0_50/d__15_ xsel_50_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_14 XI11_6/XI0/XI0_50/d__14_ xsel_50_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_13 XI11_6/XI0/XI0_50/d__13_ xsel_50_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_12 XI11_6/XI0/XI0_50/d__12_ xsel_50_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_11 XI11_6/XI0/XI0_50/d__11_ xsel_50_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_10 XI11_6/XI0/XI0_50/d__10_ xsel_50_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_9 XI11_6/XI0/XI0_50/d__9_ xsel_50_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_8 XI11_6/XI0/XI0_50/d__8_ xsel_50_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_7 XI11_6/XI0/XI0_50/d__7_ xsel_50_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_6 XI11_6/XI0/XI0_50/d__6_ xsel_50_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_5 XI11_6/XI0/XI0_50/d__5_ xsel_50_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_4 XI11_6/XI0/XI0_50/d__4_ xsel_50_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_3 XI11_6/XI0/XI0_50/d__3_ xsel_50_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_2 XI11_6/XI0/XI0_50/d__2_ xsel_50_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_1 XI11_6/XI0/XI0_50/d__1_ xsel_50_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_50/MN1_0 XI11_6/XI0/XI0_50/d__0_ xsel_50_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_15 XI11_6/net21_0_ xsel_49_ XI11_6/XI0/XI0_49/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_14 XI11_6/net21_1_ xsel_49_ XI11_6/XI0/XI0_49/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_13 XI11_6/net21_2_ xsel_49_ XI11_6/XI0/XI0_49/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_12 XI11_6/net21_3_ xsel_49_ XI11_6/XI0/XI0_49/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_11 XI11_6/net21_4_ xsel_49_ XI11_6/XI0/XI0_49/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_10 XI11_6/net21_5_ xsel_49_ XI11_6/XI0/XI0_49/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_9 XI11_6/net21_6_ xsel_49_ XI11_6/XI0/XI0_49/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_8 XI11_6/net21_7_ xsel_49_ XI11_6/XI0/XI0_49/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_7 XI11_6/net21_8_ xsel_49_ XI11_6/XI0/XI0_49/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_6 XI11_6/net21_9_ xsel_49_ XI11_6/XI0/XI0_49/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_5 XI11_6/net21_10_ xsel_49_ XI11_6/XI0/XI0_49/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_4 XI11_6/net21_11_ xsel_49_ XI11_6/XI0/XI0_49/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_3 XI11_6/net21_12_ xsel_49_ XI11_6/XI0/XI0_49/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_2 XI11_6/net21_13_ xsel_49_ XI11_6/XI0/XI0_49/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_1 XI11_6/net21_14_ xsel_49_ XI11_6/XI0/XI0_49/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN0_0 XI11_6/net21_15_ xsel_49_ XI11_6/XI0/XI0_49/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_15 XI11_6/XI0/XI0_49/d__15_ xsel_49_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_14 XI11_6/XI0/XI0_49/d__14_ xsel_49_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_13 XI11_6/XI0/XI0_49/d__13_ xsel_49_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_12 XI11_6/XI0/XI0_49/d__12_ xsel_49_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_11 XI11_6/XI0/XI0_49/d__11_ xsel_49_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_10 XI11_6/XI0/XI0_49/d__10_ xsel_49_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_9 XI11_6/XI0/XI0_49/d__9_ xsel_49_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_8 XI11_6/XI0/XI0_49/d__8_ xsel_49_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_7 XI11_6/XI0/XI0_49/d__7_ xsel_49_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_6 XI11_6/XI0/XI0_49/d__6_ xsel_49_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_5 XI11_6/XI0/XI0_49/d__5_ xsel_49_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_4 XI11_6/XI0/XI0_49/d__4_ xsel_49_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_3 XI11_6/XI0/XI0_49/d__3_ xsel_49_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_2 XI11_6/XI0/XI0_49/d__2_ xsel_49_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_1 XI11_6/XI0/XI0_49/d__1_ xsel_49_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_49/MN1_0 XI11_6/XI0/XI0_49/d__0_ xsel_49_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_15 XI11_6/net21_0_ xsel_48_ XI11_6/XI0/XI0_48/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_14 XI11_6/net21_1_ xsel_48_ XI11_6/XI0/XI0_48/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_13 XI11_6/net21_2_ xsel_48_ XI11_6/XI0/XI0_48/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_12 XI11_6/net21_3_ xsel_48_ XI11_6/XI0/XI0_48/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_11 XI11_6/net21_4_ xsel_48_ XI11_6/XI0/XI0_48/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_10 XI11_6/net21_5_ xsel_48_ XI11_6/XI0/XI0_48/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_9 XI11_6/net21_6_ xsel_48_ XI11_6/XI0/XI0_48/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_8 XI11_6/net21_7_ xsel_48_ XI11_6/XI0/XI0_48/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_7 XI11_6/net21_8_ xsel_48_ XI11_6/XI0/XI0_48/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_6 XI11_6/net21_9_ xsel_48_ XI11_6/XI0/XI0_48/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_5 XI11_6/net21_10_ xsel_48_ XI11_6/XI0/XI0_48/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_4 XI11_6/net21_11_ xsel_48_ XI11_6/XI0/XI0_48/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_3 XI11_6/net21_12_ xsel_48_ XI11_6/XI0/XI0_48/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_2 XI11_6/net21_13_ xsel_48_ XI11_6/XI0/XI0_48/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_1 XI11_6/net21_14_ xsel_48_ XI11_6/XI0/XI0_48/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN0_0 XI11_6/net21_15_ xsel_48_ XI11_6/XI0/XI0_48/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_15 XI11_6/XI0/XI0_48/d__15_ xsel_48_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_14 XI11_6/XI0/XI0_48/d__14_ xsel_48_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_13 XI11_6/XI0/XI0_48/d__13_ xsel_48_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_12 XI11_6/XI0/XI0_48/d__12_ xsel_48_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_11 XI11_6/XI0/XI0_48/d__11_ xsel_48_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_10 XI11_6/XI0/XI0_48/d__10_ xsel_48_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_9 XI11_6/XI0/XI0_48/d__9_ xsel_48_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_8 XI11_6/XI0/XI0_48/d__8_ xsel_48_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_7 XI11_6/XI0/XI0_48/d__7_ xsel_48_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_6 XI11_6/XI0/XI0_48/d__6_ xsel_48_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_5 XI11_6/XI0/XI0_48/d__5_ xsel_48_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_4 XI11_6/XI0/XI0_48/d__4_ xsel_48_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_3 XI11_6/XI0/XI0_48/d__3_ xsel_48_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_2 XI11_6/XI0/XI0_48/d__2_ xsel_48_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_1 XI11_6/XI0/XI0_48/d__1_ xsel_48_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_48/MN1_0 XI11_6/XI0/XI0_48/d__0_ xsel_48_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_15 XI11_6/net21_0_ xsel_47_ XI11_6/XI0/XI0_47/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_14 XI11_6/net21_1_ xsel_47_ XI11_6/XI0/XI0_47/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_13 XI11_6/net21_2_ xsel_47_ XI11_6/XI0/XI0_47/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_12 XI11_6/net21_3_ xsel_47_ XI11_6/XI0/XI0_47/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_11 XI11_6/net21_4_ xsel_47_ XI11_6/XI0/XI0_47/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_10 XI11_6/net21_5_ xsel_47_ XI11_6/XI0/XI0_47/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_9 XI11_6/net21_6_ xsel_47_ XI11_6/XI0/XI0_47/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_8 XI11_6/net21_7_ xsel_47_ XI11_6/XI0/XI0_47/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_7 XI11_6/net21_8_ xsel_47_ XI11_6/XI0/XI0_47/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_6 XI11_6/net21_9_ xsel_47_ XI11_6/XI0/XI0_47/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_5 XI11_6/net21_10_ xsel_47_ XI11_6/XI0/XI0_47/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_4 XI11_6/net21_11_ xsel_47_ XI11_6/XI0/XI0_47/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_3 XI11_6/net21_12_ xsel_47_ XI11_6/XI0/XI0_47/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_2 XI11_6/net21_13_ xsel_47_ XI11_6/XI0/XI0_47/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_1 XI11_6/net21_14_ xsel_47_ XI11_6/XI0/XI0_47/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN0_0 XI11_6/net21_15_ xsel_47_ XI11_6/XI0/XI0_47/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_15 XI11_6/XI0/XI0_47/d__15_ xsel_47_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_14 XI11_6/XI0/XI0_47/d__14_ xsel_47_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_13 XI11_6/XI0/XI0_47/d__13_ xsel_47_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_12 XI11_6/XI0/XI0_47/d__12_ xsel_47_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_11 XI11_6/XI0/XI0_47/d__11_ xsel_47_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_10 XI11_6/XI0/XI0_47/d__10_ xsel_47_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_9 XI11_6/XI0/XI0_47/d__9_ xsel_47_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_8 XI11_6/XI0/XI0_47/d__8_ xsel_47_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_7 XI11_6/XI0/XI0_47/d__7_ xsel_47_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_6 XI11_6/XI0/XI0_47/d__6_ xsel_47_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_5 XI11_6/XI0/XI0_47/d__5_ xsel_47_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_4 XI11_6/XI0/XI0_47/d__4_ xsel_47_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_3 XI11_6/XI0/XI0_47/d__3_ xsel_47_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_2 XI11_6/XI0/XI0_47/d__2_ xsel_47_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_1 XI11_6/XI0/XI0_47/d__1_ xsel_47_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_47/MN1_0 XI11_6/XI0/XI0_47/d__0_ xsel_47_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_15 XI11_6/net21_0_ xsel_46_ XI11_6/XI0/XI0_46/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_14 XI11_6/net21_1_ xsel_46_ XI11_6/XI0/XI0_46/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_13 XI11_6/net21_2_ xsel_46_ XI11_6/XI0/XI0_46/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_12 XI11_6/net21_3_ xsel_46_ XI11_6/XI0/XI0_46/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_11 XI11_6/net21_4_ xsel_46_ XI11_6/XI0/XI0_46/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_10 XI11_6/net21_5_ xsel_46_ XI11_6/XI0/XI0_46/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_9 XI11_6/net21_6_ xsel_46_ XI11_6/XI0/XI0_46/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_8 XI11_6/net21_7_ xsel_46_ XI11_6/XI0/XI0_46/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_7 XI11_6/net21_8_ xsel_46_ XI11_6/XI0/XI0_46/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_6 XI11_6/net21_9_ xsel_46_ XI11_6/XI0/XI0_46/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_5 XI11_6/net21_10_ xsel_46_ XI11_6/XI0/XI0_46/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_4 XI11_6/net21_11_ xsel_46_ XI11_6/XI0/XI0_46/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_3 XI11_6/net21_12_ xsel_46_ XI11_6/XI0/XI0_46/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_2 XI11_6/net21_13_ xsel_46_ XI11_6/XI0/XI0_46/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_1 XI11_6/net21_14_ xsel_46_ XI11_6/XI0/XI0_46/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN0_0 XI11_6/net21_15_ xsel_46_ XI11_6/XI0/XI0_46/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_15 XI11_6/XI0/XI0_46/d__15_ xsel_46_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_14 XI11_6/XI0/XI0_46/d__14_ xsel_46_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_13 XI11_6/XI0/XI0_46/d__13_ xsel_46_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_12 XI11_6/XI0/XI0_46/d__12_ xsel_46_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_11 XI11_6/XI0/XI0_46/d__11_ xsel_46_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_10 XI11_6/XI0/XI0_46/d__10_ xsel_46_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_9 XI11_6/XI0/XI0_46/d__9_ xsel_46_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_8 XI11_6/XI0/XI0_46/d__8_ xsel_46_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_7 XI11_6/XI0/XI0_46/d__7_ xsel_46_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_6 XI11_6/XI0/XI0_46/d__6_ xsel_46_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_5 XI11_6/XI0/XI0_46/d__5_ xsel_46_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_4 XI11_6/XI0/XI0_46/d__4_ xsel_46_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_3 XI11_6/XI0/XI0_46/d__3_ xsel_46_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_2 XI11_6/XI0/XI0_46/d__2_ xsel_46_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_1 XI11_6/XI0/XI0_46/d__1_ xsel_46_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_46/MN1_0 XI11_6/XI0/XI0_46/d__0_ xsel_46_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_15 XI11_6/net21_0_ xsel_45_ XI11_6/XI0/XI0_45/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_14 XI11_6/net21_1_ xsel_45_ XI11_6/XI0/XI0_45/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_13 XI11_6/net21_2_ xsel_45_ XI11_6/XI0/XI0_45/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_12 XI11_6/net21_3_ xsel_45_ XI11_6/XI0/XI0_45/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_11 XI11_6/net21_4_ xsel_45_ XI11_6/XI0/XI0_45/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_10 XI11_6/net21_5_ xsel_45_ XI11_6/XI0/XI0_45/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_9 XI11_6/net21_6_ xsel_45_ XI11_6/XI0/XI0_45/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_8 XI11_6/net21_7_ xsel_45_ XI11_6/XI0/XI0_45/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_7 XI11_6/net21_8_ xsel_45_ XI11_6/XI0/XI0_45/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_6 XI11_6/net21_9_ xsel_45_ XI11_6/XI0/XI0_45/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_5 XI11_6/net21_10_ xsel_45_ XI11_6/XI0/XI0_45/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_4 XI11_6/net21_11_ xsel_45_ XI11_6/XI0/XI0_45/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_3 XI11_6/net21_12_ xsel_45_ XI11_6/XI0/XI0_45/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_2 XI11_6/net21_13_ xsel_45_ XI11_6/XI0/XI0_45/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_1 XI11_6/net21_14_ xsel_45_ XI11_6/XI0/XI0_45/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN0_0 XI11_6/net21_15_ xsel_45_ XI11_6/XI0/XI0_45/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_15 XI11_6/XI0/XI0_45/d__15_ xsel_45_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_14 XI11_6/XI0/XI0_45/d__14_ xsel_45_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_13 XI11_6/XI0/XI0_45/d__13_ xsel_45_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_12 XI11_6/XI0/XI0_45/d__12_ xsel_45_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_11 XI11_6/XI0/XI0_45/d__11_ xsel_45_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_10 XI11_6/XI0/XI0_45/d__10_ xsel_45_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_9 XI11_6/XI0/XI0_45/d__9_ xsel_45_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_8 XI11_6/XI0/XI0_45/d__8_ xsel_45_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_7 XI11_6/XI0/XI0_45/d__7_ xsel_45_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_6 XI11_6/XI0/XI0_45/d__6_ xsel_45_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_5 XI11_6/XI0/XI0_45/d__5_ xsel_45_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_4 XI11_6/XI0/XI0_45/d__4_ xsel_45_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_3 XI11_6/XI0/XI0_45/d__3_ xsel_45_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_2 XI11_6/XI0/XI0_45/d__2_ xsel_45_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_1 XI11_6/XI0/XI0_45/d__1_ xsel_45_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_45/MN1_0 XI11_6/XI0/XI0_45/d__0_ xsel_45_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_15 XI11_6/net21_0_ xsel_44_ XI11_6/XI0/XI0_44/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_14 XI11_6/net21_1_ xsel_44_ XI11_6/XI0/XI0_44/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_13 XI11_6/net21_2_ xsel_44_ XI11_6/XI0/XI0_44/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_12 XI11_6/net21_3_ xsel_44_ XI11_6/XI0/XI0_44/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_11 XI11_6/net21_4_ xsel_44_ XI11_6/XI0/XI0_44/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_10 XI11_6/net21_5_ xsel_44_ XI11_6/XI0/XI0_44/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_9 XI11_6/net21_6_ xsel_44_ XI11_6/XI0/XI0_44/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_8 XI11_6/net21_7_ xsel_44_ XI11_6/XI0/XI0_44/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_7 XI11_6/net21_8_ xsel_44_ XI11_6/XI0/XI0_44/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_6 XI11_6/net21_9_ xsel_44_ XI11_6/XI0/XI0_44/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_5 XI11_6/net21_10_ xsel_44_ XI11_6/XI0/XI0_44/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_4 XI11_6/net21_11_ xsel_44_ XI11_6/XI0/XI0_44/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_3 XI11_6/net21_12_ xsel_44_ XI11_6/XI0/XI0_44/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_2 XI11_6/net21_13_ xsel_44_ XI11_6/XI0/XI0_44/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_1 XI11_6/net21_14_ xsel_44_ XI11_6/XI0/XI0_44/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN0_0 XI11_6/net21_15_ xsel_44_ XI11_6/XI0/XI0_44/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_15 XI11_6/XI0/XI0_44/d__15_ xsel_44_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_14 XI11_6/XI0/XI0_44/d__14_ xsel_44_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_13 XI11_6/XI0/XI0_44/d__13_ xsel_44_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_12 XI11_6/XI0/XI0_44/d__12_ xsel_44_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_11 XI11_6/XI0/XI0_44/d__11_ xsel_44_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_10 XI11_6/XI0/XI0_44/d__10_ xsel_44_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_9 XI11_6/XI0/XI0_44/d__9_ xsel_44_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_8 XI11_6/XI0/XI0_44/d__8_ xsel_44_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_7 XI11_6/XI0/XI0_44/d__7_ xsel_44_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_6 XI11_6/XI0/XI0_44/d__6_ xsel_44_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_5 XI11_6/XI0/XI0_44/d__5_ xsel_44_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_4 XI11_6/XI0/XI0_44/d__4_ xsel_44_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_3 XI11_6/XI0/XI0_44/d__3_ xsel_44_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_2 XI11_6/XI0/XI0_44/d__2_ xsel_44_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_1 XI11_6/XI0/XI0_44/d__1_ xsel_44_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_44/MN1_0 XI11_6/XI0/XI0_44/d__0_ xsel_44_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_15 XI11_6/net21_0_ xsel_43_ XI11_6/XI0/XI0_43/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_14 XI11_6/net21_1_ xsel_43_ XI11_6/XI0/XI0_43/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_13 XI11_6/net21_2_ xsel_43_ XI11_6/XI0/XI0_43/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_12 XI11_6/net21_3_ xsel_43_ XI11_6/XI0/XI0_43/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_11 XI11_6/net21_4_ xsel_43_ XI11_6/XI0/XI0_43/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_10 XI11_6/net21_5_ xsel_43_ XI11_6/XI0/XI0_43/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_9 XI11_6/net21_6_ xsel_43_ XI11_6/XI0/XI0_43/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_8 XI11_6/net21_7_ xsel_43_ XI11_6/XI0/XI0_43/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_7 XI11_6/net21_8_ xsel_43_ XI11_6/XI0/XI0_43/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_6 XI11_6/net21_9_ xsel_43_ XI11_6/XI0/XI0_43/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_5 XI11_6/net21_10_ xsel_43_ XI11_6/XI0/XI0_43/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_4 XI11_6/net21_11_ xsel_43_ XI11_6/XI0/XI0_43/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_3 XI11_6/net21_12_ xsel_43_ XI11_6/XI0/XI0_43/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_2 XI11_6/net21_13_ xsel_43_ XI11_6/XI0/XI0_43/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_1 XI11_6/net21_14_ xsel_43_ XI11_6/XI0/XI0_43/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN0_0 XI11_6/net21_15_ xsel_43_ XI11_6/XI0/XI0_43/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_15 XI11_6/XI0/XI0_43/d__15_ xsel_43_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_14 XI11_6/XI0/XI0_43/d__14_ xsel_43_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_13 XI11_6/XI0/XI0_43/d__13_ xsel_43_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_12 XI11_6/XI0/XI0_43/d__12_ xsel_43_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_11 XI11_6/XI0/XI0_43/d__11_ xsel_43_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_10 XI11_6/XI0/XI0_43/d__10_ xsel_43_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_9 XI11_6/XI0/XI0_43/d__9_ xsel_43_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_8 XI11_6/XI0/XI0_43/d__8_ xsel_43_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_7 XI11_6/XI0/XI0_43/d__7_ xsel_43_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_6 XI11_6/XI0/XI0_43/d__6_ xsel_43_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_5 XI11_6/XI0/XI0_43/d__5_ xsel_43_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_4 XI11_6/XI0/XI0_43/d__4_ xsel_43_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_3 XI11_6/XI0/XI0_43/d__3_ xsel_43_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_2 XI11_6/XI0/XI0_43/d__2_ xsel_43_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_1 XI11_6/XI0/XI0_43/d__1_ xsel_43_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_43/MN1_0 XI11_6/XI0/XI0_43/d__0_ xsel_43_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_15 XI11_6/net21_0_ xsel_42_ XI11_6/XI0/XI0_42/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_14 XI11_6/net21_1_ xsel_42_ XI11_6/XI0/XI0_42/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_13 XI11_6/net21_2_ xsel_42_ XI11_6/XI0/XI0_42/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_12 XI11_6/net21_3_ xsel_42_ XI11_6/XI0/XI0_42/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_11 XI11_6/net21_4_ xsel_42_ XI11_6/XI0/XI0_42/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_10 XI11_6/net21_5_ xsel_42_ XI11_6/XI0/XI0_42/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_9 XI11_6/net21_6_ xsel_42_ XI11_6/XI0/XI0_42/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_8 XI11_6/net21_7_ xsel_42_ XI11_6/XI0/XI0_42/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_7 XI11_6/net21_8_ xsel_42_ XI11_6/XI0/XI0_42/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_6 XI11_6/net21_9_ xsel_42_ XI11_6/XI0/XI0_42/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_5 XI11_6/net21_10_ xsel_42_ XI11_6/XI0/XI0_42/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_4 XI11_6/net21_11_ xsel_42_ XI11_6/XI0/XI0_42/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_3 XI11_6/net21_12_ xsel_42_ XI11_6/XI0/XI0_42/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_2 XI11_6/net21_13_ xsel_42_ XI11_6/XI0/XI0_42/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_1 XI11_6/net21_14_ xsel_42_ XI11_6/XI0/XI0_42/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN0_0 XI11_6/net21_15_ xsel_42_ XI11_6/XI0/XI0_42/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_15 XI11_6/XI0/XI0_42/d__15_ xsel_42_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_14 XI11_6/XI0/XI0_42/d__14_ xsel_42_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_13 XI11_6/XI0/XI0_42/d__13_ xsel_42_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_12 XI11_6/XI0/XI0_42/d__12_ xsel_42_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_11 XI11_6/XI0/XI0_42/d__11_ xsel_42_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_10 XI11_6/XI0/XI0_42/d__10_ xsel_42_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_9 XI11_6/XI0/XI0_42/d__9_ xsel_42_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_8 XI11_6/XI0/XI0_42/d__8_ xsel_42_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_7 XI11_6/XI0/XI0_42/d__7_ xsel_42_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_6 XI11_6/XI0/XI0_42/d__6_ xsel_42_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_5 XI11_6/XI0/XI0_42/d__5_ xsel_42_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_4 XI11_6/XI0/XI0_42/d__4_ xsel_42_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_3 XI11_6/XI0/XI0_42/d__3_ xsel_42_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_2 XI11_6/XI0/XI0_42/d__2_ xsel_42_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_1 XI11_6/XI0/XI0_42/d__1_ xsel_42_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_42/MN1_0 XI11_6/XI0/XI0_42/d__0_ xsel_42_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_15 XI11_6/net21_0_ xsel_41_ XI11_6/XI0/XI0_41/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_14 XI11_6/net21_1_ xsel_41_ XI11_6/XI0/XI0_41/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_13 XI11_6/net21_2_ xsel_41_ XI11_6/XI0/XI0_41/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_12 XI11_6/net21_3_ xsel_41_ XI11_6/XI0/XI0_41/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_11 XI11_6/net21_4_ xsel_41_ XI11_6/XI0/XI0_41/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_10 XI11_6/net21_5_ xsel_41_ XI11_6/XI0/XI0_41/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_9 XI11_6/net21_6_ xsel_41_ XI11_6/XI0/XI0_41/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_8 XI11_6/net21_7_ xsel_41_ XI11_6/XI0/XI0_41/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_7 XI11_6/net21_8_ xsel_41_ XI11_6/XI0/XI0_41/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_6 XI11_6/net21_9_ xsel_41_ XI11_6/XI0/XI0_41/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_5 XI11_6/net21_10_ xsel_41_ XI11_6/XI0/XI0_41/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_4 XI11_6/net21_11_ xsel_41_ XI11_6/XI0/XI0_41/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_3 XI11_6/net21_12_ xsel_41_ XI11_6/XI0/XI0_41/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_2 XI11_6/net21_13_ xsel_41_ XI11_6/XI0/XI0_41/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_1 XI11_6/net21_14_ xsel_41_ XI11_6/XI0/XI0_41/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN0_0 XI11_6/net21_15_ xsel_41_ XI11_6/XI0/XI0_41/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_15 XI11_6/XI0/XI0_41/d__15_ xsel_41_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_14 XI11_6/XI0/XI0_41/d__14_ xsel_41_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_13 XI11_6/XI0/XI0_41/d__13_ xsel_41_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_12 XI11_6/XI0/XI0_41/d__12_ xsel_41_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_11 XI11_6/XI0/XI0_41/d__11_ xsel_41_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_10 XI11_6/XI0/XI0_41/d__10_ xsel_41_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_9 XI11_6/XI0/XI0_41/d__9_ xsel_41_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_8 XI11_6/XI0/XI0_41/d__8_ xsel_41_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_7 XI11_6/XI0/XI0_41/d__7_ xsel_41_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_6 XI11_6/XI0/XI0_41/d__6_ xsel_41_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_5 XI11_6/XI0/XI0_41/d__5_ xsel_41_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_4 XI11_6/XI0/XI0_41/d__4_ xsel_41_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_3 XI11_6/XI0/XI0_41/d__3_ xsel_41_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_2 XI11_6/XI0/XI0_41/d__2_ xsel_41_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_1 XI11_6/XI0/XI0_41/d__1_ xsel_41_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_41/MN1_0 XI11_6/XI0/XI0_41/d__0_ xsel_41_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_15 XI11_6/net21_0_ xsel_40_ XI11_6/XI0/XI0_40/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_14 XI11_6/net21_1_ xsel_40_ XI11_6/XI0/XI0_40/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_13 XI11_6/net21_2_ xsel_40_ XI11_6/XI0/XI0_40/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_12 XI11_6/net21_3_ xsel_40_ XI11_6/XI0/XI0_40/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_11 XI11_6/net21_4_ xsel_40_ XI11_6/XI0/XI0_40/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_10 XI11_6/net21_5_ xsel_40_ XI11_6/XI0/XI0_40/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_9 XI11_6/net21_6_ xsel_40_ XI11_6/XI0/XI0_40/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_8 XI11_6/net21_7_ xsel_40_ XI11_6/XI0/XI0_40/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_7 XI11_6/net21_8_ xsel_40_ XI11_6/XI0/XI0_40/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_6 XI11_6/net21_9_ xsel_40_ XI11_6/XI0/XI0_40/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_5 XI11_6/net21_10_ xsel_40_ XI11_6/XI0/XI0_40/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_4 XI11_6/net21_11_ xsel_40_ XI11_6/XI0/XI0_40/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_3 XI11_6/net21_12_ xsel_40_ XI11_6/XI0/XI0_40/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_2 XI11_6/net21_13_ xsel_40_ XI11_6/XI0/XI0_40/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_1 XI11_6/net21_14_ xsel_40_ XI11_6/XI0/XI0_40/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN0_0 XI11_6/net21_15_ xsel_40_ XI11_6/XI0/XI0_40/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_15 XI11_6/XI0/XI0_40/d__15_ xsel_40_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_14 XI11_6/XI0/XI0_40/d__14_ xsel_40_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_13 XI11_6/XI0/XI0_40/d__13_ xsel_40_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_12 XI11_6/XI0/XI0_40/d__12_ xsel_40_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_11 XI11_6/XI0/XI0_40/d__11_ xsel_40_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_10 XI11_6/XI0/XI0_40/d__10_ xsel_40_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_9 XI11_6/XI0/XI0_40/d__9_ xsel_40_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_8 XI11_6/XI0/XI0_40/d__8_ xsel_40_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_7 XI11_6/XI0/XI0_40/d__7_ xsel_40_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_6 XI11_6/XI0/XI0_40/d__6_ xsel_40_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_5 XI11_6/XI0/XI0_40/d__5_ xsel_40_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_4 XI11_6/XI0/XI0_40/d__4_ xsel_40_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_3 XI11_6/XI0/XI0_40/d__3_ xsel_40_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_2 XI11_6/XI0/XI0_40/d__2_ xsel_40_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_1 XI11_6/XI0/XI0_40/d__1_ xsel_40_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_40/MN1_0 XI11_6/XI0/XI0_40/d__0_ xsel_40_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_15 XI11_6/net21_0_ xsel_39_ XI11_6/XI0/XI0_39/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_14 XI11_6/net21_1_ xsel_39_ XI11_6/XI0/XI0_39/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_13 XI11_6/net21_2_ xsel_39_ XI11_6/XI0/XI0_39/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_12 XI11_6/net21_3_ xsel_39_ XI11_6/XI0/XI0_39/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_11 XI11_6/net21_4_ xsel_39_ XI11_6/XI0/XI0_39/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_10 XI11_6/net21_5_ xsel_39_ XI11_6/XI0/XI0_39/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_9 XI11_6/net21_6_ xsel_39_ XI11_6/XI0/XI0_39/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_8 XI11_6/net21_7_ xsel_39_ XI11_6/XI0/XI0_39/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_7 XI11_6/net21_8_ xsel_39_ XI11_6/XI0/XI0_39/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_6 XI11_6/net21_9_ xsel_39_ XI11_6/XI0/XI0_39/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_5 XI11_6/net21_10_ xsel_39_ XI11_6/XI0/XI0_39/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_4 XI11_6/net21_11_ xsel_39_ XI11_6/XI0/XI0_39/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_3 XI11_6/net21_12_ xsel_39_ XI11_6/XI0/XI0_39/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_2 XI11_6/net21_13_ xsel_39_ XI11_6/XI0/XI0_39/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_1 XI11_6/net21_14_ xsel_39_ XI11_6/XI0/XI0_39/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN0_0 XI11_6/net21_15_ xsel_39_ XI11_6/XI0/XI0_39/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_15 XI11_6/XI0/XI0_39/d__15_ xsel_39_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_14 XI11_6/XI0/XI0_39/d__14_ xsel_39_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_13 XI11_6/XI0/XI0_39/d__13_ xsel_39_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_12 XI11_6/XI0/XI0_39/d__12_ xsel_39_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_11 XI11_6/XI0/XI0_39/d__11_ xsel_39_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_10 XI11_6/XI0/XI0_39/d__10_ xsel_39_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_9 XI11_6/XI0/XI0_39/d__9_ xsel_39_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_8 XI11_6/XI0/XI0_39/d__8_ xsel_39_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_7 XI11_6/XI0/XI0_39/d__7_ xsel_39_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_6 XI11_6/XI0/XI0_39/d__6_ xsel_39_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_5 XI11_6/XI0/XI0_39/d__5_ xsel_39_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_4 XI11_6/XI0/XI0_39/d__4_ xsel_39_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_3 XI11_6/XI0/XI0_39/d__3_ xsel_39_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_2 XI11_6/XI0/XI0_39/d__2_ xsel_39_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_1 XI11_6/XI0/XI0_39/d__1_ xsel_39_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_39/MN1_0 XI11_6/XI0/XI0_39/d__0_ xsel_39_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_15 XI11_6/net21_0_ xsel_38_ XI11_6/XI0/XI0_38/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_14 XI11_6/net21_1_ xsel_38_ XI11_6/XI0/XI0_38/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_13 XI11_6/net21_2_ xsel_38_ XI11_6/XI0/XI0_38/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_12 XI11_6/net21_3_ xsel_38_ XI11_6/XI0/XI0_38/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_11 XI11_6/net21_4_ xsel_38_ XI11_6/XI0/XI0_38/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_10 XI11_6/net21_5_ xsel_38_ XI11_6/XI0/XI0_38/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_9 XI11_6/net21_6_ xsel_38_ XI11_6/XI0/XI0_38/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_8 XI11_6/net21_7_ xsel_38_ XI11_6/XI0/XI0_38/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_7 XI11_6/net21_8_ xsel_38_ XI11_6/XI0/XI0_38/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_6 XI11_6/net21_9_ xsel_38_ XI11_6/XI0/XI0_38/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_5 XI11_6/net21_10_ xsel_38_ XI11_6/XI0/XI0_38/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_4 XI11_6/net21_11_ xsel_38_ XI11_6/XI0/XI0_38/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_3 XI11_6/net21_12_ xsel_38_ XI11_6/XI0/XI0_38/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_2 XI11_6/net21_13_ xsel_38_ XI11_6/XI0/XI0_38/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_1 XI11_6/net21_14_ xsel_38_ XI11_6/XI0/XI0_38/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN0_0 XI11_6/net21_15_ xsel_38_ XI11_6/XI0/XI0_38/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_15 XI11_6/XI0/XI0_38/d__15_ xsel_38_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_14 XI11_6/XI0/XI0_38/d__14_ xsel_38_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_13 XI11_6/XI0/XI0_38/d__13_ xsel_38_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_12 XI11_6/XI0/XI0_38/d__12_ xsel_38_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_11 XI11_6/XI0/XI0_38/d__11_ xsel_38_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_10 XI11_6/XI0/XI0_38/d__10_ xsel_38_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_9 XI11_6/XI0/XI0_38/d__9_ xsel_38_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_8 XI11_6/XI0/XI0_38/d__8_ xsel_38_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_7 XI11_6/XI0/XI0_38/d__7_ xsel_38_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_6 XI11_6/XI0/XI0_38/d__6_ xsel_38_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_5 XI11_6/XI0/XI0_38/d__5_ xsel_38_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_4 XI11_6/XI0/XI0_38/d__4_ xsel_38_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_3 XI11_6/XI0/XI0_38/d__3_ xsel_38_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_2 XI11_6/XI0/XI0_38/d__2_ xsel_38_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_1 XI11_6/XI0/XI0_38/d__1_ xsel_38_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_38/MN1_0 XI11_6/XI0/XI0_38/d__0_ xsel_38_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_15 XI11_6/net21_0_ xsel_37_ XI11_6/XI0/XI0_37/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_14 XI11_6/net21_1_ xsel_37_ XI11_6/XI0/XI0_37/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_13 XI11_6/net21_2_ xsel_37_ XI11_6/XI0/XI0_37/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_12 XI11_6/net21_3_ xsel_37_ XI11_6/XI0/XI0_37/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_11 XI11_6/net21_4_ xsel_37_ XI11_6/XI0/XI0_37/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_10 XI11_6/net21_5_ xsel_37_ XI11_6/XI0/XI0_37/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_9 XI11_6/net21_6_ xsel_37_ XI11_6/XI0/XI0_37/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_8 XI11_6/net21_7_ xsel_37_ XI11_6/XI0/XI0_37/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_7 XI11_6/net21_8_ xsel_37_ XI11_6/XI0/XI0_37/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_6 XI11_6/net21_9_ xsel_37_ XI11_6/XI0/XI0_37/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_5 XI11_6/net21_10_ xsel_37_ XI11_6/XI0/XI0_37/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_4 XI11_6/net21_11_ xsel_37_ XI11_6/XI0/XI0_37/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_3 XI11_6/net21_12_ xsel_37_ XI11_6/XI0/XI0_37/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_2 XI11_6/net21_13_ xsel_37_ XI11_6/XI0/XI0_37/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_1 XI11_6/net21_14_ xsel_37_ XI11_6/XI0/XI0_37/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN0_0 XI11_6/net21_15_ xsel_37_ XI11_6/XI0/XI0_37/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_15 XI11_6/XI0/XI0_37/d__15_ xsel_37_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_14 XI11_6/XI0/XI0_37/d__14_ xsel_37_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_13 XI11_6/XI0/XI0_37/d__13_ xsel_37_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_12 XI11_6/XI0/XI0_37/d__12_ xsel_37_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_11 XI11_6/XI0/XI0_37/d__11_ xsel_37_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_10 XI11_6/XI0/XI0_37/d__10_ xsel_37_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_9 XI11_6/XI0/XI0_37/d__9_ xsel_37_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_8 XI11_6/XI0/XI0_37/d__8_ xsel_37_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_7 XI11_6/XI0/XI0_37/d__7_ xsel_37_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_6 XI11_6/XI0/XI0_37/d__6_ xsel_37_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_5 XI11_6/XI0/XI0_37/d__5_ xsel_37_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_4 XI11_6/XI0/XI0_37/d__4_ xsel_37_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_3 XI11_6/XI0/XI0_37/d__3_ xsel_37_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_2 XI11_6/XI0/XI0_37/d__2_ xsel_37_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_1 XI11_6/XI0/XI0_37/d__1_ xsel_37_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_37/MN1_0 XI11_6/XI0/XI0_37/d__0_ xsel_37_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_15 XI11_6/net21_0_ xsel_36_ XI11_6/XI0/XI0_36/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_14 XI11_6/net21_1_ xsel_36_ XI11_6/XI0/XI0_36/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_13 XI11_6/net21_2_ xsel_36_ XI11_6/XI0/XI0_36/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_12 XI11_6/net21_3_ xsel_36_ XI11_6/XI0/XI0_36/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_11 XI11_6/net21_4_ xsel_36_ XI11_6/XI0/XI0_36/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_10 XI11_6/net21_5_ xsel_36_ XI11_6/XI0/XI0_36/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_9 XI11_6/net21_6_ xsel_36_ XI11_6/XI0/XI0_36/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_8 XI11_6/net21_7_ xsel_36_ XI11_6/XI0/XI0_36/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_7 XI11_6/net21_8_ xsel_36_ XI11_6/XI0/XI0_36/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_6 XI11_6/net21_9_ xsel_36_ XI11_6/XI0/XI0_36/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_5 XI11_6/net21_10_ xsel_36_ XI11_6/XI0/XI0_36/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_4 XI11_6/net21_11_ xsel_36_ XI11_6/XI0/XI0_36/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_3 XI11_6/net21_12_ xsel_36_ XI11_6/XI0/XI0_36/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_2 XI11_6/net21_13_ xsel_36_ XI11_6/XI0/XI0_36/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_1 XI11_6/net21_14_ xsel_36_ XI11_6/XI0/XI0_36/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN0_0 XI11_6/net21_15_ xsel_36_ XI11_6/XI0/XI0_36/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_15 XI11_6/XI0/XI0_36/d__15_ xsel_36_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_14 XI11_6/XI0/XI0_36/d__14_ xsel_36_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_13 XI11_6/XI0/XI0_36/d__13_ xsel_36_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_12 XI11_6/XI0/XI0_36/d__12_ xsel_36_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_11 XI11_6/XI0/XI0_36/d__11_ xsel_36_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_10 XI11_6/XI0/XI0_36/d__10_ xsel_36_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_9 XI11_6/XI0/XI0_36/d__9_ xsel_36_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_8 XI11_6/XI0/XI0_36/d__8_ xsel_36_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_7 XI11_6/XI0/XI0_36/d__7_ xsel_36_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_6 XI11_6/XI0/XI0_36/d__6_ xsel_36_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_5 XI11_6/XI0/XI0_36/d__5_ xsel_36_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_4 XI11_6/XI0/XI0_36/d__4_ xsel_36_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_3 XI11_6/XI0/XI0_36/d__3_ xsel_36_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_2 XI11_6/XI0/XI0_36/d__2_ xsel_36_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_1 XI11_6/XI0/XI0_36/d__1_ xsel_36_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_36/MN1_0 XI11_6/XI0/XI0_36/d__0_ xsel_36_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_15 XI11_6/net21_0_ xsel_35_ XI11_6/XI0/XI0_35/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_14 XI11_6/net21_1_ xsel_35_ XI11_6/XI0/XI0_35/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_13 XI11_6/net21_2_ xsel_35_ XI11_6/XI0/XI0_35/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_12 XI11_6/net21_3_ xsel_35_ XI11_6/XI0/XI0_35/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_11 XI11_6/net21_4_ xsel_35_ XI11_6/XI0/XI0_35/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_10 XI11_6/net21_5_ xsel_35_ XI11_6/XI0/XI0_35/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_9 XI11_6/net21_6_ xsel_35_ XI11_6/XI0/XI0_35/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_8 XI11_6/net21_7_ xsel_35_ XI11_6/XI0/XI0_35/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_7 XI11_6/net21_8_ xsel_35_ XI11_6/XI0/XI0_35/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_6 XI11_6/net21_9_ xsel_35_ XI11_6/XI0/XI0_35/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_5 XI11_6/net21_10_ xsel_35_ XI11_6/XI0/XI0_35/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_4 XI11_6/net21_11_ xsel_35_ XI11_6/XI0/XI0_35/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_3 XI11_6/net21_12_ xsel_35_ XI11_6/XI0/XI0_35/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_2 XI11_6/net21_13_ xsel_35_ XI11_6/XI0/XI0_35/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_1 XI11_6/net21_14_ xsel_35_ XI11_6/XI0/XI0_35/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN0_0 XI11_6/net21_15_ xsel_35_ XI11_6/XI0/XI0_35/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_15 XI11_6/XI0/XI0_35/d__15_ xsel_35_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_14 XI11_6/XI0/XI0_35/d__14_ xsel_35_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_13 XI11_6/XI0/XI0_35/d__13_ xsel_35_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_12 XI11_6/XI0/XI0_35/d__12_ xsel_35_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_11 XI11_6/XI0/XI0_35/d__11_ xsel_35_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_10 XI11_6/XI0/XI0_35/d__10_ xsel_35_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_9 XI11_6/XI0/XI0_35/d__9_ xsel_35_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_8 XI11_6/XI0/XI0_35/d__8_ xsel_35_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_7 XI11_6/XI0/XI0_35/d__7_ xsel_35_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_6 XI11_6/XI0/XI0_35/d__6_ xsel_35_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_5 XI11_6/XI0/XI0_35/d__5_ xsel_35_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_4 XI11_6/XI0/XI0_35/d__4_ xsel_35_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_3 XI11_6/XI0/XI0_35/d__3_ xsel_35_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_2 XI11_6/XI0/XI0_35/d__2_ xsel_35_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_1 XI11_6/XI0/XI0_35/d__1_ xsel_35_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_35/MN1_0 XI11_6/XI0/XI0_35/d__0_ xsel_35_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_15 XI11_6/net21_0_ xsel_34_ XI11_6/XI0/XI0_34/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_14 XI11_6/net21_1_ xsel_34_ XI11_6/XI0/XI0_34/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_13 XI11_6/net21_2_ xsel_34_ XI11_6/XI0/XI0_34/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_12 XI11_6/net21_3_ xsel_34_ XI11_6/XI0/XI0_34/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_11 XI11_6/net21_4_ xsel_34_ XI11_6/XI0/XI0_34/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_10 XI11_6/net21_5_ xsel_34_ XI11_6/XI0/XI0_34/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_9 XI11_6/net21_6_ xsel_34_ XI11_6/XI0/XI0_34/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_8 XI11_6/net21_7_ xsel_34_ XI11_6/XI0/XI0_34/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_7 XI11_6/net21_8_ xsel_34_ XI11_6/XI0/XI0_34/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_6 XI11_6/net21_9_ xsel_34_ XI11_6/XI0/XI0_34/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_5 XI11_6/net21_10_ xsel_34_ XI11_6/XI0/XI0_34/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_4 XI11_6/net21_11_ xsel_34_ XI11_6/XI0/XI0_34/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_3 XI11_6/net21_12_ xsel_34_ XI11_6/XI0/XI0_34/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_2 XI11_6/net21_13_ xsel_34_ XI11_6/XI0/XI0_34/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_1 XI11_6/net21_14_ xsel_34_ XI11_6/XI0/XI0_34/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN0_0 XI11_6/net21_15_ xsel_34_ XI11_6/XI0/XI0_34/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_15 XI11_6/XI0/XI0_34/d__15_ xsel_34_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_14 XI11_6/XI0/XI0_34/d__14_ xsel_34_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_13 XI11_6/XI0/XI0_34/d__13_ xsel_34_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_12 XI11_6/XI0/XI0_34/d__12_ xsel_34_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_11 XI11_6/XI0/XI0_34/d__11_ xsel_34_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_10 XI11_6/XI0/XI0_34/d__10_ xsel_34_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_9 XI11_6/XI0/XI0_34/d__9_ xsel_34_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_8 XI11_6/XI0/XI0_34/d__8_ xsel_34_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_7 XI11_6/XI0/XI0_34/d__7_ xsel_34_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_6 XI11_6/XI0/XI0_34/d__6_ xsel_34_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_5 XI11_6/XI0/XI0_34/d__5_ xsel_34_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_4 XI11_6/XI0/XI0_34/d__4_ xsel_34_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_3 XI11_6/XI0/XI0_34/d__3_ xsel_34_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_2 XI11_6/XI0/XI0_34/d__2_ xsel_34_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_1 XI11_6/XI0/XI0_34/d__1_ xsel_34_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_34/MN1_0 XI11_6/XI0/XI0_34/d__0_ xsel_34_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_15 XI11_6/net21_0_ xsel_33_ XI11_6/XI0/XI0_33/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_14 XI11_6/net21_1_ xsel_33_ XI11_6/XI0/XI0_33/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_13 XI11_6/net21_2_ xsel_33_ XI11_6/XI0/XI0_33/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_12 XI11_6/net21_3_ xsel_33_ XI11_6/XI0/XI0_33/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_11 XI11_6/net21_4_ xsel_33_ XI11_6/XI0/XI0_33/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_10 XI11_6/net21_5_ xsel_33_ XI11_6/XI0/XI0_33/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_9 XI11_6/net21_6_ xsel_33_ XI11_6/XI0/XI0_33/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_8 XI11_6/net21_7_ xsel_33_ XI11_6/XI0/XI0_33/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_7 XI11_6/net21_8_ xsel_33_ XI11_6/XI0/XI0_33/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_6 XI11_6/net21_9_ xsel_33_ XI11_6/XI0/XI0_33/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_5 XI11_6/net21_10_ xsel_33_ XI11_6/XI0/XI0_33/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_4 XI11_6/net21_11_ xsel_33_ XI11_6/XI0/XI0_33/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_3 XI11_6/net21_12_ xsel_33_ XI11_6/XI0/XI0_33/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_2 XI11_6/net21_13_ xsel_33_ XI11_6/XI0/XI0_33/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_1 XI11_6/net21_14_ xsel_33_ XI11_6/XI0/XI0_33/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN0_0 XI11_6/net21_15_ xsel_33_ XI11_6/XI0/XI0_33/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_15 XI11_6/XI0/XI0_33/d__15_ xsel_33_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_14 XI11_6/XI0/XI0_33/d__14_ xsel_33_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_13 XI11_6/XI0/XI0_33/d__13_ xsel_33_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_12 XI11_6/XI0/XI0_33/d__12_ xsel_33_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_11 XI11_6/XI0/XI0_33/d__11_ xsel_33_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_10 XI11_6/XI0/XI0_33/d__10_ xsel_33_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_9 XI11_6/XI0/XI0_33/d__9_ xsel_33_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_8 XI11_6/XI0/XI0_33/d__8_ xsel_33_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_7 XI11_6/XI0/XI0_33/d__7_ xsel_33_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_6 XI11_6/XI0/XI0_33/d__6_ xsel_33_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_5 XI11_6/XI0/XI0_33/d__5_ xsel_33_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_4 XI11_6/XI0/XI0_33/d__4_ xsel_33_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_3 XI11_6/XI0/XI0_33/d__3_ xsel_33_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_2 XI11_6/XI0/XI0_33/d__2_ xsel_33_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_1 XI11_6/XI0/XI0_33/d__1_ xsel_33_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_33/MN1_0 XI11_6/XI0/XI0_33/d__0_ xsel_33_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_15 XI11_6/net21_0_ xsel_32_ XI11_6/XI0/XI0_32/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_14 XI11_6/net21_1_ xsel_32_ XI11_6/XI0/XI0_32/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_13 XI11_6/net21_2_ xsel_32_ XI11_6/XI0/XI0_32/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_12 XI11_6/net21_3_ xsel_32_ XI11_6/XI0/XI0_32/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_11 XI11_6/net21_4_ xsel_32_ XI11_6/XI0/XI0_32/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_10 XI11_6/net21_5_ xsel_32_ XI11_6/XI0/XI0_32/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_9 XI11_6/net21_6_ xsel_32_ XI11_6/XI0/XI0_32/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_8 XI11_6/net21_7_ xsel_32_ XI11_6/XI0/XI0_32/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_7 XI11_6/net21_8_ xsel_32_ XI11_6/XI0/XI0_32/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_6 XI11_6/net21_9_ xsel_32_ XI11_6/XI0/XI0_32/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_5 XI11_6/net21_10_ xsel_32_ XI11_6/XI0/XI0_32/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_4 XI11_6/net21_11_ xsel_32_ XI11_6/XI0/XI0_32/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_3 XI11_6/net21_12_ xsel_32_ XI11_6/XI0/XI0_32/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_2 XI11_6/net21_13_ xsel_32_ XI11_6/XI0/XI0_32/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_1 XI11_6/net21_14_ xsel_32_ XI11_6/XI0/XI0_32/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN0_0 XI11_6/net21_15_ xsel_32_ XI11_6/XI0/XI0_32/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_15 XI11_6/XI0/XI0_32/d__15_ xsel_32_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_14 XI11_6/XI0/XI0_32/d__14_ xsel_32_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_13 XI11_6/XI0/XI0_32/d__13_ xsel_32_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_12 XI11_6/XI0/XI0_32/d__12_ xsel_32_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_11 XI11_6/XI0/XI0_32/d__11_ xsel_32_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_10 XI11_6/XI0/XI0_32/d__10_ xsel_32_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_9 XI11_6/XI0/XI0_32/d__9_ xsel_32_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_8 XI11_6/XI0/XI0_32/d__8_ xsel_32_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_7 XI11_6/XI0/XI0_32/d__7_ xsel_32_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_6 XI11_6/XI0/XI0_32/d__6_ xsel_32_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_5 XI11_6/XI0/XI0_32/d__5_ xsel_32_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_4 XI11_6/XI0/XI0_32/d__4_ xsel_32_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_3 XI11_6/XI0/XI0_32/d__3_ xsel_32_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_2 XI11_6/XI0/XI0_32/d__2_ xsel_32_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_1 XI11_6/XI0/XI0_32/d__1_ xsel_32_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_32/MN1_0 XI11_6/XI0/XI0_32/d__0_ xsel_32_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_15 XI11_6/net21_0_ xsel_31_ XI11_6/XI0/XI0_31/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_14 XI11_6/net21_1_ xsel_31_ XI11_6/XI0/XI0_31/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_13 XI11_6/net21_2_ xsel_31_ XI11_6/XI0/XI0_31/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_12 XI11_6/net21_3_ xsel_31_ XI11_6/XI0/XI0_31/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_11 XI11_6/net21_4_ xsel_31_ XI11_6/XI0/XI0_31/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_10 XI11_6/net21_5_ xsel_31_ XI11_6/XI0/XI0_31/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_9 XI11_6/net21_6_ xsel_31_ XI11_6/XI0/XI0_31/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_8 XI11_6/net21_7_ xsel_31_ XI11_6/XI0/XI0_31/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_7 XI11_6/net21_8_ xsel_31_ XI11_6/XI0/XI0_31/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_6 XI11_6/net21_9_ xsel_31_ XI11_6/XI0/XI0_31/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_5 XI11_6/net21_10_ xsel_31_ XI11_6/XI0/XI0_31/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_4 XI11_6/net21_11_ xsel_31_ XI11_6/XI0/XI0_31/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_3 XI11_6/net21_12_ xsel_31_ XI11_6/XI0/XI0_31/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_2 XI11_6/net21_13_ xsel_31_ XI11_6/XI0/XI0_31/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_1 XI11_6/net21_14_ xsel_31_ XI11_6/XI0/XI0_31/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN0_0 XI11_6/net21_15_ xsel_31_ XI11_6/XI0/XI0_31/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_15 XI11_6/XI0/XI0_31/d__15_ xsel_31_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_14 XI11_6/XI0/XI0_31/d__14_ xsel_31_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_13 XI11_6/XI0/XI0_31/d__13_ xsel_31_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_12 XI11_6/XI0/XI0_31/d__12_ xsel_31_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_11 XI11_6/XI0/XI0_31/d__11_ xsel_31_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_10 XI11_6/XI0/XI0_31/d__10_ xsel_31_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_9 XI11_6/XI0/XI0_31/d__9_ xsel_31_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_8 XI11_6/XI0/XI0_31/d__8_ xsel_31_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_7 XI11_6/XI0/XI0_31/d__7_ xsel_31_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_6 XI11_6/XI0/XI0_31/d__6_ xsel_31_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_5 XI11_6/XI0/XI0_31/d__5_ xsel_31_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_4 XI11_6/XI0/XI0_31/d__4_ xsel_31_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_3 XI11_6/XI0/XI0_31/d__3_ xsel_31_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_2 XI11_6/XI0/XI0_31/d__2_ xsel_31_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_1 XI11_6/XI0/XI0_31/d__1_ xsel_31_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_31/MN1_0 XI11_6/XI0/XI0_31/d__0_ xsel_31_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_15 XI11_6/net21_0_ xsel_30_ XI11_6/XI0/XI0_30/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_14 XI11_6/net21_1_ xsel_30_ XI11_6/XI0/XI0_30/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_13 XI11_6/net21_2_ xsel_30_ XI11_6/XI0/XI0_30/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_12 XI11_6/net21_3_ xsel_30_ XI11_6/XI0/XI0_30/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_11 XI11_6/net21_4_ xsel_30_ XI11_6/XI0/XI0_30/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_10 XI11_6/net21_5_ xsel_30_ XI11_6/XI0/XI0_30/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_9 XI11_6/net21_6_ xsel_30_ XI11_6/XI0/XI0_30/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_8 XI11_6/net21_7_ xsel_30_ XI11_6/XI0/XI0_30/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_7 XI11_6/net21_8_ xsel_30_ XI11_6/XI0/XI0_30/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_6 XI11_6/net21_9_ xsel_30_ XI11_6/XI0/XI0_30/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_5 XI11_6/net21_10_ xsel_30_ XI11_6/XI0/XI0_30/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_4 XI11_6/net21_11_ xsel_30_ XI11_6/XI0/XI0_30/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_3 XI11_6/net21_12_ xsel_30_ XI11_6/XI0/XI0_30/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_2 XI11_6/net21_13_ xsel_30_ XI11_6/XI0/XI0_30/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_1 XI11_6/net21_14_ xsel_30_ XI11_6/XI0/XI0_30/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN0_0 XI11_6/net21_15_ xsel_30_ XI11_6/XI0/XI0_30/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_15 XI11_6/XI0/XI0_30/d__15_ xsel_30_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_14 XI11_6/XI0/XI0_30/d__14_ xsel_30_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_13 XI11_6/XI0/XI0_30/d__13_ xsel_30_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_12 XI11_6/XI0/XI0_30/d__12_ xsel_30_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_11 XI11_6/XI0/XI0_30/d__11_ xsel_30_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_10 XI11_6/XI0/XI0_30/d__10_ xsel_30_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_9 XI11_6/XI0/XI0_30/d__9_ xsel_30_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_8 XI11_6/XI0/XI0_30/d__8_ xsel_30_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_7 XI11_6/XI0/XI0_30/d__7_ xsel_30_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_6 XI11_6/XI0/XI0_30/d__6_ xsel_30_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_5 XI11_6/XI0/XI0_30/d__5_ xsel_30_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_4 XI11_6/XI0/XI0_30/d__4_ xsel_30_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_3 XI11_6/XI0/XI0_30/d__3_ xsel_30_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_2 XI11_6/XI0/XI0_30/d__2_ xsel_30_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_1 XI11_6/XI0/XI0_30/d__1_ xsel_30_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_30/MN1_0 XI11_6/XI0/XI0_30/d__0_ xsel_30_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_15 XI11_6/net21_0_ xsel_29_ XI11_6/XI0/XI0_29/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_14 XI11_6/net21_1_ xsel_29_ XI11_6/XI0/XI0_29/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_13 XI11_6/net21_2_ xsel_29_ XI11_6/XI0/XI0_29/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_12 XI11_6/net21_3_ xsel_29_ XI11_6/XI0/XI0_29/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_11 XI11_6/net21_4_ xsel_29_ XI11_6/XI0/XI0_29/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_10 XI11_6/net21_5_ xsel_29_ XI11_6/XI0/XI0_29/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_9 XI11_6/net21_6_ xsel_29_ XI11_6/XI0/XI0_29/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_8 XI11_6/net21_7_ xsel_29_ XI11_6/XI0/XI0_29/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_7 XI11_6/net21_8_ xsel_29_ XI11_6/XI0/XI0_29/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_6 XI11_6/net21_9_ xsel_29_ XI11_6/XI0/XI0_29/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_5 XI11_6/net21_10_ xsel_29_ XI11_6/XI0/XI0_29/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_4 XI11_6/net21_11_ xsel_29_ XI11_6/XI0/XI0_29/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_3 XI11_6/net21_12_ xsel_29_ XI11_6/XI0/XI0_29/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_2 XI11_6/net21_13_ xsel_29_ XI11_6/XI0/XI0_29/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_1 XI11_6/net21_14_ xsel_29_ XI11_6/XI0/XI0_29/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN0_0 XI11_6/net21_15_ xsel_29_ XI11_6/XI0/XI0_29/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_15 XI11_6/XI0/XI0_29/d__15_ xsel_29_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_14 XI11_6/XI0/XI0_29/d__14_ xsel_29_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_13 XI11_6/XI0/XI0_29/d__13_ xsel_29_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_12 XI11_6/XI0/XI0_29/d__12_ xsel_29_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_11 XI11_6/XI0/XI0_29/d__11_ xsel_29_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_10 XI11_6/XI0/XI0_29/d__10_ xsel_29_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_9 XI11_6/XI0/XI0_29/d__9_ xsel_29_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_8 XI11_6/XI0/XI0_29/d__8_ xsel_29_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_7 XI11_6/XI0/XI0_29/d__7_ xsel_29_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_6 XI11_6/XI0/XI0_29/d__6_ xsel_29_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_5 XI11_6/XI0/XI0_29/d__5_ xsel_29_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_4 XI11_6/XI0/XI0_29/d__4_ xsel_29_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_3 XI11_6/XI0/XI0_29/d__3_ xsel_29_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_2 XI11_6/XI0/XI0_29/d__2_ xsel_29_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_1 XI11_6/XI0/XI0_29/d__1_ xsel_29_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_29/MN1_0 XI11_6/XI0/XI0_29/d__0_ xsel_29_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_15 XI11_6/net21_0_ xsel_28_ XI11_6/XI0/XI0_28/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_14 XI11_6/net21_1_ xsel_28_ XI11_6/XI0/XI0_28/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_13 XI11_6/net21_2_ xsel_28_ XI11_6/XI0/XI0_28/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_12 XI11_6/net21_3_ xsel_28_ XI11_6/XI0/XI0_28/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_11 XI11_6/net21_4_ xsel_28_ XI11_6/XI0/XI0_28/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_10 XI11_6/net21_5_ xsel_28_ XI11_6/XI0/XI0_28/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_9 XI11_6/net21_6_ xsel_28_ XI11_6/XI0/XI0_28/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_8 XI11_6/net21_7_ xsel_28_ XI11_6/XI0/XI0_28/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_7 XI11_6/net21_8_ xsel_28_ XI11_6/XI0/XI0_28/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_6 XI11_6/net21_9_ xsel_28_ XI11_6/XI0/XI0_28/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_5 XI11_6/net21_10_ xsel_28_ XI11_6/XI0/XI0_28/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_4 XI11_6/net21_11_ xsel_28_ XI11_6/XI0/XI0_28/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_3 XI11_6/net21_12_ xsel_28_ XI11_6/XI0/XI0_28/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_2 XI11_6/net21_13_ xsel_28_ XI11_6/XI0/XI0_28/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_1 XI11_6/net21_14_ xsel_28_ XI11_6/XI0/XI0_28/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN0_0 XI11_6/net21_15_ xsel_28_ XI11_6/XI0/XI0_28/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_15 XI11_6/XI0/XI0_28/d__15_ xsel_28_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_14 XI11_6/XI0/XI0_28/d__14_ xsel_28_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_13 XI11_6/XI0/XI0_28/d__13_ xsel_28_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_12 XI11_6/XI0/XI0_28/d__12_ xsel_28_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_11 XI11_6/XI0/XI0_28/d__11_ xsel_28_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_10 XI11_6/XI0/XI0_28/d__10_ xsel_28_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_9 XI11_6/XI0/XI0_28/d__9_ xsel_28_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_8 XI11_6/XI0/XI0_28/d__8_ xsel_28_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_7 XI11_6/XI0/XI0_28/d__7_ xsel_28_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_6 XI11_6/XI0/XI0_28/d__6_ xsel_28_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_5 XI11_6/XI0/XI0_28/d__5_ xsel_28_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_4 XI11_6/XI0/XI0_28/d__4_ xsel_28_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_3 XI11_6/XI0/XI0_28/d__3_ xsel_28_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_2 XI11_6/XI0/XI0_28/d__2_ xsel_28_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_1 XI11_6/XI0/XI0_28/d__1_ xsel_28_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_28/MN1_0 XI11_6/XI0/XI0_28/d__0_ xsel_28_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_15 XI11_6/net21_0_ xsel_27_ XI11_6/XI0/XI0_27/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_14 XI11_6/net21_1_ xsel_27_ XI11_6/XI0/XI0_27/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_13 XI11_6/net21_2_ xsel_27_ XI11_6/XI0/XI0_27/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_12 XI11_6/net21_3_ xsel_27_ XI11_6/XI0/XI0_27/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_11 XI11_6/net21_4_ xsel_27_ XI11_6/XI0/XI0_27/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_10 XI11_6/net21_5_ xsel_27_ XI11_6/XI0/XI0_27/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_9 XI11_6/net21_6_ xsel_27_ XI11_6/XI0/XI0_27/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_8 XI11_6/net21_7_ xsel_27_ XI11_6/XI0/XI0_27/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_7 XI11_6/net21_8_ xsel_27_ XI11_6/XI0/XI0_27/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_6 XI11_6/net21_9_ xsel_27_ XI11_6/XI0/XI0_27/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_5 XI11_6/net21_10_ xsel_27_ XI11_6/XI0/XI0_27/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_4 XI11_6/net21_11_ xsel_27_ XI11_6/XI0/XI0_27/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_3 XI11_6/net21_12_ xsel_27_ XI11_6/XI0/XI0_27/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_2 XI11_6/net21_13_ xsel_27_ XI11_6/XI0/XI0_27/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_1 XI11_6/net21_14_ xsel_27_ XI11_6/XI0/XI0_27/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN0_0 XI11_6/net21_15_ xsel_27_ XI11_6/XI0/XI0_27/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_15 XI11_6/XI0/XI0_27/d__15_ xsel_27_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_14 XI11_6/XI0/XI0_27/d__14_ xsel_27_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_13 XI11_6/XI0/XI0_27/d__13_ xsel_27_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_12 XI11_6/XI0/XI0_27/d__12_ xsel_27_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_11 XI11_6/XI0/XI0_27/d__11_ xsel_27_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_10 XI11_6/XI0/XI0_27/d__10_ xsel_27_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_9 XI11_6/XI0/XI0_27/d__9_ xsel_27_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_8 XI11_6/XI0/XI0_27/d__8_ xsel_27_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_7 XI11_6/XI0/XI0_27/d__7_ xsel_27_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_6 XI11_6/XI0/XI0_27/d__6_ xsel_27_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_5 XI11_6/XI0/XI0_27/d__5_ xsel_27_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_4 XI11_6/XI0/XI0_27/d__4_ xsel_27_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_3 XI11_6/XI0/XI0_27/d__3_ xsel_27_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_2 XI11_6/XI0/XI0_27/d__2_ xsel_27_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_1 XI11_6/XI0/XI0_27/d__1_ xsel_27_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_27/MN1_0 XI11_6/XI0/XI0_27/d__0_ xsel_27_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_15 XI11_6/net21_0_ xsel_26_ XI11_6/XI0/XI0_26/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_14 XI11_6/net21_1_ xsel_26_ XI11_6/XI0/XI0_26/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_13 XI11_6/net21_2_ xsel_26_ XI11_6/XI0/XI0_26/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_12 XI11_6/net21_3_ xsel_26_ XI11_6/XI0/XI0_26/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_11 XI11_6/net21_4_ xsel_26_ XI11_6/XI0/XI0_26/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_10 XI11_6/net21_5_ xsel_26_ XI11_6/XI0/XI0_26/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_9 XI11_6/net21_6_ xsel_26_ XI11_6/XI0/XI0_26/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_8 XI11_6/net21_7_ xsel_26_ XI11_6/XI0/XI0_26/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_7 XI11_6/net21_8_ xsel_26_ XI11_6/XI0/XI0_26/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_6 XI11_6/net21_9_ xsel_26_ XI11_6/XI0/XI0_26/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_5 XI11_6/net21_10_ xsel_26_ XI11_6/XI0/XI0_26/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_4 XI11_6/net21_11_ xsel_26_ XI11_6/XI0/XI0_26/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_3 XI11_6/net21_12_ xsel_26_ XI11_6/XI0/XI0_26/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_2 XI11_6/net21_13_ xsel_26_ XI11_6/XI0/XI0_26/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_1 XI11_6/net21_14_ xsel_26_ XI11_6/XI0/XI0_26/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN0_0 XI11_6/net21_15_ xsel_26_ XI11_6/XI0/XI0_26/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_15 XI11_6/XI0/XI0_26/d__15_ xsel_26_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_14 XI11_6/XI0/XI0_26/d__14_ xsel_26_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_13 XI11_6/XI0/XI0_26/d__13_ xsel_26_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_12 XI11_6/XI0/XI0_26/d__12_ xsel_26_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_11 XI11_6/XI0/XI0_26/d__11_ xsel_26_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_10 XI11_6/XI0/XI0_26/d__10_ xsel_26_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_9 XI11_6/XI0/XI0_26/d__9_ xsel_26_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_8 XI11_6/XI0/XI0_26/d__8_ xsel_26_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_7 XI11_6/XI0/XI0_26/d__7_ xsel_26_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_6 XI11_6/XI0/XI0_26/d__6_ xsel_26_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_5 XI11_6/XI0/XI0_26/d__5_ xsel_26_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_4 XI11_6/XI0/XI0_26/d__4_ xsel_26_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_3 XI11_6/XI0/XI0_26/d__3_ xsel_26_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_2 XI11_6/XI0/XI0_26/d__2_ xsel_26_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_1 XI11_6/XI0/XI0_26/d__1_ xsel_26_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_26/MN1_0 XI11_6/XI0/XI0_26/d__0_ xsel_26_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_15 XI11_6/net21_0_ xsel_25_ XI11_6/XI0/XI0_25/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_14 XI11_6/net21_1_ xsel_25_ XI11_6/XI0/XI0_25/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_13 XI11_6/net21_2_ xsel_25_ XI11_6/XI0/XI0_25/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_12 XI11_6/net21_3_ xsel_25_ XI11_6/XI0/XI0_25/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_11 XI11_6/net21_4_ xsel_25_ XI11_6/XI0/XI0_25/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_10 XI11_6/net21_5_ xsel_25_ XI11_6/XI0/XI0_25/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_9 XI11_6/net21_6_ xsel_25_ XI11_6/XI0/XI0_25/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_8 XI11_6/net21_7_ xsel_25_ XI11_6/XI0/XI0_25/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_7 XI11_6/net21_8_ xsel_25_ XI11_6/XI0/XI0_25/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_6 XI11_6/net21_9_ xsel_25_ XI11_6/XI0/XI0_25/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_5 XI11_6/net21_10_ xsel_25_ XI11_6/XI0/XI0_25/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_4 XI11_6/net21_11_ xsel_25_ XI11_6/XI0/XI0_25/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_3 XI11_6/net21_12_ xsel_25_ XI11_6/XI0/XI0_25/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_2 XI11_6/net21_13_ xsel_25_ XI11_6/XI0/XI0_25/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_1 XI11_6/net21_14_ xsel_25_ XI11_6/XI0/XI0_25/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN0_0 XI11_6/net21_15_ xsel_25_ XI11_6/XI0/XI0_25/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_15 XI11_6/XI0/XI0_25/d__15_ xsel_25_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_14 XI11_6/XI0/XI0_25/d__14_ xsel_25_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_13 XI11_6/XI0/XI0_25/d__13_ xsel_25_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_12 XI11_6/XI0/XI0_25/d__12_ xsel_25_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_11 XI11_6/XI0/XI0_25/d__11_ xsel_25_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_10 XI11_6/XI0/XI0_25/d__10_ xsel_25_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_9 XI11_6/XI0/XI0_25/d__9_ xsel_25_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_8 XI11_6/XI0/XI0_25/d__8_ xsel_25_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_7 XI11_6/XI0/XI0_25/d__7_ xsel_25_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_6 XI11_6/XI0/XI0_25/d__6_ xsel_25_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_5 XI11_6/XI0/XI0_25/d__5_ xsel_25_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_4 XI11_6/XI0/XI0_25/d__4_ xsel_25_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_3 XI11_6/XI0/XI0_25/d__3_ xsel_25_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_2 XI11_6/XI0/XI0_25/d__2_ xsel_25_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_1 XI11_6/XI0/XI0_25/d__1_ xsel_25_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_25/MN1_0 XI11_6/XI0/XI0_25/d__0_ xsel_25_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_15 XI11_6/net21_0_ xsel_24_ XI11_6/XI0/XI0_24/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_14 XI11_6/net21_1_ xsel_24_ XI11_6/XI0/XI0_24/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_13 XI11_6/net21_2_ xsel_24_ XI11_6/XI0/XI0_24/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_12 XI11_6/net21_3_ xsel_24_ XI11_6/XI0/XI0_24/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_11 XI11_6/net21_4_ xsel_24_ XI11_6/XI0/XI0_24/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_10 XI11_6/net21_5_ xsel_24_ XI11_6/XI0/XI0_24/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_9 XI11_6/net21_6_ xsel_24_ XI11_6/XI0/XI0_24/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_8 XI11_6/net21_7_ xsel_24_ XI11_6/XI0/XI0_24/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_7 XI11_6/net21_8_ xsel_24_ XI11_6/XI0/XI0_24/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_6 XI11_6/net21_9_ xsel_24_ XI11_6/XI0/XI0_24/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_5 XI11_6/net21_10_ xsel_24_ XI11_6/XI0/XI0_24/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_4 XI11_6/net21_11_ xsel_24_ XI11_6/XI0/XI0_24/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_3 XI11_6/net21_12_ xsel_24_ XI11_6/XI0/XI0_24/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_2 XI11_6/net21_13_ xsel_24_ XI11_6/XI0/XI0_24/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_1 XI11_6/net21_14_ xsel_24_ XI11_6/XI0/XI0_24/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN0_0 XI11_6/net21_15_ xsel_24_ XI11_6/XI0/XI0_24/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_15 XI11_6/XI0/XI0_24/d__15_ xsel_24_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_14 XI11_6/XI0/XI0_24/d__14_ xsel_24_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_13 XI11_6/XI0/XI0_24/d__13_ xsel_24_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_12 XI11_6/XI0/XI0_24/d__12_ xsel_24_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_11 XI11_6/XI0/XI0_24/d__11_ xsel_24_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_10 XI11_6/XI0/XI0_24/d__10_ xsel_24_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_9 XI11_6/XI0/XI0_24/d__9_ xsel_24_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_8 XI11_6/XI0/XI0_24/d__8_ xsel_24_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_7 XI11_6/XI0/XI0_24/d__7_ xsel_24_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_6 XI11_6/XI0/XI0_24/d__6_ xsel_24_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_5 XI11_6/XI0/XI0_24/d__5_ xsel_24_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_4 XI11_6/XI0/XI0_24/d__4_ xsel_24_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_3 XI11_6/XI0/XI0_24/d__3_ xsel_24_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_2 XI11_6/XI0/XI0_24/d__2_ xsel_24_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_1 XI11_6/XI0/XI0_24/d__1_ xsel_24_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_24/MN1_0 XI11_6/XI0/XI0_24/d__0_ xsel_24_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_15 XI11_6/net21_0_ xsel_23_ XI11_6/XI0/XI0_23/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_14 XI11_6/net21_1_ xsel_23_ XI11_6/XI0/XI0_23/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_13 XI11_6/net21_2_ xsel_23_ XI11_6/XI0/XI0_23/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_12 XI11_6/net21_3_ xsel_23_ XI11_6/XI0/XI0_23/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_11 XI11_6/net21_4_ xsel_23_ XI11_6/XI0/XI0_23/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_10 XI11_6/net21_5_ xsel_23_ XI11_6/XI0/XI0_23/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_9 XI11_6/net21_6_ xsel_23_ XI11_6/XI0/XI0_23/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_8 XI11_6/net21_7_ xsel_23_ XI11_6/XI0/XI0_23/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_7 XI11_6/net21_8_ xsel_23_ XI11_6/XI0/XI0_23/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_6 XI11_6/net21_9_ xsel_23_ XI11_6/XI0/XI0_23/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_5 XI11_6/net21_10_ xsel_23_ XI11_6/XI0/XI0_23/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_4 XI11_6/net21_11_ xsel_23_ XI11_6/XI0/XI0_23/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_3 XI11_6/net21_12_ xsel_23_ XI11_6/XI0/XI0_23/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_2 XI11_6/net21_13_ xsel_23_ XI11_6/XI0/XI0_23/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_1 XI11_6/net21_14_ xsel_23_ XI11_6/XI0/XI0_23/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN0_0 XI11_6/net21_15_ xsel_23_ XI11_6/XI0/XI0_23/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_15 XI11_6/XI0/XI0_23/d__15_ xsel_23_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_14 XI11_6/XI0/XI0_23/d__14_ xsel_23_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_13 XI11_6/XI0/XI0_23/d__13_ xsel_23_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_12 XI11_6/XI0/XI0_23/d__12_ xsel_23_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_11 XI11_6/XI0/XI0_23/d__11_ xsel_23_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_10 XI11_6/XI0/XI0_23/d__10_ xsel_23_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_9 XI11_6/XI0/XI0_23/d__9_ xsel_23_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_8 XI11_6/XI0/XI0_23/d__8_ xsel_23_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_7 XI11_6/XI0/XI0_23/d__7_ xsel_23_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_6 XI11_6/XI0/XI0_23/d__6_ xsel_23_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_5 XI11_6/XI0/XI0_23/d__5_ xsel_23_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_4 XI11_6/XI0/XI0_23/d__4_ xsel_23_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_3 XI11_6/XI0/XI0_23/d__3_ xsel_23_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_2 XI11_6/XI0/XI0_23/d__2_ xsel_23_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_1 XI11_6/XI0/XI0_23/d__1_ xsel_23_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_23/MN1_0 XI11_6/XI0/XI0_23/d__0_ xsel_23_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_15 XI11_6/net21_0_ xsel_22_ XI11_6/XI0/XI0_22/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_14 XI11_6/net21_1_ xsel_22_ XI11_6/XI0/XI0_22/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_13 XI11_6/net21_2_ xsel_22_ XI11_6/XI0/XI0_22/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_12 XI11_6/net21_3_ xsel_22_ XI11_6/XI0/XI0_22/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_11 XI11_6/net21_4_ xsel_22_ XI11_6/XI0/XI0_22/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_10 XI11_6/net21_5_ xsel_22_ XI11_6/XI0/XI0_22/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_9 XI11_6/net21_6_ xsel_22_ XI11_6/XI0/XI0_22/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_8 XI11_6/net21_7_ xsel_22_ XI11_6/XI0/XI0_22/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_7 XI11_6/net21_8_ xsel_22_ XI11_6/XI0/XI0_22/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_6 XI11_6/net21_9_ xsel_22_ XI11_6/XI0/XI0_22/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_5 XI11_6/net21_10_ xsel_22_ XI11_6/XI0/XI0_22/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_4 XI11_6/net21_11_ xsel_22_ XI11_6/XI0/XI0_22/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_3 XI11_6/net21_12_ xsel_22_ XI11_6/XI0/XI0_22/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_2 XI11_6/net21_13_ xsel_22_ XI11_6/XI0/XI0_22/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_1 XI11_6/net21_14_ xsel_22_ XI11_6/XI0/XI0_22/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN0_0 XI11_6/net21_15_ xsel_22_ XI11_6/XI0/XI0_22/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_15 XI11_6/XI0/XI0_22/d__15_ xsel_22_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_14 XI11_6/XI0/XI0_22/d__14_ xsel_22_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_13 XI11_6/XI0/XI0_22/d__13_ xsel_22_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_12 XI11_6/XI0/XI0_22/d__12_ xsel_22_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_11 XI11_6/XI0/XI0_22/d__11_ xsel_22_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_10 XI11_6/XI0/XI0_22/d__10_ xsel_22_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_9 XI11_6/XI0/XI0_22/d__9_ xsel_22_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_8 XI11_6/XI0/XI0_22/d__8_ xsel_22_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_7 XI11_6/XI0/XI0_22/d__7_ xsel_22_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_6 XI11_6/XI0/XI0_22/d__6_ xsel_22_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_5 XI11_6/XI0/XI0_22/d__5_ xsel_22_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_4 XI11_6/XI0/XI0_22/d__4_ xsel_22_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_3 XI11_6/XI0/XI0_22/d__3_ xsel_22_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_2 XI11_6/XI0/XI0_22/d__2_ xsel_22_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_1 XI11_6/XI0/XI0_22/d__1_ xsel_22_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_22/MN1_0 XI11_6/XI0/XI0_22/d__0_ xsel_22_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_15 XI11_6/net21_0_ xsel_21_ XI11_6/XI0/XI0_21/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_14 XI11_6/net21_1_ xsel_21_ XI11_6/XI0/XI0_21/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_13 XI11_6/net21_2_ xsel_21_ XI11_6/XI0/XI0_21/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_12 XI11_6/net21_3_ xsel_21_ XI11_6/XI0/XI0_21/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_11 XI11_6/net21_4_ xsel_21_ XI11_6/XI0/XI0_21/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_10 XI11_6/net21_5_ xsel_21_ XI11_6/XI0/XI0_21/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_9 XI11_6/net21_6_ xsel_21_ XI11_6/XI0/XI0_21/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_8 XI11_6/net21_7_ xsel_21_ XI11_6/XI0/XI0_21/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_7 XI11_6/net21_8_ xsel_21_ XI11_6/XI0/XI0_21/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_6 XI11_6/net21_9_ xsel_21_ XI11_6/XI0/XI0_21/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_5 XI11_6/net21_10_ xsel_21_ XI11_6/XI0/XI0_21/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_4 XI11_6/net21_11_ xsel_21_ XI11_6/XI0/XI0_21/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_3 XI11_6/net21_12_ xsel_21_ XI11_6/XI0/XI0_21/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_2 XI11_6/net21_13_ xsel_21_ XI11_6/XI0/XI0_21/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_1 XI11_6/net21_14_ xsel_21_ XI11_6/XI0/XI0_21/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN0_0 XI11_6/net21_15_ xsel_21_ XI11_6/XI0/XI0_21/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_15 XI11_6/XI0/XI0_21/d__15_ xsel_21_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_14 XI11_6/XI0/XI0_21/d__14_ xsel_21_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_13 XI11_6/XI0/XI0_21/d__13_ xsel_21_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_12 XI11_6/XI0/XI0_21/d__12_ xsel_21_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_11 XI11_6/XI0/XI0_21/d__11_ xsel_21_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_10 XI11_6/XI0/XI0_21/d__10_ xsel_21_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_9 XI11_6/XI0/XI0_21/d__9_ xsel_21_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_8 XI11_6/XI0/XI0_21/d__8_ xsel_21_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_7 XI11_6/XI0/XI0_21/d__7_ xsel_21_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_6 XI11_6/XI0/XI0_21/d__6_ xsel_21_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_5 XI11_6/XI0/XI0_21/d__5_ xsel_21_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_4 XI11_6/XI0/XI0_21/d__4_ xsel_21_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_3 XI11_6/XI0/XI0_21/d__3_ xsel_21_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_2 XI11_6/XI0/XI0_21/d__2_ xsel_21_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_1 XI11_6/XI0/XI0_21/d__1_ xsel_21_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_21/MN1_0 XI11_6/XI0/XI0_21/d__0_ xsel_21_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_15 XI11_6/net21_0_ xsel_20_ XI11_6/XI0/XI0_20/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_14 XI11_6/net21_1_ xsel_20_ XI11_6/XI0/XI0_20/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_13 XI11_6/net21_2_ xsel_20_ XI11_6/XI0/XI0_20/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_12 XI11_6/net21_3_ xsel_20_ XI11_6/XI0/XI0_20/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_11 XI11_6/net21_4_ xsel_20_ XI11_6/XI0/XI0_20/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_10 XI11_6/net21_5_ xsel_20_ XI11_6/XI0/XI0_20/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_9 XI11_6/net21_6_ xsel_20_ XI11_6/XI0/XI0_20/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_8 XI11_6/net21_7_ xsel_20_ XI11_6/XI0/XI0_20/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_7 XI11_6/net21_8_ xsel_20_ XI11_6/XI0/XI0_20/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_6 XI11_6/net21_9_ xsel_20_ XI11_6/XI0/XI0_20/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_5 XI11_6/net21_10_ xsel_20_ XI11_6/XI0/XI0_20/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_4 XI11_6/net21_11_ xsel_20_ XI11_6/XI0/XI0_20/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_3 XI11_6/net21_12_ xsel_20_ XI11_6/XI0/XI0_20/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_2 XI11_6/net21_13_ xsel_20_ XI11_6/XI0/XI0_20/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_1 XI11_6/net21_14_ xsel_20_ XI11_6/XI0/XI0_20/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN0_0 XI11_6/net21_15_ xsel_20_ XI11_6/XI0/XI0_20/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_15 XI11_6/XI0/XI0_20/d__15_ xsel_20_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_14 XI11_6/XI0/XI0_20/d__14_ xsel_20_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_13 XI11_6/XI0/XI0_20/d__13_ xsel_20_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_12 XI11_6/XI0/XI0_20/d__12_ xsel_20_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_11 XI11_6/XI0/XI0_20/d__11_ xsel_20_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_10 XI11_6/XI0/XI0_20/d__10_ xsel_20_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_9 XI11_6/XI0/XI0_20/d__9_ xsel_20_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_8 XI11_6/XI0/XI0_20/d__8_ xsel_20_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_7 XI11_6/XI0/XI0_20/d__7_ xsel_20_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_6 XI11_6/XI0/XI0_20/d__6_ xsel_20_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_5 XI11_6/XI0/XI0_20/d__5_ xsel_20_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_4 XI11_6/XI0/XI0_20/d__4_ xsel_20_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_3 XI11_6/XI0/XI0_20/d__3_ xsel_20_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_2 XI11_6/XI0/XI0_20/d__2_ xsel_20_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_1 XI11_6/XI0/XI0_20/d__1_ xsel_20_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_20/MN1_0 XI11_6/XI0/XI0_20/d__0_ xsel_20_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_15 XI11_6/net21_0_ xsel_19_ XI11_6/XI0/XI0_19/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_14 XI11_6/net21_1_ xsel_19_ XI11_6/XI0/XI0_19/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_13 XI11_6/net21_2_ xsel_19_ XI11_6/XI0/XI0_19/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_12 XI11_6/net21_3_ xsel_19_ XI11_6/XI0/XI0_19/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_11 XI11_6/net21_4_ xsel_19_ XI11_6/XI0/XI0_19/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_10 XI11_6/net21_5_ xsel_19_ XI11_6/XI0/XI0_19/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_9 XI11_6/net21_6_ xsel_19_ XI11_6/XI0/XI0_19/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_8 XI11_6/net21_7_ xsel_19_ XI11_6/XI0/XI0_19/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_7 XI11_6/net21_8_ xsel_19_ XI11_6/XI0/XI0_19/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_6 XI11_6/net21_9_ xsel_19_ XI11_6/XI0/XI0_19/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_5 XI11_6/net21_10_ xsel_19_ XI11_6/XI0/XI0_19/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_4 XI11_6/net21_11_ xsel_19_ XI11_6/XI0/XI0_19/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_3 XI11_6/net21_12_ xsel_19_ XI11_6/XI0/XI0_19/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_2 XI11_6/net21_13_ xsel_19_ XI11_6/XI0/XI0_19/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_1 XI11_6/net21_14_ xsel_19_ XI11_6/XI0/XI0_19/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN0_0 XI11_6/net21_15_ xsel_19_ XI11_6/XI0/XI0_19/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_15 XI11_6/XI0/XI0_19/d__15_ xsel_19_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_14 XI11_6/XI0/XI0_19/d__14_ xsel_19_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_13 XI11_6/XI0/XI0_19/d__13_ xsel_19_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_12 XI11_6/XI0/XI0_19/d__12_ xsel_19_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_11 XI11_6/XI0/XI0_19/d__11_ xsel_19_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_10 XI11_6/XI0/XI0_19/d__10_ xsel_19_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_9 XI11_6/XI0/XI0_19/d__9_ xsel_19_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_8 XI11_6/XI0/XI0_19/d__8_ xsel_19_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_7 XI11_6/XI0/XI0_19/d__7_ xsel_19_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_6 XI11_6/XI0/XI0_19/d__6_ xsel_19_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_5 XI11_6/XI0/XI0_19/d__5_ xsel_19_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_4 XI11_6/XI0/XI0_19/d__4_ xsel_19_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_3 XI11_6/XI0/XI0_19/d__3_ xsel_19_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_2 XI11_6/XI0/XI0_19/d__2_ xsel_19_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_1 XI11_6/XI0/XI0_19/d__1_ xsel_19_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_19/MN1_0 XI11_6/XI0/XI0_19/d__0_ xsel_19_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_15 XI11_6/net21_0_ xsel_18_ XI11_6/XI0/XI0_18/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_14 XI11_6/net21_1_ xsel_18_ XI11_6/XI0/XI0_18/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_13 XI11_6/net21_2_ xsel_18_ XI11_6/XI0/XI0_18/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_12 XI11_6/net21_3_ xsel_18_ XI11_6/XI0/XI0_18/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_11 XI11_6/net21_4_ xsel_18_ XI11_6/XI0/XI0_18/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_10 XI11_6/net21_5_ xsel_18_ XI11_6/XI0/XI0_18/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_9 XI11_6/net21_6_ xsel_18_ XI11_6/XI0/XI0_18/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_8 XI11_6/net21_7_ xsel_18_ XI11_6/XI0/XI0_18/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_7 XI11_6/net21_8_ xsel_18_ XI11_6/XI0/XI0_18/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_6 XI11_6/net21_9_ xsel_18_ XI11_6/XI0/XI0_18/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_5 XI11_6/net21_10_ xsel_18_ XI11_6/XI0/XI0_18/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_4 XI11_6/net21_11_ xsel_18_ XI11_6/XI0/XI0_18/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_3 XI11_6/net21_12_ xsel_18_ XI11_6/XI0/XI0_18/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_2 XI11_6/net21_13_ xsel_18_ XI11_6/XI0/XI0_18/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_1 XI11_6/net21_14_ xsel_18_ XI11_6/XI0/XI0_18/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN0_0 XI11_6/net21_15_ xsel_18_ XI11_6/XI0/XI0_18/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_15 XI11_6/XI0/XI0_18/d__15_ xsel_18_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_14 XI11_6/XI0/XI0_18/d__14_ xsel_18_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_13 XI11_6/XI0/XI0_18/d__13_ xsel_18_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_12 XI11_6/XI0/XI0_18/d__12_ xsel_18_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_11 XI11_6/XI0/XI0_18/d__11_ xsel_18_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_10 XI11_6/XI0/XI0_18/d__10_ xsel_18_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_9 XI11_6/XI0/XI0_18/d__9_ xsel_18_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_8 XI11_6/XI0/XI0_18/d__8_ xsel_18_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_7 XI11_6/XI0/XI0_18/d__7_ xsel_18_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_6 XI11_6/XI0/XI0_18/d__6_ xsel_18_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_5 XI11_6/XI0/XI0_18/d__5_ xsel_18_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_4 XI11_6/XI0/XI0_18/d__4_ xsel_18_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_3 XI11_6/XI0/XI0_18/d__3_ xsel_18_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_2 XI11_6/XI0/XI0_18/d__2_ xsel_18_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_1 XI11_6/XI0/XI0_18/d__1_ xsel_18_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_18/MN1_0 XI11_6/XI0/XI0_18/d__0_ xsel_18_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_15 XI11_6/net21_0_ xsel_17_ XI11_6/XI0/XI0_17/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_14 XI11_6/net21_1_ xsel_17_ XI11_6/XI0/XI0_17/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_13 XI11_6/net21_2_ xsel_17_ XI11_6/XI0/XI0_17/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_12 XI11_6/net21_3_ xsel_17_ XI11_6/XI0/XI0_17/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_11 XI11_6/net21_4_ xsel_17_ XI11_6/XI0/XI0_17/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_10 XI11_6/net21_5_ xsel_17_ XI11_6/XI0/XI0_17/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_9 XI11_6/net21_6_ xsel_17_ XI11_6/XI0/XI0_17/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_8 XI11_6/net21_7_ xsel_17_ XI11_6/XI0/XI0_17/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_7 XI11_6/net21_8_ xsel_17_ XI11_6/XI0/XI0_17/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_6 XI11_6/net21_9_ xsel_17_ XI11_6/XI0/XI0_17/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_5 XI11_6/net21_10_ xsel_17_ XI11_6/XI0/XI0_17/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_4 XI11_6/net21_11_ xsel_17_ XI11_6/XI0/XI0_17/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_3 XI11_6/net21_12_ xsel_17_ XI11_6/XI0/XI0_17/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_2 XI11_6/net21_13_ xsel_17_ XI11_6/XI0/XI0_17/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_1 XI11_6/net21_14_ xsel_17_ XI11_6/XI0/XI0_17/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN0_0 XI11_6/net21_15_ xsel_17_ XI11_6/XI0/XI0_17/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_15 XI11_6/XI0/XI0_17/d__15_ xsel_17_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_14 XI11_6/XI0/XI0_17/d__14_ xsel_17_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_13 XI11_6/XI0/XI0_17/d__13_ xsel_17_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_12 XI11_6/XI0/XI0_17/d__12_ xsel_17_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_11 XI11_6/XI0/XI0_17/d__11_ xsel_17_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_10 XI11_6/XI0/XI0_17/d__10_ xsel_17_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_9 XI11_6/XI0/XI0_17/d__9_ xsel_17_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_8 XI11_6/XI0/XI0_17/d__8_ xsel_17_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_7 XI11_6/XI0/XI0_17/d__7_ xsel_17_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_6 XI11_6/XI0/XI0_17/d__6_ xsel_17_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_5 XI11_6/XI0/XI0_17/d__5_ xsel_17_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_4 XI11_6/XI0/XI0_17/d__4_ xsel_17_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_3 XI11_6/XI0/XI0_17/d__3_ xsel_17_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_2 XI11_6/XI0/XI0_17/d__2_ xsel_17_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_1 XI11_6/XI0/XI0_17/d__1_ xsel_17_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_17/MN1_0 XI11_6/XI0/XI0_17/d__0_ xsel_17_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_15 XI11_6/net21_0_ xsel_16_ XI11_6/XI0/XI0_16/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_14 XI11_6/net21_1_ xsel_16_ XI11_6/XI0/XI0_16/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_13 XI11_6/net21_2_ xsel_16_ XI11_6/XI0/XI0_16/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_12 XI11_6/net21_3_ xsel_16_ XI11_6/XI0/XI0_16/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_11 XI11_6/net21_4_ xsel_16_ XI11_6/XI0/XI0_16/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_10 XI11_6/net21_5_ xsel_16_ XI11_6/XI0/XI0_16/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_9 XI11_6/net21_6_ xsel_16_ XI11_6/XI0/XI0_16/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_8 XI11_6/net21_7_ xsel_16_ XI11_6/XI0/XI0_16/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_7 XI11_6/net21_8_ xsel_16_ XI11_6/XI0/XI0_16/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_6 XI11_6/net21_9_ xsel_16_ XI11_6/XI0/XI0_16/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_5 XI11_6/net21_10_ xsel_16_ XI11_6/XI0/XI0_16/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_4 XI11_6/net21_11_ xsel_16_ XI11_6/XI0/XI0_16/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_3 XI11_6/net21_12_ xsel_16_ XI11_6/XI0/XI0_16/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_2 XI11_6/net21_13_ xsel_16_ XI11_6/XI0/XI0_16/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_1 XI11_6/net21_14_ xsel_16_ XI11_6/XI0/XI0_16/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN0_0 XI11_6/net21_15_ xsel_16_ XI11_6/XI0/XI0_16/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_15 XI11_6/XI0/XI0_16/d__15_ xsel_16_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_14 XI11_6/XI0/XI0_16/d__14_ xsel_16_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_13 XI11_6/XI0/XI0_16/d__13_ xsel_16_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_12 XI11_6/XI0/XI0_16/d__12_ xsel_16_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_11 XI11_6/XI0/XI0_16/d__11_ xsel_16_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_10 XI11_6/XI0/XI0_16/d__10_ xsel_16_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_9 XI11_6/XI0/XI0_16/d__9_ xsel_16_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_8 XI11_6/XI0/XI0_16/d__8_ xsel_16_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_7 XI11_6/XI0/XI0_16/d__7_ xsel_16_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_6 XI11_6/XI0/XI0_16/d__6_ xsel_16_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_5 XI11_6/XI0/XI0_16/d__5_ xsel_16_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_4 XI11_6/XI0/XI0_16/d__4_ xsel_16_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_3 XI11_6/XI0/XI0_16/d__3_ xsel_16_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_2 XI11_6/XI0/XI0_16/d__2_ xsel_16_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_1 XI11_6/XI0/XI0_16/d__1_ xsel_16_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_16/MN1_0 XI11_6/XI0/XI0_16/d__0_ xsel_16_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_15 XI11_6/net21_0_ xsel_15_ XI11_6/XI0/XI0_15/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_14 XI11_6/net21_1_ xsel_15_ XI11_6/XI0/XI0_15/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_13 XI11_6/net21_2_ xsel_15_ XI11_6/XI0/XI0_15/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_12 XI11_6/net21_3_ xsel_15_ XI11_6/XI0/XI0_15/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_11 XI11_6/net21_4_ xsel_15_ XI11_6/XI0/XI0_15/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_10 XI11_6/net21_5_ xsel_15_ XI11_6/XI0/XI0_15/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_9 XI11_6/net21_6_ xsel_15_ XI11_6/XI0/XI0_15/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_8 XI11_6/net21_7_ xsel_15_ XI11_6/XI0/XI0_15/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_7 XI11_6/net21_8_ xsel_15_ XI11_6/XI0/XI0_15/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_6 XI11_6/net21_9_ xsel_15_ XI11_6/XI0/XI0_15/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_5 XI11_6/net21_10_ xsel_15_ XI11_6/XI0/XI0_15/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_4 XI11_6/net21_11_ xsel_15_ XI11_6/XI0/XI0_15/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_3 XI11_6/net21_12_ xsel_15_ XI11_6/XI0/XI0_15/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_2 XI11_6/net21_13_ xsel_15_ XI11_6/XI0/XI0_15/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_1 XI11_6/net21_14_ xsel_15_ XI11_6/XI0/XI0_15/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN0_0 XI11_6/net21_15_ xsel_15_ XI11_6/XI0/XI0_15/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_15 XI11_6/XI0/XI0_15/d__15_ xsel_15_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_14 XI11_6/XI0/XI0_15/d__14_ xsel_15_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_13 XI11_6/XI0/XI0_15/d__13_ xsel_15_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_12 XI11_6/XI0/XI0_15/d__12_ xsel_15_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_11 XI11_6/XI0/XI0_15/d__11_ xsel_15_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_10 XI11_6/XI0/XI0_15/d__10_ xsel_15_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_9 XI11_6/XI0/XI0_15/d__9_ xsel_15_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_8 XI11_6/XI0/XI0_15/d__8_ xsel_15_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_7 XI11_6/XI0/XI0_15/d__7_ xsel_15_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_6 XI11_6/XI0/XI0_15/d__6_ xsel_15_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_5 XI11_6/XI0/XI0_15/d__5_ xsel_15_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_4 XI11_6/XI0/XI0_15/d__4_ xsel_15_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_3 XI11_6/XI0/XI0_15/d__3_ xsel_15_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_2 XI11_6/XI0/XI0_15/d__2_ xsel_15_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_1 XI11_6/XI0/XI0_15/d__1_ xsel_15_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_15/MN1_0 XI11_6/XI0/XI0_15/d__0_ xsel_15_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_15 XI11_6/net21_0_ xsel_14_ XI11_6/XI0/XI0_14/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_14 XI11_6/net21_1_ xsel_14_ XI11_6/XI0/XI0_14/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_13 XI11_6/net21_2_ xsel_14_ XI11_6/XI0/XI0_14/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_12 XI11_6/net21_3_ xsel_14_ XI11_6/XI0/XI0_14/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_11 XI11_6/net21_4_ xsel_14_ XI11_6/XI0/XI0_14/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_10 XI11_6/net21_5_ xsel_14_ XI11_6/XI0/XI0_14/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_9 XI11_6/net21_6_ xsel_14_ XI11_6/XI0/XI0_14/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_8 XI11_6/net21_7_ xsel_14_ XI11_6/XI0/XI0_14/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_7 XI11_6/net21_8_ xsel_14_ XI11_6/XI0/XI0_14/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_6 XI11_6/net21_9_ xsel_14_ XI11_6/XI0/XI0_14/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_5 XI11_6/net21_10_ xsel_14_ XI11_6/XI0/XI0_14/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_4 XI11_6/net21_11_ xsel_14_ XI11_6/XI0/XI0_14/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_3 XI11_6/net21_12_ xsel_14_ XI11_6/XI0/XI0_14/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_2 XI11_6/net21_13_ xsel_14_ XI11_6/XI0/XI0_14/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_1 XI11_6/net21_14_ xsel_14_ XI11_6/XI0/XI0_14/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN0_0 XI11_6/net21_15_ xsel_14_ XI11_6/XI0/XI0_14/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_15 XI11_6/XI0/XI0_14/d__15_ xsel_14_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_14 XI11_6/XI0/XI0_14/d__14_ xsel_14_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_13 XI11_6/XI0/XI0_14/d__13_ xsel_14_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_12 XI11_6/XI0/XI0_14/d__12_ xsel_14_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_11 XI11_6/XI0/XI0_14/d__11_ xsel_14_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_10 XI11_6/XI0/XI0_14/d__10_ xsel_14_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_9 XI11_6/XI0/XI0_14/d__9_ xsel_14_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_8 XI11_6/XI0/XI0_14/d__8_ xsel_14_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_7 XI11_6/XI0/XI0_14/d__7_ xsel_14_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_6 XI11_6/XI0/XI0_14/d__6_ xsel_14_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_5 XI11_6/XI0/XI0_14/d__5_ xsel_14_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_4 XI11_6/XI0/XI0_14/d__4_ xsel_14_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_3 XI11_6/XI0/XI0_14/d__3_ xsel_14_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_2 XI11_6/XI0/XI0_14/d__2_ xsel_14_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_1 XI11_6/XI0/XI0_14/d__1_ xsel_14_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_14/MN1_0 XI11_6/XI0/XI0_14/d__0_ xsel_14_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_15 XI11_6/net21_0_ xsel_13_ XI11_6/XI0/XI0_13/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_14 XI11_6/net21_1_ xsel_13_ XI11_6/XI0/XI0_13/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_13 XI11_6/net21_2_ xsel_13_ XI11_6/XI0/XI0_13/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_12 XI11_6/net21_3_ xsel_13_ XI11_6/XI0/XI0_13/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_11 XI11_6/net21_4_ xsel_13_ XI11_6/XI0/XI0_13/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_10 XI11_6/net21_5_ xsel_13_ XI11_6/XI0/XI0_13/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_9 XI11_6/net21_6_ xsel_13_ XI11_6/XI0/XI0_13/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_8 XI11_6/net21_7_ xsel_13_ XI11_6/XI0/XI0_13/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_7 XI11_6/net21_8_ xsel_13_ XI11_6/XI0/XI0_13/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_6 XI11_6/net21_9_ xsel_13_ XI11_6/XI0/XI0_13/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_5 XI11_6/net21_10_ xsel_13_ XI11_6/XI0/XI0_13/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_4 XI11_6/net21_11_ xsel_13_ XI11_6/XI0/XI0_13/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_3 XI11_6/net21_12_ xsel_13_ XI11_6/XI0/XI0_13/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_2 XI11_6/net21_13_ xsel_13_ XI11_6/XI0/XI0_13/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_1 XI11_6/net21_14_ xsel_13_ XI11_6/XI0/XI0_13/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN0_0 XI11_6/net21_15_ xsel_13_ XI11_6/XI0/XI0_13/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_15 XI11_6/XI0/XI0_13/d__15_ xsel_13_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_14 XI11_6/XI0/XI0_13/d__14_ xsel_13_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_13 XI11_6/XI0/XI0_13/d__13_ xsel_13_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_12 XI11_6/XI0/XI0_13/d__12_ xsel_13_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_11 XI11_6/XI0/XI0_13/d__11_ xsel_13_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_10 XI11_6/XI0/XI0_13/d__10_ xsel_13_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_9 XI11_6/XI0/XI0_13/d__9_ xsel_13_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_8 XI11_6/XI0/XI0_13/d__8_ xsel_13_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_7 XI11_6/XI0/XI0_13/d__7_ xsel_13_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_6 XI11_6/XI0/XI0_13/d__6_ xsel_13_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_5 XI11_6/XI0/XI0_13/d__5_ xsel_13_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_4 XI11_6/XI0/XI0_13/d__4_ xsel_13_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_3 XI11_6/XI0/XI0_13/d__3_ xsel_13_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_2 XI11_6/XI0/XI0_13/d__2_ xsel_13_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_1 XI11_6/XI0/XI0_13/d__1_ xsel_13_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_13/MN1_0 XI11_6/XI0/XI0_13/d__0_ xsel_13_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_15 XI11_6/net21_0_ xsel_12_ XI11_6/XI0/XI0_12/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_14 XI11_6/net21_1_ xsel_12_ XI11_6/XI0/XI0_12/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_13 XI11_6/net21_2_ xsel_12_ XI11_6/XI0/XI0_12/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_12 XI11_6/net21_3_ xsel_12_ XI11_6/XI0/XI0_12/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_11 XI11_6/net21_4_ xsel_12_ XI11_6/XI0/XI0_12/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_10 XI11_6/net21_5_ xsel_12_ XI11_6/XI0/XI0_12/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_9 XI11_6/net21_6_ xsel_12_ XI11_6/XI0/XI0_12/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_8 XI11_6/net21_7_ xsel_12_ XI11_6/XI0/XI0_12/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_7 XI11_6/net21_8_ xsel_12_ XI11_6/XI0/XI0_12/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_6 XI11_6/net21_9_ xsel_12_ XI11_6/XI0/XI0_12/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_5 XI11_6/net21_10_ xsel_12_ XI11_6/XI0/XI0_12/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_4 XI11_6/net21_11_ xsel_12_ XI11_6/XI0/XI0_12/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_3 XI11_6/net21_12_ xsel_12_ XI11_6/XI0/XI0_12/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_2 XI11_6/net21_13_ xsel_12_ XI11_6/XI0/XI0_12/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_1 XI11_6/net21_14_ xsel_12_ XI11_6/XI0/XI0_12/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN0_0 XI11_6/net21_15_ xsel_12_ XI11_6/XI0/XI0_12/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_15 XI11_6/XI0/XI0_12/d__15_ xsel_12_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_14 XI11_6/XI0/XI0_12/d__14_ xsel_12_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_13 XI11_6/XI0/XI0_12/d__13_ xsel_12_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_12 XI11_6/XI0/XI0_12/d__12_ xsel_12_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_11 XI11_6/XI0/XI0_12/d__11_ xsel_12_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_10 XI11_6/XI0/XI0_12/d__10_ xsel_12_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_9 XI11_6/XI0/XI0_12/d__9_ xsel_12_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_8 XI11_6/XI0/XI0_12/d__8_ xsel_12_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_7 XI11_6/XI0/XI0_12/d__7_ xsel_12_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_6 XI11_6/XI0/XI0_12/d__6_ xsel_12_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_5 XI11_6/XI0/XI0_12/d__5_ xsel_12_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_4 XI11_6/XI0/XI0_12/d__4_ xsel_12_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_3 XI11_6/XI0/XI0_12/d__3_ xsel_12_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_2 XI11_6/XI0/XI0_12/d__2_ xsel_12_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_1 XI11_6/XI0/XI0_12/d__1_ xsel_12_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_12/MN1_0 XI11_6/XI0/XI0_12/d__0_ xsel_12_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_15 XI11_6/net21_0_ xsel_11_ XI11_6/XI0/XI0_11/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_14 XI11_6/net21_1_ xsel_11_ XI11_6/XI0/XI0_11/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_13 XI11_6/net21_2_ xsel_11_ XI11_6/XI0/XI0_11/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_12 XI11_6/net21_3_ xsel_11_ XI11_6/XI0/XI0_11/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_11 XI11_6/net21_4_ xsel_11_ XI11_6/XI0/XI0_11/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_10 XI11_6/net21_5_ xsel_11_ XI11_6/XI0/XI0_11/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_9 XI11_6/net21_6_ xsel_11_ XI11_6/XI0/XI0_11/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_8 XI11_6/net21_7_ xsel_11_ XI11_6/XI0/XI0_11/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_7 XI11_6/net21_8_ xsel_11_ XI11_6/XI0/XI0_11/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_6 XI11_6/net21_9_ xsel_11_ XI11_6/XI0/XI0_11/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_5 XI11_6/net21_10_ xsel_11_ XI11_6/XI0/XI0_11/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_4 XI11_6/net21_11_ xsel_11_ XI11_6/XI0/XI0_11/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_3 XI11_6/net21_12_ xsel_11_ XI11_6/XI0/XI0_11/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_2 XI11_6/net21_13_ xsel_11_ XI11_6/XI0/XI0_11/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_1 XI11_6/net21_14_ xsel_11_ XI11_6/XI0/XI0_11/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN0_0 XI11_6/net21_15_ xsel_11_ XI11_6/XI0/XI0_11/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_15 XI11_6/XI0/XI0_11/d__15_ xsel_11_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_14 XI11_6/XI0/XI0_11/d__14_ xsel_11_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_13 XI11_6/XI0/XI0_11/d__13_ xsel_11_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_12 XI11_6/XI0/XI0_11/d__12_ xsel_11_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_11 XI11_6/XI0/XI0_11/d__11_ xsel_11_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_10 XI11_6/XI0/XI0_11/d__10_ xsel_11_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_9 XI11_6/XI0/XI0_11/d__9_ xsel_11_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_8 XI11_6/XI0/XI0_11/d__8_ xsel_11_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_7 XI11_6/XI0/XI0_11/d__7_ xsel_11_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_6 XI11_6/XI0/XI0_11/d__6_ xsel_11_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_5 XI11_6/XI0/XI0_11/d__5_ xsel_11_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_4 XI11_6/XI0/XI0_11/d__4_ xsel_11_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_3 XI11_6/XI0/XI0_11/d__3_ xsel_11_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_2 XI11_6/XI0/XI0_11/d__2_ xsel_11_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_1 XI11_6/XI0/XI0_11/d__1_ xsel_11_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_11/MN1_0 XI11_6/XI0/XI0_11/d__0_ xsel_11_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_15 XI11_6/net21_0_ xsel_10_ XI11_6/XI0/XI0_10/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_14 XI11_6/net21_1_ xsel_10_ XI11_6/XI0/XI0_10/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_13 XI11_6/net21_2_ xsel_10_ XI11_6/XI0/XI0_10/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_12 XI11_6/net21_3_ xsel_10_ XI11_6/XI0/XI0_10/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_11 XI11_6/net21_4_ xsel_10_ XI11_6/XI0/XI0_10/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_10 XI11_6/net21_5_ xsel_10_ XI11_6/XI0/XI0_10/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_9 XI11_6/net21_6_ xsel_10_ XI11_6/XI0/XI0_10/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_8 XI11_6/net21_7_ xsel_10_ XI11_6/XI0/XI0_10/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_7 XI11_6/net21_8_ xsel_10_ XI11_6/XI0/XI0_10/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_6 XI11_6/net21_9_ xsel_10_ XI11_6/XI0/XI0_10/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_5 XI11_6/net21_10_ xsel_10_ XI11_6/XI0/XI0_10/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_4 XI11_6/net21_11_ xsel_10_ XI11_6/XI0/XI0_10/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_3 XI11_6/net21_12_ xsel_10_ XI11_6/XI0/XI0_10/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_2 XI11_6/net21_13_ xsel_10_ XI11_6/XI0/XI0_10/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_1 XI11_6/net21_14_ xsel_10_ XI11_6/XI0/XI0_10/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN0_0 XI11_6/net21_15_ xsel_10_ XI11_6/XI0/XI0_10/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_15 XI11_6/XI0/XI0_10/d__15_ xsel_10_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_14 XI11_6/XI0/XI0_10/d__14_ xsel_10_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_13 XI11_6/XI0/XI0_10/d__13_ xsel_10_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_12 XI11_6/XI0/XI0_10/d__12_ xsel_10_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_11 XI11_6/XI0/XI0_10/d__11_ xsel_10_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_10 XI11_6/XI0/XI0_10/d__10_ xsel_10_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_9 XI11_6/XI0/XI0_10/d__9_ xsel_10_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_8 XI11_6/XI0/XI0_10/d__8_ xsel_10_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_7 XI11_6/XI0/XI0_10/d__7_ xsel_10_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_6 XI11_6/XI0/XI0_10/d__6_ xsel_10_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_5 XI11_6/XI0/XI0_10/d__5_ xsel_10_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_4 XI11_6/XI0/XI0_10/d__4_ xsel_10_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_3 XI11_6/XI0/XI0_10/d__3_ xsel_10_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_2 XI11_6/XI0/XI0_10/d__2_ xsel_10_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_1 XI11_6/XI0/XI0_10/d__1_ xsel_10_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_10/MN1_0 XI11_6/XI0/XI0_10/d__0_ xsel_10_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_15 XI11_6/net21_0_ xsel_9_ XI11_6/XI0/XI0_9/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_14 XI11_6/net21_1_ xsel_9_ XI11_6/XI0/XI0_9/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_13 XI11_6/net21_2_ xsel_9_ XI11_6/XI0/XI0_9/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_12 XI11_6/net21_3_ xsel_9_ XI11_6/XI0/XI0_9/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_11 XI11_6/net21_4_ xsel_9_ XI11_6/XI0/XI0_9/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_10 XI11_6/net21_5_ xsel_9_ XI11_6/XI0/XI0_9/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_9 XI11_6/net21_6_ xsel_9_ XI11_6/XI0/XI0_9/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_8 XI11_6/net21_7_ xsel_9_ XI11_6/XI0/XI0_9/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_7 XI11_6/net21_8_ xsel_9_ XI11_6/XI0/XI0_9/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_6 XI11_6/net21_9_ xsel_9_ XI11_6/XI0/XI0_9/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_5 XI11_6/net21_10_ xsel_9_ XI11_6/XI0/XI0_9/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_4 XI11_6/net21_11_ xsel_9_ XI11_6/XI0/XI0_9/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_3 XI11_6/net21_12_ xsel_9_ XI11_6/XI0/XI0_9/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_2 XI11_6/net21_13_ xsel_9_ XI11_6/XI0/XI0_9/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_1 XI11_6/net21_14_ xsel_9_ XI11_6/XI0/XI0_9/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN0_0 XI11_6/net21_15_ xsel_9_ XI11_6/XI0/XI0_9/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_15 XI11_6/XI0/XI0_9/d__15_ xsel_9_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_14 XI11_6/XI0/XI0_9/d__14_ xsel_9_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_13 XI11_6/XI0/XI0_9/d__13_ xsel_9_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_12 XI11_6/XI0/XI0_9/d__12_ xsel_9_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_11 XI11_6/XI0/XI0_9/d__11_ xsel_9_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_10 XI11_6/XI0/XI0_9/d__10_ xsel_9_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_9 XI11_6/XI0/XI0_9/d__9_ xsel_9_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_8 XI11_6/XI0/XI0_9/d__8_ xsel_9_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_7 XI11_6/XI0/XI0_9/d__7_ xsel_9_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_6 XI11_6/XI0/XI0_9/d__6_ xsel_9_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_5 XI11_6/XI0/XI0_9/d__5_ xsel_9_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_4 XI11_6/XI0/XI0_9/d__4_ xsel_9_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_3 XI11_6/XI0/XI0_9/d__3_ xsel_9_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_2 XI11_6/XI0/XI0_9/d__2_ xsel_9_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_1 XI11_6/XI0/XI0_9/d__1_ xsel_9_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_9/MN1_0 XI11_6/XI0/XI0_9/d__0_ xsel_9_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_15 XI11_6/net21_0_ xsel_8_ XI11_6/XI0/XI0_8/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_14 XI11_6/net21_1_ xsel_8_ XI11_6/XI0/XI0_8/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_13 XI11_6/net21_2_ xsel_8_ XI11_6/XI0/XI0_8/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_12 XI11_6/net21_3_ xsel_8_ XI11_6/XI0/XI0_8/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_11 XI11_6/net21_4_ xsel_8_ XI11_6/XI0/XI0_8/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_10 XI11_6/net21_5_ xsel_8_ XI11_6/XI0/XI0_8/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_9 XI11_6/net21_6_ xsel_8_ XI11_6/XI0/XI0_8/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_8 XI11_6/net21_7_ xsel_8_ XI11_6/XI0/XI0_8/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_7 XI11_6/net21_8_ xsel_8_ XI11_6/XI0/XI0_8/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_6 XI11_6/net21_9_ xsel_8_ XI11_6/XI0/XI0_8/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_5 XI11_6/net21_10_ xsel_8_ XI11_6/XI0/XI0_8/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_4 XI11_6/net21_11_ xsel_8_ XI11_6/XI0/XI0_8/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_3 XI11_6/net21_12_ xsel_8_ XI11_6/XI0/XI0_8/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_2 XI11_6/net21_13_ xsel_8_ XI11_6/XI0/XI0_8/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_1 XI11_6/net21_14_ xsel_8_ XI11_6/XI0/XI0_8/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN0_0 XI11_6/net21_15_ xsel_8_ XI11_6/XI0/XI0_8/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_15 XI11_6/XI0/XI0_8/d__15_ xsel_8_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_14 XI11_6/XI0/XI0_8/d__14_ xsel_8_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_13 XI11_6/XI0/XI0_8/d__13_ xsel_8_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_12 XI11_6/XI0/XI0_8/d__12_ xsel_8_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_11 XI11_6/XI0/XI0_8/d__11_ xsel_8_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_10 XI11_6/XI0/XI0_8/d__10_ xsel_8_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_9 XI11_6/XI0/XI0_8/d__9_ xsel_8_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_8 XI11_6/XI0/XI0_8/d__8_ xsel_8_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_7 XI11_6/XI0/XI0_8/d__7_ xsel_8_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_6 XI11_6/XI0/XI0_8/d__6_ xsel_8_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_5 XI11_6/XI0/XI0_8/d__5_ xsel_8_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_4 XI11_6/XI0/XI0_8/d__4_ xsel_8_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_3 XI11_6/XI0/XI0_8/d__3_ xsel_8_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_2 XI11_6/XI0/XI0_8/d__2_ xsel_8_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_1 XI11_6/XI0/XI0_8/d__1_ xsel_8_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_8/MN1_0 XI11_6/XI0/XI0_8/d__0_ xsel_8_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_15 XI11_6/net21_0_ xsel_7_ XI11_6/XI0/XI0_7/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_14 XI11_6/net21_1_ xsel_7_ XI11_6/XI0/XI0_7/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_13 XI11_6/net21_2_ xsel_7_ XI11_6/XI0/XI0_7/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_12 XI11_6/net21_3_ xsel_7_ XI11_6/XI0/XI0_7/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_11 XI11_6/net21_4_ xsel_7_ XI11_6/XI0/XI0_7/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_10 XI11_6/net21_5_ xsel_7_ XI11_6/XI0/XI0_7/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_9 XI11_6/net21_6_ xsel_7_ XI11_6/XI0/XI0_7/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_8 XI11_6/net21_7_ xsel_7_ XI11_6/XI0/XI0_7/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_7 XI11_6/net21_8_ xsel_7_ XI11_6/XI0/XI0_7/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_6 XI11_6/net21_9_ xsel_7_ XI11_6/XI0/XI0_7/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_5 XI11_6/net21_10_ xsel_7_ XI11_6/XI0/XI0_7/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_4 XI11_6/net21_11_ xsel_7_ XI11_6/XI0/XI0_7/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_3 XI11_6/net21_12_ xsel_7_ XI11_6/XI0/XI0_7/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_2 XI11_6/net21_13_ xsel_7_ XI11_6/XI0/XI0_7/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_1 XI11_6/net21_14_ xsel_7_ XI11_6/XI0/XI0_7/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN0_0 XI11_6/net21_15_ xsel_7_ XI11_6/XI0/XI0_7/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_15 XI11_6/XI0/XI0_7/d__15_ xsel_7_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_14 XI11_6/XI0/XI0_7/d__14_ xsel_7_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_13 XI11_6/XI0/XI0_7/d__13_ xsel_7_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_12 XI11_6/XI0/XI0_7/d__12_ xsel_7_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_11 XI11_6/XI0/XI0_7/d__11_ xsel_7_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_10 XI11_6/XI0/XI0_7/d__10_ xsel_7_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_9 XI11_6/XI0/XI0_7/d__9_ xsel_7_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_8 XI11_6/XI0/XI0_7/d__8_ xsel_7_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_7 XI11_6/XI0/XI0_7/d__7_ xsel_7_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_6 XI11_6/XI0/XI0_7/d__6_ xsel_7_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_5 XI11_6/XI0/XI0_7/d__5_ xsel_7_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_4 XI11_6/XI0/XI0_7/d__4_ xsel_7_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_3 XI11_6/XI0/XI0_7/d__3_ xsel_7_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_2 XI11_6/XI0/XI0_7/d__2_ xsel_7_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_1 XI11_6/XI0/XI0_7/d__1_ xsel_7_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_7/MN1_0 XI11_6/XI0/XI0_7/d__0_ xsel_7_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_15 XI11_6/net21_0_ xsel_6_ XI11_6/XI0/XI0_6/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_14 XI11_6/net21_1_ xsel_6_ XI11_6/XI0/XI0_6/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_13 XI11_6/net21_2_ xsel_6_ XI11_6/XI0/XI0_6/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_12 XI11_6/net21_3_ xsel_6_ XI11_6/XI0/XI0_6/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_11 XI11_6/net21_4_ xsel_6_ XI11_6/XI0/XI0_6/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_10 XI11_6/net21_5_ xsel_6_ XI11_6/XI0/XI0_6/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_9 XI11_6/net21_6_ xsel_6_ XI11_6/XI0/XI0_6/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_8 XI11_6/net21_7_ xsel_6_ XI11_6/XI0/XI0_6/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_7 XI11_6/net21_8_ xsel_6_ XI11_6/XI0/XI0_6/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_6 XI11_6/net21_9_ xsel_6_ XI11_6/XI0/XI0_6/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_5 XI11_6/net21_10_ xsel_6_ XI11_6/XI0/XI0_6/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_4 XI11_6/net21_11_ xsel_6_ XI11_6/XI0/XI0_6/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_3 XI11_6/net21_12_ xsel_6_ XI11_6/XI0/XI0_6/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_2 XI11_6/net21_13_ xsel_6_ XI11_6/XI0/XI0_6/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_1 XI11_6/net21_14_ xsel_6_ XI11_6/XI0/XI0_6/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN0_0 XI11_6/net21_15_ xsel_6_ XI11_6/XI0/XI0_6/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_15 XI11_6/XI0/XI0_6/d__15_ xsel_6_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_14 XI11_6/XI0/XI0_6/d__14_ xsel_6_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_13 XI11_6/XI0/XI0_6/d__13_ xsel_6_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_12 XI11_6/XI0/XI0_6/d__12_ xsel_6_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_11 XI11_6/XI0/XI0_6/d__11_ xsel_6_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_10 XI11_6/XI0/XI0_6/d__10_ xsel_6_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_9 XI11_6/XI0/XI0_6/d__9_ xsel_6_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_8 XI11_6/XI0/XI0_6/d__8_ xsel_6_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_7 XI11_6/XI0/XI0_6/d__7_ xsel_6_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_6 XI11_6/XI0/XI0_6/d__6_ xsel_6_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_5 XI11_6/XI0/XI0_6/d__5_ xsel_6_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_4 XI11_6/XI0/XI0_6/d__4_ xsel_6_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_3 XI11_6/XI0/XI0_6/d__3_ xsel_6_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_2 XI11_6/XI0/XI0_6/d__2_ xsel_6_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_1 XI11_6/XI0/XI0_6/d__1_ xsel_6_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_6/MN1_0 XI11_6/XI0/XI0_6/d__0_ xsel_6_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_15 XI11_6/net21_0_ xsel_5_ XI11_6/XI0/XI0_5/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_14 XI11_6/net21_1_ xsel_5_ XI11_6/XI0/XI0_5/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_13 XI11_6/net21_2_ xsel_5_ XI11_6/XI0/XI0_5/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_12 XI11_6/net21_3_ xsel_5_ XI11_6/XI0/XI0_5/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_11 XI11_6/net21_4_ xsel_5_ XI11_6/XI0/XI0_5/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_10 XI11_6/net21_5_ xsel_5_ XI11_6/XI0/XI0_5/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_9 XI11_6/net21_6_ xsel_5_ XI11_6/XI0/XI0_5/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_8 XI11_6/net21_7_ xsel_5_ XI11_6/XI0/XI0_5/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_7 XI11_6/net21_8_ xsel_5_ XI11_6/XI0/XI0_5/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_6 XI11_6/net21_9_ xsel_5_ XI11_6/XI0/XI0_5/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_5 XI11_6/net21_10_ xsel_5_ XI11_6/XI0/XI0_5/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_4 XI11_6/net21_11_ xsel_5_ XI11_6/XI0/XI0_5/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_3 XI11_6/net21_12_ xsel_5_ XI11_6/XI0/XI0_5/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_2 XI11_6/net21_13_ xsel_5_ XI11_6/XI0/XI0_5/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_1 XI11_6/net21_14_ xsel_5_ XI11_6/XI0/XI0_5/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN0_0 XI11_6/net21_15_ xsel_5_ XI11_6/XI0/XI0_5/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_15 XI11_6/XI0/XI0_5/d__15_ xsel_5_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_14 XI11_6/XI0/XI0_5/d__14_ xsel_5_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_13 XI11_6/XI0/XI0_5/d__13_ xsel_5_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_12 XI11_6/XI0/XI0_5/d__12_ xsel_5_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_11 XI11_6/XI0/XI0_5/d__11_ xsel_5_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_10 XI11_6/XI0/XI0_5/d__10_ xsel_5_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_9 XI11_6/XI0/XI0_5/d__9_ xsel_5_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_8 XI11_6/XI0/XI0_5/d__8_ xsel_5_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_7 XI11_6/XI0/XI0_5/d__7_ xsel_5_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_6 XI11_6/XI0/XI0_5/d__6_ xsel_5_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_5 XI11_6/XI0/XI0_5/d__5_ xsel_5_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_4 XI11_6/XI0/XI0_5/d__4_ xsel_5_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_3 XI11_6/XI0/XI0_5/d__3_ xsel_5_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_2 XI11_6/XI0/XI0_5/d__2_ xsel_5_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_1 XI11_6/XI0/XI0_5/d__1_ xsel_5_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_5/MN1_0 XI11_6/XI0/XI0_5/d__0_ xsel_5_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_15 XI11_6/net21_0_ xsel_4_ XI11_6/XI0/XI0_4/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_14 XI11_6/net21_1_ xsel_4_ XI11_6/XI0/XI0_4/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_13 XI11_6/net21_2_ xsel_4_ XI11_6/XI0/XI0_4/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_12 XI11_6/net21_3_ xsel_4_ XI11_6/XI0/XI0_4/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_11 XI11_6/net21_4_ xsel_4_ XI11_6/XI0/XI0_4/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_10 XI11_6/net21_5_ xsel_4_ XI11_6/XI0/XI0_4/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_9 XI11_6/net21_6_ xsel_4_ XI11_6/XI0/XI0_4/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_8 XI11_6/net21_7_ xsel_4_ XI11_6/XI0/XI0_4/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_7 XI11_6/net21_8_ xsel_4_ XI11_6/XI0/XI0_4/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_6 XI11_6/net21_9_ xsel_4_ XI11_6/XI0/XI0_4/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_5 XI11_6/net21_10_ xsel_4_ XI11_6/XI0/XI0_4/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_4 XI11_6/net21_11_ xsel_4_ XI11_6/XI0/XI0_4/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_3 XI11_6/net21_12_ xsel_4_ XI11_6/XI0/XI0_4/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_2 XI11_6/net21_13_ xsel_4_ XI11_6/XI0/XI0_4/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_1 XI11_6/net21_14_ xsel_4_ XI11_6/XI0/XI0_4/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN0_0 XI11_6/net21_15_ xsel_4_ XI11_6/XI0/XI0_4/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_15 XI11_6/XI0/XI0_4/d__15_ xsel_4_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_14 XI11_6/XI0/XI0_4/d__14_ xsel_4_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_13 XI11_6/XI0/XI0_4/d__13_ xsel_4_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_12 XI11_6/XI0/XI0_4/d__12_ xsel_4_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_11 XI11_6/XI0/XI0_4/d__11_ xsel_4_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_10 XI11_6/XI0/XI0_4/d__10_ xsel_4_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_9 XI11_6/XI0/XI0_4/d__9_ xsel_4_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_8 XI11_6/XI0/XI0_4/d__8_ xsel_4_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_7 XI11_6/XI0/XI0_4/d__7_ xsel_4_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_6 XI11_6/XI0/XI0_4/d__6_ xsel_4_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_5 XI11_6/XI0/XI0_4/d__5_ xsel_4_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_4 XI11_6/XI0/XI0_4/d__4_ xsel_4_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_3 XI11_6/XI0/XI0_4/d__3_ xsel_4_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_2 XI11_6/XI0/XI0_4/d__2_ xsel_4_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_1 XI11_6/XI0/XI0_4/d__1_ xsel_4_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_4/MN1_0 XI11_6/XI0/XI0_4/d__0_ xsel_4_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_15 XI11_6/net21_0_ xsel_3_ XI11_6/XI0/XI0_3/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_14 XI11_6/net21_1_ xsel_3_ XI11_6/XI0/XI0_3/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_13 XI11_6/net21_2_ xsel_3_ XI11_6/XI0/XI0_3/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_12 XI11_6/net21_3_ xsel_3_ XI11_6/XI0/XI0_3/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_11 XI11_6/net21_4_ xsel_3_ XI11_6/XI0/XI0_3/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_10 XI11_6/net21_5_ xsel_3_ XI11_6/XI0/XI0_3/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_9 XI11_6/net21_6_ xsel_3_ XI11_6/XI0/XI0_3/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_8 XI11_6/net21_7_ xsel_3_ XI11_6/XI0/XI0_3/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_7 XI11_6/net21_8_ xsel_3_ XI11_6/XI0/XI0_3/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_6 XI11_6/net21_9_ xsel_3_ XI11_6/XI0/XI0_3/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_5 XI11_6/net21_10_ xsel_3_ XI11_6/XI0/XI0_3/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_4 XI11_6/net21_11_ xsel_3_ XI11_6/XI0/XI0_3/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_3 XI11_6/net21_12_ xsel_3_ XI11_6/XI0/XI0_3/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_2 XI11_6/net21_13_ xsel_3_ XI11_6/XI0/XI0_3/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_1 XI11_6/net21_14_ xsel_3_ XI11_6/XI0/XI0_3/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN0_0 XI11_6/net21_15_ xsel_3_ XI11_6/XI0/XI0_3/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_15 XI11_6/XI0/XI0_3/d__15_ xsel_3_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_14 XI11_6/XI0/XI0_3/d__14_ xsel_3_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_13 XI11_6/XI0/XI0_3/d__13_ xsel_3_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_12 XI11_6/XI0/XI0_3/d__12_ xsel_3_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_11 XI11_6/XI0/XI0_3/d__11_ xsel_3_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_10 XI11_6/XI0/XI0_3/d__10_ xsel_3_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_9 XI11_6/XI0/XI0_3/d__9_ xsel_3_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_8 XI11_6/XI0/XI0_3/d__8_ xsel_3_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_7 XI11_6/XI0/XI0_3/d__7_ xsel_3_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_6 XI11_6/XI0/XI0_3/d__6_ xsel_3_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_5 XI11_6/XI0/XI0_3/d__5_ xsel_3_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_4 XI11_6/XI0/XI0_3/d__4_ xsel_3_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_3 XI11_6/XI0/XI0_3/d__3_ xsel_3_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_2 XI11_6/XI0/XI0_3/d__2_ xsel_3_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_1 XI11_6/XI0/XI0_3/d__1_ xsel_3_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_3/MN1_0 XI11_6/XI0/XI0_3/d__0_ xsel_3_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_15 XI11_6/net21_0_ xsel_2_ XI11_6/XI0/XI0_2/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_14 XI11_6/net21_1_ xsel_2_ XI11_6/XI0/XI0_2/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_13 XI11_6/net21_2_ xsel_2_ XI11_6/XI0/XI0_2/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_12 XI11_6/net21_3_ xsel_2_ XI11_6/XI0/XI0_2/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_11 XI11_6/net21_4_ xsel_2_ XI11_6/XI0/XI0_2/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_10 XI11_6/net21_5_ xsel_2_ XI11_6/XI0/XI0_2/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_9 XI11_6/net21_6_ xsel_2_ XI11_6/XI0/XI0_2/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_8 XI11_6/net21_7_ xsel_2_ XI11_6/XI0/XI0_2/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_7 XI11_6/net21_8_ xsel_2_ XI11_6/XI0/XI0_2/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_6 XI11_6/net21_9_ xsel_2_ XI11_6/XI0/XI0_2/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_5 XI11_6/net21_10_ xsel_2_ XI11_6/XI0/XI0_2/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_4 XI11_6/net21_11_ xsel_2_ XI11_6/XI0/XI0_2/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_3 XI11_6/net21_12_ xsel_2_ XI11_6/XI0/XI0_2/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_2 XI11_6/net21_13_ xsel_2_ XI11_6/XI0/XI0_2/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_1 XI11_6/net21_14_ xsel_2_ XI11_6/XI0/XI0_2/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN0_0 XI11_6/net21_15_ xsel_2_ XI11_6/XI0/XI0_2/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_15 XI11_6/XI0/XI0_2/d__15_ xsel_2_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_14 XI11_6/XI0/XI0_2/d__14_ xsel_2_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_13 XI11_6/XI0/XI0_2/d__13_ xsel_2_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_12 XI11_6/XI0/XI0_2/d__12_ xsel_2_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_11 XI11_6/XI0/XI0_2/d__11_ xsel_2_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_10 XI11_6/XI0/XI0_2/d__10_ xsel_2_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_9 XI11_6/XI0/XI0_2/d__9_ xsel_2_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_8 XI11_6/XI0/XI0_2/d__8_ xsel_2_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_7 XI11_6/XI0/XI0_2/d__7_ xsel_2_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_6 XI11_6/XI0/XI0_2/d__6_ xsel_2_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_5 XI11_6/XI0/XI0_2/d__5_ xsel_2_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_4 XI11_6/XI0/XI0_2/d__4_ xsel_2_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_3 XI11_6/XI0/XI0_2/d__3_ xsel_2_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_2 XI11_6/XI0/XI0_2/d__2_ xsel_2_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_1 XI11_6/XI0/XI0_2/d__1_ xsel_2_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_2/MN1_0 XI11_6/XI0/XI0_2/d__0_ xsel_2_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_15 XI11_6/net21_0_ xsel_1_ XI11_6/XI0/XI0_1/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_14 XI11_6/net21_1_ xsel_1_ XI11_6/XI0/XI0_1/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_13 XI11_6/net21_2_ xsel_1_ XI11_6/XI0/XI0_1/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_12 XI11_6/net21_3_ xsel_1_ XI11_6/XI0/XI0_1/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_11 XI11_6/net21_4_ xsel_1_ XI11_6/XI0/XI0_1/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_10 XI11_6/net21_5_ xsel_1_ XI11_6/XI0/XI0_1/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_9 XI11_6/net21_6_ xsel_1_ XI11_6/XI0/XI0_1/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_8 XI11_6/net21_7_ xsel_1_ XI11_6/XI0/XI0_1/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_7 XI11_6/net21_8_ xsel_1_ XI11_6/XI0/XI0_1/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_6 XI11_6/net21_9_ xsel_1_ XI11_6/XI0/XI0_1/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_5 XI11_6/net21_10_ xsel_1_ XI11_6/XI0/XI0_1/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_4 XI11_6/net21_11_ xsel_1_ XI11_6/XI0/XI0_1/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_3 XI11_6/net21_12_ xsel_1_ XI11_6/XI0/XI0_1/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_2 XI11_6/net21_13_ xsel_1_ XI11_6/XI0/XI0_1/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_1 XI11_6/net21_14_ xsel_1_ XI11_6/XI0/XI0_1/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN0_0 XI11_6/net21_15_ xsel_1_ XI11_6/XI0/XI0_1/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_15 XI11_6/XI0/XI0_1/d__15_ xsel_1_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_14 XI11_6/XI0/XI0_1/d__14_ xsel_1_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_13 XI11_6/XI0/XI0_1/d__13_ xsel_1_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_12 XI11_6/XI0/XI0_1/d__12_ xsel_1_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_11 XI11_6/XI0/XI0_1/d__11_ xsel_1_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_10 XI11_6/XI0/XI0_1/d__10_ xsel_1_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_9 XI11_6/XI0/XI0_1/d__9_ xsel_1_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_8 XI11_6/XI0/XI0_1/d__8_ xsel_1_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_7 XI11_6/XI0/XI0_1/d__7_ xsel_1_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_6 XI11_6/XI0/XI0_1/d__6_ xsel_1_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_5 XI11_6/XI0/XI0_1/d__5_ xsel_1_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_4 XI11_6/XI0/XI0_1/d__4_ xsel_1_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_3 XI11_6/XI0/XI0_1/d__3_ xsel_1_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_2 XI11_6/XI0/XI0_1/d__2_ xsel_1_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_1 XI11_6/XI0/XI0_1/d__1_ xsel_1_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_1/MN1_0 XI11_6/XI0/XI0_1/d__0_ xsel_1_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_15 XI11_6/net21_0_ xsel_0_ XI11_6/XI0/XI0_0/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_14 XI11_6/net21_1_ xsel_0_ XI11_6/XI0/XI0_0/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_13 XI11_6/net21_2_ xsel_0_ XI11_6/XI0/XI0_0/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_12 XI11_6/net21_3_ xsel_0_ XI11_6/XI0/XI0_0/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_11 XI11_6/net21_4_ xsel_0_ XI11_6/XI0/XI0_0/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_10 XI11_6/net21_5_ xsel_0_ XI11_6/XI0/XI0_0/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_9 XI11_6/net21_6_ xsel_0_ XI11_6/XI0/XI0_0/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_8 XI11_6/net21_7_ xsel_0_ XI11_6/XI0/XI0_0/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_7 XI11_6/net21_8_ xsel_0_ XI11_6/XI0/XI0_0/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_6 XI11_6/net21_9_ xsel_0_ XI11_6/XI0/XI0_0/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_5 XI11_6/net21_10_ xsel_0_ XI11_6/XI0/XI0_0/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_4 XI11_6/net21_11_ xsel_0_ XI11_6/XI0/XI0_0/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_3 XI11_6/net21_12_ xsel_0_ XI11_6/XI0/XI0_0/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_2 XI11_6/net21_13_ xsel_0_ XI11_6/XI0/XI0_0/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_1 XI11_6/net21_14_ xsel_0_ XI11_6/XI0/XI0_0/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN0_0 XI11_6/net21_15_ xsel_0_ XI11_6/XI0/XI0_0/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_15 XI11_6/XI0/XI0_0/d__15_ xsel_0_ XI11_6/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_14 XI11_6/XI0/XI0_0/d__14_ xsel_0_ XI11_6/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_13 XI11_6/XI0/XI0_0/d__13_ xsel_0_ XI11_6/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_12 XI11_6/XI0/XI0_0/d__12_ xsel_0_ XI11_6/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_11 XI11_6/XI0/XI0_0/d__11_ xsel_0_ XI11_6/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_10 XI11_6/XI0/XI0_0/d__10_ xsel_0_ XI11_6/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_9 XI11_6/XI0/XI0_0/d__9_ xsel_0_ XI11_6/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_8 XI11_6/XI0/XI0_0/d__8_ xsel_0_ XI11_6/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_7 XI11_6/XI0/XI0_0/d__7_ xsel_0_ XI11_6/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_6 XI11_6/XI0/XI0_0/d__6_ xsel_0_ XI11_6/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_5 XI11_6/XI0/XI0_0/d__5_ xsel_0_ XI11_6/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_4 XI11_6/XI0/XI0_0/d__4_ xsel_0_ XI11_6/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_3 XI11_6/XI0/XI0_0/d__3_ xsel_0_ XI11_6/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_2 XI11_6/XI0/XI0_0/d__2_ xsel_0_ XI11_6/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_1 XI11_6/XI0/XI0_0/d__1_ xsel_0_ XI11_6/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_6/XI0/XI0_0/MN1_0 XI11_6/XI0/XI0_0/d__0_ xsel_0_ XI11_6/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI2/MN0_15 XI11_5/net21_0_ ysel_15_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_14 XI11_5/net21_1_ ysel_14_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_13 XI11_5/net21_2_ ysel_13_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_12 XI11_5/net21_3_ ysel_12_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_11 XI11_5/net21_4_ ysel_11_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_10 XI11_5/net21_5_ ysel_10_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_9 XI11_5/net21_6_ ysel_9_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_8 XI11_5/net21_7_ ysel_8_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_7 XI11_5/net21_8_ ysel_7_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_6 XI11_5/net21_9_ ysel_6_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_5 XI11_5/net21_10_ ysel_5_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_4 XI11_5/net21_11_ ysel_4_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_3 XI11_5/net21_12_ ysel_3_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_2 XI11_5/net21_13_ ysel_2_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_1 XI11_5/net21_14_ ysel_1_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN0_0 XI11_5/net21_15_ ysel_0_ XI11_5/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_15 XI11_5/net20_0_ ysel_15_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_14 XI11_5/net20_1_ ysel_14_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_13 XI11_5/net20_2_ ysel_13_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_12 XI11_5/net20_3_ ysel_12_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_11 XI11_5/net20_4_ ysel_11_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_10 XI11_5/net20_5_ ysel_10_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_9 XI11_5/net20_6_ ysel_9_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_8 XI11_5/net20_7_ ysel_8_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_7 XI11_5/net20_8_ ysel_7_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_6 XI11_5/net20_9_ ysel_6_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_5 XI11_5/net20_10_ ysel_5_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_4 XI11_5/net20_11_ ysel_4_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_3 XI11_5/net20_12_ ysel_3_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_2 XI11_5/net20_13_ ysel_2_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_1 XI11_5/net20_14_ ysel_1_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI2/MN1_0 XI11_5/net20_15_ ysel_0_ XI11_5/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_5/XI4/MN8 vdd XI11_5/XI4/net8 XI11_5/net12 vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_5/XI4/MP0 XI11_5/net9 XI11_5/XI4/net23 vdd vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_5/XI4/MP4 XI11_5/net12 XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI4/MP1 XI11_5/net9 XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI4/MP5 XI11_5/net12 XI11_5/preck XI11_5/net9 vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI4/MN7 vdd XI11_5/XI4/net090 DOUT_5_ vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_5/XI4/MP3 gnd XI11_5/XI4/net089 XI11_5/net12 gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_5/XI4/MN5 XI11_5/net9 XI11_5/XI4/net0103 gnd gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_5/XI4/MN4 XI11_5/XI4/data_out_ XI11_5/XI4/net32 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_5/XI4/MN0 XI11_5/XI4/data_out XI11_5/XI4/net52 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_5/XI4/MN9 gnd XI11_5/XI4/net0112 DOUT_5_ gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_5/XI1_15/MP2 XI11_5/net20_0_ XI11_5/preck XI11_5/net21_0_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_15/MP1 XI11_5/net20_0_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_15/MP0 XI11_5/net21_0_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_14/MP2 XI11_5/net20_1_ XI11_5/preck XI11_5/net21_1_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_14/MP1 XI11_5/net20_1_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_14/MP0 XI11_5/net21_1_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_13/MP2 XI11_5/net20_2_ XI11_5/preck XI11_5/net21_2_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_13/MP1 XI11_5/net20_2_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_13/MP0 XI11_5/net21_2_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_12/MP2 XI11_5/net20_3_ XI11_5/preck XI11_5/net21_3_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_12/MP1 XI11_5/net20_3_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_12/MP0 XI11_5/net21_3_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_11/MP2 XI11_5/net20_4_ XI11_5/preck XI11_5/net21_4_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_11/MP1 XI11_5/net20_4_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_11/MP0 XI11_5/net21_4_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_10/MP2 XI11_5/net20_5_ XI11_5/preck XI11_5/net21_5_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_10/MP1 XI11_5/net20_5_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_10/MP0 XI11_5/net21_5_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_9/MP2 XI11_5/net20_6_ XI11_5/preck XI11_5/net21_6_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_9/MP1 XI11_5/net20_6_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_9/MP0 XI11_5/net21_6_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_8/MP2 XI11_5/net20_7_ XI11_5/preck XI11_5/net21_7_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_8/MP1 XI11_5/net20_7_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_8/MP0 XI11_5/net21_7_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_7/MP2 XI11_5/net20_8_ XI11_5/preck XI11_5/net21_8_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_7/MP1 XI11_5/net20_8_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_7/MP0 XI11_5/net21_8_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_6/MP2 XI11_5/net20_9_ XI11_5/preck XI11_5/net21_9_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_6/MP1 XI11_5/net20_9_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_6/MP0 XI11_5/net21_9_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_5/MP2 XI11_5/net20_10_ XI11_5/preck XI11_5/net21_10_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_5/MP1 XI11_5/net20_10_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_5/MP0 XI11_5/net21_10_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_4/MP2 XI11_5/net20_11_ XI11_5/preck XI11_5/net21_11_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_4/MP1 XI11_5/net20_11_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_4/MP0 XI11_5/net21_11_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_3/MP2 XI11_5/net20_12_ XI11_5/preck XI11_5/net21_12_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_3/MP1 XI11_5/net20_12_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_3/MP0 XI11_5/net21_12_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_2/MP2 XI11_5/net20_13_ XI11_5/preck XI11_5/net21_13_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_2/MP1 XI11_5/net20_13_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_2/MP0 XI11_5/net21_13_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_1/MP2 XI11_5/net20_14_ XI11_5/preck XI11_5/net21_14_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_1/MP1 XI11_5/net20_14_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_1/MP0 XI11_5/net21_14_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_0/MP2 XI11_5/net20_15_ XI11_5/preck XI11_5/net21_15_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_5/XI1_0/MP1 XI11_5/net20_15_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI1_0/MP0 XI11_5/net21_15_ XI11_5/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_5/XI0/MN0_15 gnd gnd XI11_5/net21_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_14 gnd gnd XI11_5/net21_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_13 gnd gnd XI11_5/net21_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_12 gnd gnd XI11_5/net21_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_11 gnd gnd XI11_5/net21_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_10 gnd gnd XI11_5/net21_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_9 gnd gnd XI11_5/net21_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_8 gnd gnd XI11_5/net21_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_7 gnd gnd XI11_5/net21_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_6 gnd gnd XI11_5/net21_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_5 gnd gnd XI11_5/net21_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_4 gnd gnd XI11_5/net21_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_3 gnd gnd XI11_5/net21_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_2 gnd gnd XI11_5/net21_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_1 gnd gnd XI11_5/net21_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN0_0 gnd gnd XI11_5/net21_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_15 gnd gnd XI11_5/net20_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_14 gnd gnd XI11_5/net20_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_13 gnd gnd XI11_5/net20_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_12 gnd gnd XI11_5/net20_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_11 gnd gnd XI11_5/net20_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_10 gnd gnd XI11_5/net20_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_9 gnd gnd XI11_5/net20_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_8 gnd gnd XI11_5/net20_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_7 gnd gnd XI11_5/net20_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_6 gnd gnd XI11_5/net20_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_5 gnd gnd XI11_5/net20_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_4 gnd gnd XI11_5/net20_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_3 gnd gnd XI11_5/net20_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_2 gnd gnd XI11_5/net20_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_1 gnd gnd XI11_5/net20_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/MN1_0 gnd gnd XI11_5/net20_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_15 XI11_5/net21_0_ xsel_63_ XI11_5/XI0/XI0_63/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_14 XI11_5/net21_1_ xsel_63_ XI11_5/XI0/XI0_63/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_13 XI11_5/net21_2_ xsel_63_ XI11_5/XI0/XI0_63/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_12 XI11_5/net21_3_ xsel_63_ XI11_5/XI0/XI0_63/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_11 XI11_5/net21_4_ xsel_63_ XI11_5/XI0/XI0_63/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_10 XI11_5/net21_5_ xsel_63_ XI11_5/XI0/XI0_63/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_9 XI11_5/net21_6_ xsel_63_ XI11_5/XI0/XI0_63/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_8 XI11_5/net21_7_ xsel_63_ XI11_5/XI0/XI0_63/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_7 XI11_5/net21_8_ xsel_63_ XI11_5/XI0/XI0_63/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_6 XI11_5/net21_9_ xsel_63_ XI11_5/XI0/XI0_63/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_5 XI11_5/net21_10_ xsel_63_ XI11_5/XI0/XI0_63/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_4 XI11_5/net21_11_ xsel_63_ XI11_5/XI0/XI0_63/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_3 XI11_5/net21_12_ xsel_63_ XI11_5/XI0/XI0_63/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_2 XI11_5/net21_13_ xsel_63_ XI11_5/XI0/XI0_63/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_1 XI11_5/net21_14_ xsel_63_ XI11_5/XI0/XI0_63/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN0_0 XI11_5/net21_15_ xsel_63_ XI11_5/XI0/XI0_63/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_15 XI11_5/XI0/XI0_63/d__15_ xsel_63_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_14 XI11_5/XI0/XI0_63/d__14_ xsel_63_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_13 XI11_5/XI0/XI0_63/d__13_ xsel_63_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_12 XI11_5/XI0/XI0_63/d__12_ xsel_63_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_11 XI11_5/XI0/XI0_63/d__11_ xsel_63_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_10 XI11_5/XI0/XI0_63/d__10_ xsel_63_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_9 XI11_5/XI0/XI0_63/d__9_ xsel_63_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_8 XI11_5/XI0/XI0_63/d__8_ xsel_63_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_7 XI11_5/XI0/XI0_63/d__7_ xsel_63_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_6 XI11_5/XI0/XI0_63/d__6_ xsel_63_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_5 XI11_5/XI0/XI0_63/d__5_ xsel_63_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_4 XI11_5/XI0/XI0_63/d__4_ xsel_63_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_3 XI11_5/XI0/XI0_63/d__3_ xsel_63_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_2 XI11_5/XI0/XI0_63/d__2_ xsel_63_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_1 XI11_5/XI0/XI0_63/d__1_ xsel_63_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_63/MN1_0 XI11_5/XI0/XI0_63/d__0_ xsel_63_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_15 XI11_5/net21_0_ xsel_62_ XI11_5/XI0/XI0_62/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_14 XI11_5/net21_1_ xsel_62_ XI11_5/XI0/XI0_62/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_13 XI11_5/net21_2_ xsel_62_ XI11_5/XI0/XI0_62/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_12 XI11_5/net21_3_ xsel_62_ XI11_5/XI0/XI0_62/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_11 XI11_5/net21_4_ xsel_62_ XI11_5/XI0/XI0_62/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_10 XI11_5/net21_5_ xsel_62_ XI11_5/XI0/XI0_62/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_9 XI11_5/net21_6_ xsel_62_ XI11_5/XI0/XI0_62/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_8 XI11_5/net21_7_ xsel_62_ XI11_5/XI0/XI0_62/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_7 XI11_5/net21_8_ xsel_62_ XI11_5/XI0/XI0_62/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_6 XI11_5/net21_9_ xsel_62_ XI11_5/XI0/XI0_62/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_5 XI11_5/net21_10_ xsel_62_ XI11_5/XI0/XI0_62/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_4 XI11_5/net21_11_ xsel_62_ XI11_5/XI0/XI0_62/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_3 XI11_5/net21_12_ xsel_62_ XI11_5/XI0/XI0_62/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_2 XI11_5/net21_13_ xsel_62_ XI11_5/XI0/XI0_62/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_1 XI11_5/net21_14_ xsel_62_ XI11_5/XI0/XI0_62/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN0_0 XI11_5/net21_15_ xsel_62_ XI11_5/XI0/XI0_62/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_15 XI11_5/XI0/XI0_62/d__15_ xsel_62_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_14 XI11_5/XI0/XI0_62/d__14_ xsel_62_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_13 XI11_5/XI0/XI0_62/d__13_ xsel_62_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_12 XI11_5/XI0/XI0_62/d__12_ xsel_62_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_11 XI11_5/XI0/XI0_62/d__11_ xsel_62_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_10 XI11_5/XI0/XI0_62/d__10_ xsel_62_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_9 XI11_5/XI0/XI0_62/d__9_ xsel_62_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_8 XI11_5/XI0/XI0_62/d__8_ xsel_62_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_7 XI11_5/XI0/XI0_62/d__7_ xsel_62_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_6 XI11_5/XI0/XI0_62/d__6_ xsel_62_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_5 XI11_5/XI0/XI0_62/d__5_ xsel_62_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_4 XI11_5/XI0/XI0_62/d__4_ xsel_62_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_3 XI11_5/XI0/XI0_62/d__3_ xsel_62_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_2 XI11_5/XI0/XI0_62/d__2_ xsel_62_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_1 XI11_5/XI0/XI0_62/d__1_ xsel_62_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_62/MN1_0 XI11_5/XI0/XI0_62/d__0_ xsel_62_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_15 XI11_5/net21_0_ xsel_61_ XI11_5/XI0/XI0_61/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_14 XI11_5/net21_1_ xsel_61_ XI11_5/XI0/XI0_61/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_13 XI11_5/net21_2_ xsel_61_ XI11_5/XI0/XI0_61/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_12 XI11_5/net21_3_ xsel_61_ XI11_5/XI0/XI0_61/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_11 XI11_5/net21_4_ xsel_61_ XI11_5/XI0/XI0_61/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_10 XI11_5/net21_5_ xsel_61_ XI11_5/XI0/XI0_61/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_9 XI11_5/net21_6_ xsel_61_ XI11_5/XI0/XI0_61/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_8 XI11_5/net21_7_ xsel_61_ XI11_5/XI0/XI0_61/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_7 XI11_5/net21_8_ xsel_61_ XI11_5/XI0/XI0_61/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_6 XI11_5/net21_9_ xsel_61_ XI11_5/XI0/XI0_61/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_5 XI11_5/net21_10_ xsel_61_ XI11_5/XI0/XI0_61/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_4 XI11_5/net21_11_ xsel_61_ XI11_5/XI0/XI0_61/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_3 XI11_5/net21_12_ xsel_61_ XI11_5/XI0/XI0_61/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_2 XI11_5/net21_13_ xsel_61_ XI11_5/XI0/XI0_61/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_1 XI11_5/net21_14_ xsel_61_ XI11_5/XI0/XI0_61/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN0_0 XI11_5/net21_15_ xsel_61_ XI11_5/XI0/XI0_61/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_15 XI11_5/XI0/XI0_61/d__15_ xsel_61_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_14 XI11_5/XI0/XI0_61/d__14_ xsel_61_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_13 XI11_5/XI0/XI0_61/d__13_ xsel_61_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_12 XI11_5/XI0/XI0_61/d__12_ xsel_61_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_11 XI11_5/XI0/XI0_61/d__11_ xsel_61_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_10 XI11_5/XI0/XI0_61/d__10_ xsel_61_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_9 XI11_5/XI0/XI0_61/d__9_ xsel_61_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_8 XI11_5/XI0/XI0_61/d__8_ xsel_61_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_7 XI11_5/XI0/XI0_61/d__7_ xsel_61_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_6 XI11_5/XI0/XI0_61/d__6_ xsel_61_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_5 XI11_5/XI0/XI0_61/d__5_ xsel_61_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_4 XI11_5/XI0/XI0_61/d__4_ xsel_61_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_3 XI11_5/XI0/XI0_61/d__3_ xsel_61_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_2 XI11_5/XI0/XI0_61/d__2_ xsel_61_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_1 XI11_5/XI0/XI0_61/d__1_ xsel_61_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_61/MN1_0 XI11_5/XI0/XI0_61/d__0_ xsel_61_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_15 XI11_5/net21_0_ xsel_60_ XI11_5/XI0/XI0_60/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_14 XI11_5/net21_1_ xsel_60_ XI11_5/XI0/XI0_60/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_13 XI11_5/net21_2_ xsel_60_ XI11_5/XI0/XI0_60/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_12 XI11_5/net21_3_ xsel_60_ XI11_5/XI0/XI0_60/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_11 XI11_5/net21_4_ xsel_60_ XI11_5/XI0/XI0_60/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_10 XI11_5/net21_5_ xsel_60_ XI11_5/XI0/XI0_60/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_9 XI11_5/net21_6_ xsel_60_ XI11_5/XI0/XI0_60/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_8 XI11_5/net21_7_ xsel_60_ XI11_5/XI0/XI0_60/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_7 XI11_5/net21_8_ xsel_60_ XI11_5/XI0/XI0_60/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_6 XI11_5/net21_9_ xsel_60_ XI11_5/XI0/XI0_60/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_5 XI11_5/net21_10_ xsel_60_ XI11_5/XI0/XI0_60/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_4 XI11_5/net21_11_ xsel_60_ XI11_5/XI0/XI0_60/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_3 XI11_5/net21_12_ xsel_60_ XI11_5/XI0/XI0_60/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_2 XI11_5/net21_13_ xsel_60_ XI11_5/XI0/XI0_60/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_1 XI11_5/net21_14_ xsel_60_ XI11_5/XI0/XI0_60/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN0_0 XI11_5/net21_15_ xsel_60_ XI11_5/XI0/XI0_60/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_15 XI11_5/XI0/XI0_60/d__15_ xsel_60_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_14 XI11_5/XI0/XI0_60/d__14_ xsel_60_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_13 XI11_5/XI0/XI0_60/d__13_ xsel_60_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_12 XI11_5/XI0/XI0_60/d__12_ xsel_60_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_11 XI11_5/XI0/XI0_60/d__11_ xsel_60_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_10 XI11_5/XI0/XI0_60/d__10_ xsel_60_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_9 XI11_5/XI0/XI0_60/d__9_ xsel_60_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_8 XI11_5/XI0/XI0_60/d__8_ xsel_60_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_7 XI11_5/XI0/XI0_60/d__7_ xsel_60_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_6 XI11_5/XI0/XI0_60/d__6_ xsel_60_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_5 XI11_5/XI0/XI0_60/d__5_ xsel_60_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_4 XI11_5/XI0/XI0_60/d__4_ xsel_60_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_3 XI11_5/XI0/XI0_60/d__3_ xsel_60_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_2 XI11_5/XI0/XI0_60/d__2_ xsel_60_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_1 XI11_5/XI0/XI0_60/d__1_ xsel_60_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_60/MN1_0 XI11_5/XI0/XI0_60/d__0_ xsel_60_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_15 XI11_5/net21_0_ xsel_59_ XI11_5/XI0/XI0_59/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_14 XI11_5/net21_1_ xsel_59_ XI11_5/XI0/XI0_59/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_13 XI11_5/net21_2_ xsel_59_ XI11_5/XI0/XI0_59/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_12 XI11_5/net21_3_ xsel_59_ XI11_5/XI0/XI0_59/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_11 XI11_5/net21_4_ xsel_59_ XI11_5/XI0/XI0_59/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_10 XI11_5/net21_5_ xsel_59_ XI11_5/XI0/XI0_59/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_9 XI11_5/net21_6_ xsel_59_ XI11_5/XI0/XI0_59/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_8 XI11_5/net21_7_ xsel_59_ XI11_5/XI0/XI0_59/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_7 XI11_5/net21_8_ xsel_59_ XI11_5/XI0/XI0_59/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_6 XI11_5/net21_9_ xsel_59_ XI11_5/XI0/XI0_59/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_5 XI11_5/net21_10_ xsel_59_ XI11_5/XI0/XI0_59/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_4 XI11_5/net21_11_ xsel_59_ XI11_5/XI0/XI0_59/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_3 XI11_5/net21_12_ xsel_59_ XI11_5/XI0/XI0_59/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_2 XI11_5/net21_13_ xsel_59_ XI11_5/XI0/XI0_59/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_1 XI11_5/net21_14_ xsel_59_ XI11_5/XI0/XI0_59/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN0_0 XI11_5/net21_15_ xsel_59_ XI11_5/XI0/XI0_59/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_15 XI11_5/XI0/XI0_59/d__15_ xsel_59_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_14 XI11_5/XI0/XI0_59/d__14_ xsel_59_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_13 XI11_5/XI0/XI0_59/d__13_ xsel_59_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_12 XI11_5/XI0/XI0_59/d__12_ xsel_59_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_11 XI11_5/XI0/XI0_59/d__11_ xsel_59_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_10 XI11_5/XI0/XI0_59/d__10_ xsel_59_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_9 XI11_5/XI0/XI0_59/d__9_ xsel_59_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_8 XI11_5/XI0/XI0_59/d__8_ xsel_59_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_7 XI11_5/XI0/XI0_59/d__7_ xsel_59_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_6 XI11_5/XI0/XI0_59/d__6_ xsel_59_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_5 XI11_5/XI0/XI0_59/d__5_ xsel_59_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_4 XI11_5/XI0/XI0_59/d__4_ xsel_59_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_3 XI11_5/XI0/XI0_59/d__3_ xsel_59_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_2 XI11_5/XI0/XI0_59/d__2_ xsel_59_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_1 XI11_5/XI0/XI0_59/d__1_ xsel_59_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_59/MN1_0 XI11_5/XI0/XI0_59/d__0_ xsel_59_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_15 XI11_5/net21_0_ xsel_58_ XI11_5/XI0/XI0_58/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_14 XI11_5/net21_1_ xsel_58_ XI11_5/XI0/XI0_58/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_13 XI11_5/net21_2_ xsel_58_ XI11_5/XI0/XI0_58/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_12 XI11_5/net21_3_ xsel_58_ XI11_5/XI0/XI0_58/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_11 XI11_5/net21_4_ xsel_58_ XI11_5/XI0/XI0_58/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_10 XI11_5/net21_5_ xsel_58_ XI11_5/XI0/XI0_58/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_9 XI11_5/net21_6_ xsel_58_ XI11_5/XI0/XI0_58/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_8 XI11_5/net21_7_ xsel_58_ XI11_5/XI0/XI0_58/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_7 XI11_5/net21_8_ xsel_58_ XI11_5/XI0/XI0_58/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_6 XI11_5/net21_9_ xsel_58_ XI11_5/XI0/XI0_58/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_5 XI11_5/net21_10_ xsel_58_ XI11_5/XI0/XI0_58/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_4 XI11_5/net21_11_ xsel_58_ XI11_5/XI0/XI0_58/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_3 XI11_5/net21_12_ xsel_58_ XI11_5/XI0/XI0_58/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_2 XI11_5/net21_13_ xsel_58_ XI11_5/XI0/XI0_58/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_1 XI11_5/net21_14_ xsel_58_ XI11_5/XI0/XI0_58/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN0_0 XI11_5/net21_15_ xsel_58_ XI11_5/XI0/XI0_58/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_15 XI11_5/XI0/XI0_58/d__15_ xsel_58_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_14 XI11_5/XI0/XI0_58/d__14_ xsel_58_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_13 XI11_5/XI0/XI0_58/d__13_ xsel_58_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_12 XI11_5/XI0/XI0_58/d__12_ xsel_58_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_11 XI11_5/XI0/XI0_58/d__11_ xsel_58_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_10 XI11_5/XI0/XI0_58/d__10_ xsel_58_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_9 XI11_5/XI0/XI0_58/d__9_ xsel_58_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_8 XI11_5/XI0/XI0_58/d__8_ xsel_58_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_7 XI11_5/XI0/XI0_58/d__7_ xsel_58_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_6 XI11_5/XI0/XI0_58/d__6_ xsel_58_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_5 XI11_5/XI0/XI0_58/d__5_ xsel_58_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_4 XI11_5/XI0/XI0_58/d__4_ xsel_58_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_3 XI11_5/XI0/XI0_58/d__3_ xsel_58_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_2 XI11_5/XI0/XI0_58/d__2_ xsel_58_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_1 XI11_5/XI0/XI0_58/d__1_ xsel_58_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_58/MN1_0 XI11_5/XI0/XI0_58/d__0_ xsel_58_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_15 XI11_5/net21_0_ xsel_57_ XI11_5/XI0/XI0_57/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_14 XI11_5/net21_1_ xsel_57_ XI11_5/XI0/XI0_57/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_13 XI11_5/net21_2_ xsel_57_ XI11_5/XI0/XI0_57/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_12 XI11_5/net21_3_ xsel_57_ XI11_5/XI0/XI0_57/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_11 XI11_5/net21_4_ xsel_57_ XI11_5/XI0/XI0_57/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_10 XI11_5/net21_5_ xsel_57_ XI11_5/XI0/XI0_57/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_9 XI11_5/net21_6_ xsel_57_ XI11_5/XI0/XI0_57/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_8 XI11_5/net21_7_ xsel_57_ XI11_5/XI0/XI0_57/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_7 XI11_5/net21_8_ xsel_57_ XI11_5/XI0/XI0_57/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_6 XI11_5/net21_9_ xsel_57_ XI11_5/XI0/XI0_57/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_5 XI11_5/net21_10_ xsel_57_ XI11_5/XI0/XI0_57/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_4 XI11_5/net21_11_ xsel_57_ XI11_5/XI0/XI0_57/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_3 XI11_5/net21_12_ xsel_57_ XI11_5/XI0/XI0_57/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_2 XI11_5/net21_13_ xsel_57_ XI11_5/XI0/XI0_57/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_1 XI11_5/net21_14_ xsel_57_ XI11_5/XI0/XI0_57/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN0_0 XI11_5/net21_15_ xsel_57_ XI11_5/XI0/XI0_57/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_15 XI11_5/XI0/XI0_57/d__15_ xsel_57_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_14 XI11_5/XI0/XI0_57/d__14_ xsel_57_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_13 XI11_5/XI0/XI0_57/d__13_ xsel_57_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_12 XI11_5/XI0/XI0_57/d__12_ xsel_57_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_11 XI11_5/XI0/XI0_57/d__11_ xsel_57_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_10 XI11_5/XI0/XI0_57/d__10_ xsel_57_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_9 XI11_5/XI0/XI0_57/d__9_ xsel_57_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_8 XI11_5/XI0/XI0_57/d__8_ xsel_57_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_7 XI11_5/XI0/XI0_57/d__7_ xsel_57_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_6 XI11_5/XI0/XI0_57/d__6_ xsel_57_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_5 XI11_5/XI0/XI0_57/d__5_ xsel_57_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_4 XI11_5/XI0/XI0_57/d__4_ xsel_57_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_3 XI11_5/XI0/XI0_57/d__3_ xsel_57_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_2 XI11_5/XI0/XI0_57/d__2_ xsel_57_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_1 XI11_5/XI0/XI0_57/d__1_ xsel_57_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_57/MN1_0 XI11_5/XI0/XI0_57/d__0_ xsel_57_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_15 XI11_5/net21_0_ xsel_56_ XI11_5/XI0/XI0_56/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_14 XI11_5/net21_1_ xsel_56_ XI11_5/XI0/XI0_56/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_13 XI11_5/net21_2_ xsel_56_ XI11_5/XI0/XI0_56/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_12 XI11_5/net21_3_ xsel_56_ XI11_5/XI0/XI0_56/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_11 XI11_5/net21_4_ xsel_56_ XI11_5/XI0/XI0_56/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_10 XI11_5/net21_5_ xsel_56_ XI11_5/XI0/XI0_56/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_9 XI11_5/net21_6_ xsel_56_ XI11_5/XI0/XI0_56/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_8 XI11_5/net21_7_ xsel_56_ XI11_5/XI0/XI0_56/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_7 XI11_5/net21_8_ xsel_56_ XI11_5/XI0/XI0_56/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_6 XI11_5/net21_9_ xsel_56_ XI11_5/XI0/XI0_56/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_5 XI11_5/net21_10_ xsel_56_ XI11_5/XI0/XI0_56/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_4 XI11_5/net21_11_ xsel_56_ XI11_5/XI0/XI0_56/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_3 XI11_5/net21_12_ xsel_56_ XI11_5/XI0/XI0_56/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_2 XI11_5/net21_13_ xsel_56_ XI11_5/XI0/XI0_56/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_1 XI11_5/net21_14_ xsel_56_ XI11_5/XI0/XI0_56/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN0_0 XI11_5/net21_15_ xsel_56_ XI11_5/XI0/XI0_56/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_15 XI11_5/XI0/XI0_56/d__15_ xsel_56_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_14 XI11_5/XI0/XI0_56/d__14_ xsel_56_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_13 XI11_5/XI0/XI0_56/d__13_ xsel_56_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_12 XI11_5/XI0/XI0_56/d__12_ xsel_56_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_11 XI11_5/XI0/XI0_56/d__11_ xsel_56_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_10 XI11_5/XI0/XI0_56/d__10_ xsel_56_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_9 XI11_5/XI0/XI0_56/d__9_ xsel_56_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_8 XI11_5/XI0/XI0_56/d__8_ xsel_56_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_7 XI11_5/XI0/XI0_56/d__7_ xsel_56_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_6 XI11_5/XI0/XI0_56/d__6_ xsel_56_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_5 XI11_5/XI0/XI0_56/d__5_ xsel_56_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_4 XI11_5/XI0/XI0_56/d__4_ xsel_56_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_3 XI11_5/XI0/XI0_56/d__3_ xsel_56_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_2 XI11_5/XI0/XI0_56/d__2_ xsel_56_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_1 XI11_5/XI0/XI0_56/d__1_ xsel_56_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_56/MN1_0 XI11_5/XI0/XI0_56/d__0_ xsel_56_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_15 XI11_5/net21_0_ xsel_55_ XI11_5/XI0/XI0_55/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_14 XI11_5/net21_1_ xsel_55_ XI11_5/XI0/XI0_55/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_13 XI11_5/net21_2_ xsel_55_ XI11_5/XI0/XI0_55/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_12 XI11_5/net21_3_ xsel_55_ XI11_5/XI0/XI0_55/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_11 XI11_5/net21_4_ xsel_55_ XI11_5/XI0/XI0_55/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_10 XI11_5/net21_5_ xsel_55_ XI11_5/XI0/XI0_55/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_9 XI11_5/net21_6_ xsel_55_ XI11_5/XI0/XI0_55/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_8 XI11_5/net21_7_ xsel_55_ XI11_5/XI0/XI0_55/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_7 XI11_5/net21_8_ xsel_55_ XI11_5/XI0/XI0_55/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_6 XI11_5/net21_9_ xsel_55_ XI11_5/XI0/XI0_55/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_5 XI11_5/net21_10_ xsel_55_ XI11_5/XI0/XI0_55/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_4 XI11_5/net21_11_ xsel_55_ XI11_5/XI0/XI0_55/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_3 XI11_5/net21_12_ xsel_55_ XI11_5/XI0/XI0_55/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_2 XI11_5/net21_13_ xsel_55_ XI11_5/XI0/XI0_55/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_1 XI11_5/net21_14_ xsel_55_ XI11_5/XI0/XI0_55/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN0_0 XI11_5/net21_15_ xsel_55_ XI11_5/XI0/XI0_55/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_15 XI11_5/XI0/XI0_55/d__15_ xsel_55_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_14 XI11_5/XI0/XI0_55/d__14_ xsel_55_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_13 XI11_5/XI0/XI0_55/d__13_ xsel_55_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_12 XI11_5/XI0/XI0_55/d__12_ xsel_55_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_11 XI11_5/XI0/XI0_55/d__11_ xsel_55_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_10 XI11_5/XI0/XI0_55/d__10_ xsel_55_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_9 XI11_5/XI0/XI0_55/d__9_ xsel_55_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_8 XI11_5/XI0/XI0_55/d__8_ xsel_55_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_7 XI11_5/XI0/XI0_55/d__7_ xsel_55_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_6 XI11_5/XI0/XI0_55/d__6_ xsel_55_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_5 XI11_5/XI0/XI0_55/d__5_ xsel_55_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_4 XI11_5/XI0/XI0_55/d__4_ xsel_55_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_3 XI11_5/XI0/XI0_55/d__3_ xsel_55_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_2 XI11_5/XI0/XI0_55/d__2_ xsel_55_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_1 XI11_5/XI0/XI0_55/d__1_ xsel_55_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_55/MN1_0 XI11_5/XI0/XI0_55/d__0_ xsel_55_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_15 XI11_5/net21_0_ xsel_54_ XI11_5/XI0/XI0_54/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_14 XI11_5/net21_1_ xsel_54_ XI11_5/XI0/XI0_54/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_13 XI11_5/net21_2_ xsel_54_ XI11_5/XI0/XI0_54/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_12 XI11_5/net21_3_ xsel_54_ XI11_5/XI0/XI0_54/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_11 XI11_5/net21_4_ xsel_54_ XI11_5/XI0/XI0_54/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_10 XI11_5/net21_5_ xsel_54_ XI11_5/XI0/XI0_54/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_9 XI11_5/net21_6_ xsel_54_ XI11_5/XI0/XI0_54/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_8 XI11_5/net21_7_ xsel_54_ XI11_5/XI0/XI0_54/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_7 XI11_5/net21_8_ xsel_54_ XI11_5/XI0/XI0_54/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_6 XI11_5/net21_9_ xsel_54_ XI11_5/XI0/XI0_54/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_5 XI11_5/net21_10_ xsel_54_ XI11_5/XI0/XI0_54/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_4 XI11_5/net21_11_ xsel_54_ XI11_5/XI0/XI0_54/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_3 XI11_5/net21_12_ xsel_54_ XI11_5/XI0/XI0_54/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_2 XI11_5/net21_13_ xsel_54_ XI11_5/XI0/XI0_54/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_1 XI11_5/net21_14_ xsel_54_ XI11_5/XI0/XI0_54/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN0_0 XI11_5/net21_15_ xsel_54_ XI11_5/XI0/XI0_54/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_15 XI11_5/XI0/XI0_54/d__15_ xsel_54_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_14 XI11_5/XI0/XI0_54/d__14_ xsel_54_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_13 XI11_5/XI0/XI0_54/d__13_ xsel_54_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_12 XI11_5/XI0/XI0_54/d__12_ xsel_54_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_11 XI11_5/XI0/XI0_54/d__11_ xsel_54_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_10 XI11_5/XI0/XI0_54/d__10_ xsel_54_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_9 XI11_5/XI0/XI0_54/d__9_ xsel_54_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_8 XI11_5/XI0/XI0_54/d__8_ xsel_54_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_7 XI11_5/XI0/XI0_54/d__7_ xsel_54_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_6 XI11_5/XI0/XI0_54/d__6_ xsel_54_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_5 XI11_5/XI0/XI0_54/d__5_ xsel_54_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_4 XI11_5/XI0/XI0_54/d__4_ xsel_54_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_3 XI11_5/XI0/XI0_54/d__3_ xsel_54_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_2 XI11_5/XI0/XI0_54/d__2_ xsel_54_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_1 XI11_5/XI0/XI0_54/d__1_ xsel_54_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_54/MN1_0 XI11_5/XI0/XI0_54/d__0_ xsel_54_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_15 XI11_5/net21_0_ xsel_53_ XI11_5/XI0/XI0_53/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_14 XI11_5/net21_1_ xsel_53_ XI11_5/XI0/XI0_53/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_13 XI11_5/net21_2_ xsel_53_ XI11_5/XI0/XI0_53/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_12 XI11_5/net21_3_ xsel_53_ XI11_5/XI0/XI0_53/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_11 XI11_5/net21_4_ xsel_53_ XI11_5/XI0/XI0_53/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_10 XI11_5/net21_5_ xsel_53_ XI11_5/XI0/XI0_53/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_9 XI11_5/net21_6_ xsel_53_ XI11_5/XI0/XI0_53/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_8 XI11_5/net21_7_ xsel_53_ XI11_5/XI0/XI0_53/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_7 XI11_5/net21_8_ xsel_53_ XI11_5/XI0/XI0_53/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_6 XI11_5/net21_9_ xsel_53_ XI11_5/XI0/XI0_53/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_5 XI11_5/net21_10_ xsel_53_ XI11_5/XI0/XI0_53/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_4 XI11_5/net21_11_ xsel_53_ XI11_5/XI0/XI0_53/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_3 XI11_5/net21_12_ xsel_53_ XI11_5/XI0/XI0_53/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_2 XI11_5/net21_13_ xsel_53_ XI11_5/XI0/XI0_53/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_1 XI11_5/net21_14_ xsel_53_ XI11_5/XI0/XI0_53/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN0_0 XI11_5/net21_15_ xsel_53_ XI11_5/XI0/XI0_53/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_15 XI11_5/XI0/XI0_53/d__15_ xsel_53_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_14 XI11_5/XI0/XI0_53/d__14_ xsel_53_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_13 XI11_5/XI0/XI0_53/d__13_ xsel_53_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_12 XI11_5/XI0/XI0_53/d__12_ xsel_53_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_11 XI11_5/XI0/XI0_53/d__11_ xsel_53_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_10 XI11_5/XI0/XI0_53/d__10_ xsel_53_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_9 XI11_5/XI0/XI0_53/d__9_ xsel_53_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_8 XI11_5/XI0/XI0_53/d__8_ xsel_53_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_7 XI11_5/XI0/XI0_53/d__7_ xsel_53_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_6 XI11_5/XI0/XI0_53/d__6_ xsel_53_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_5 XI11_5/XI0/XI0_53/d__5_ xsel_53_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_4 XI11_5/XI0/XI0_53/d__4_ xsel_53_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_3 XI11_5/XI0/XI0_53/d__3_ xsel_53_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_2 XI11_5/XI0/XI0_53/d__2_ xsel_53_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_1 XI11_5/XI0/XI0_53/d__1_ xsel_53_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_53/MN1_0 XI11_5/XI0/XI0_53/d__0_ xsel_53_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_15 XI11_5/net21_0_ xsel_52_ XI11_5/XI0/XI0_52/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_14 XI11_5/net21_1_ xsel_52_ XI11_5/XI0/XI0_52/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_13 XI11_5/net21_2_ xsel_52_ XI11_5/XI0/XI0_52/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_12 XI11_5/net21_3_ xsel_52_ XI11_5/XI0/XI0_52/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_11 XI11_5/net21_4_ xsel_52_ XI11_5/XI0/XI0_52/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_10 XI11_5/net21_5_ xsel_52_ XI11_5/XI0/XI0_52/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_9 XI11_5/net21_6_ xsel_52_ XI11_5/XI0/XI0_52/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_8 XI11_5/net21_7_ xsel_52_ XI11_5/XI0/XI0_52/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_7 XI11_5/net21_8_ xsel_52_ XI11_5/XI0/XI0_52/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_6 XI11_5/net21_9_ xsel_52_ XI11_5/XI0/XI0_52/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_5 XI11_5/net21_10_ xsel_52_ XI11_5/XI0/XI0_52/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_4 XI11_5/net21_11_ xsel_52_ XI11_5/XI0/XI0_52/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_3 XI11_5/net21_12_ xsel_52_ XI11_5/XI0/XI0_52/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_2 XI11_5/net21_13_ xsel_52_ XI11_5/XI0/XI0_52/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_1 XI11_5/net21_14_ xsel_52_ XI11_5/XI0/XI0_52/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN0_0 XI11_5/net21_15_ xsel_52_ XI11_5/XI0/XI0_52/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_15 XI11_5/XI0/XI0_52/d__15_ xsel_52_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_14 XI11_5/XI0/XI0_52/d__14_ xsel_52_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_13 XI11_5/XI0/XI0_52/d__13_ xsel_52_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_12 XI11_5/XI0/XI0_52/d__12_ xsel_52_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_11 XI11_5/XI0/XI0_52/d__11_ xsel_52_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_10 XI11_5/XI0/XI0_52/d__10_ xsel_52_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_9 XI11_5/XI0/XI0_52/d__9_ xsel_52_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_8 XI11_5/XI0/XI0_52/d__8_ xsel_52_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_7 XI11_5/XI0/XI0_52/d__7_ xsel_52_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_6 XI11_5/XI0/XI0_52/d__6_ xsel_52_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_5 XI11_5/XI0/XI0_52/d__5_ xsel_52_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_4 XI11_5/XI0/XI0_52/d__4_ xsel_52_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_3 XI11_5/XI0/XI0_52/d__3_ xsel_52_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_2 XI11_5/XI0/XI0_52/d__2_ xsel_52_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_1 XI11_5/XI0/XI0_52/d__1_ xsel_52_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_52/MN1_0 XI11_5/XI0/XI0_52/d__0_ xsel_52_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_15 XI11_5/net21_0_ xsel_51_ XI11_5/XI0/XI0_51/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_14 XI11_5/net21_1_ xsel_51_ XI11_5/XI0/XI0_51/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_13 XI11_5/net21_2_ xsel_51_ XI11_5/XI0/XI0_51/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_12 XI11_5/net21_3_ xsel_51_ XI11_5/XI0/XI0_51/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_11 XI11_5/net21_4_ xsel_51_ XI11_5/XI0/XI0_51/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_10 XI11_5/net21_5_ xsel_51_ XI11_5/XI0/XI0_51/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_9 XI11_5/net21_6_ xsel_51_ XI11_5/XI0/XI0_51/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_8 XI11_5/net21_7_ xsel_51_ XI11_5/XI0/XI0_51/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_7 XI11_5/net21_8_ xsel_51_ XI11_5/XI0/XI0_51/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_6 XI11_5/net21_9_ xsel_51_ XI11_5/XI0/XI0_51/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_5 XI11_5/net21_10_ xsel_51_ XI11_5/XI0/XI0_51/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_4 XI11_5/net21_11_ xsel_51_ XI11_5/XI0/XI0_51/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_3 XI11_5/net21_12_ xsel_51_ XI11_5/XI0/XI0_51/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_2 XI11_5/net21_13_ xsel_51_ XI11_5/XI0/XI0_51/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_1 XI11_5/net21_14_ xsel_51_ XI11_5/XI0/XI0_51/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN0_0 XI11_5/net21_15_ xsel_51_ XI11_5/XI0/XI0_51/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_15 XI11_5/XI0/XI0_51/d__15_ xsel_51_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_14 XI11_5/XI0/XI0_51/d__14_ xsel_51_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_13 XI11_5/XI0/XI0_51/d__13_ xsel_51_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_12 XI11_5/XI0/XI0_51/d__12_ xsel_51_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_11 XI11_5/XI0/XI0_51/d__11_ xsel_51_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_10 XI11_5/XI0/XI0_51/d__10_ xsel_51_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_9 XI11_5/XI0/XI0_51/d__9_ xsel_51_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_8 XI11_5/XI0/XI0_51/d__8_ xsel_51_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_7 XI11_5/XI0/XI0_51/d__7_ xsel_51_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_6 XI11_5/XI0/XI0_51/d__6_ xsel_51_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_5 XI11_5/XI0/XI0_51/d__5_ xsel_51_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_4 XI11_5/XI0/XI0_51/d__4_ xsel_51_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_3 XI11_5/XI0/XI0_51/d__3_ xsel_51_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_2 XI11_5/XI0/XI0_51/d__2_ xsel_51_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_1 XI11_5/XI0/XI0_51/d__1_ xsel_51_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_51/MN1_0 XI11_5/XI0/XI0_51/d__0_ xsel_51_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_15 XI11_5/net21_0_ xsel_50_ XI11_5/XI0/XI0_50/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_14 XI11_5/net21_1_ xsel_50_ XI11_5/XI0/XI0_50/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_13 XI11_5/net21_2_ xsel_50_ XI11_5/XI0/XI0_50/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_12 XI11_5/net21_3_ xsel_50_ XI11_5/XI0/XI0_50/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_11 XI11_5/net21_4_ xsel_50_ XI11_5/XI0/XI0_50/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_10 XI11_5/net21_5_ xsel_50_ XI11_5/XI0/XI0_50/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_9 XI11_5/net21_6_ xsel_50_ XI11_5/XI0/XI0_50/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_8 XI11_5/net21_7_ xsel_50_ XI11_5/XI0/XI0_50/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_7 XI11_5/net21_8_ xsel_50_ XI11_5/XI0/XI0_50/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_6 XI11_5/net21_9_ xsel_50_ XI11_5/XI0/XI0_50/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_5 XI11_5/net21_10_ xsel_50_ XI11_5/XI0/XI0_50/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_4 XI11_5/net21_11_ xsel_50_ XI11_5/XI0/XI0_50/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_3 XI11_5/net21_12_ xsel_50_ XI11_5/XI0/XI0_50/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_2 XI11_5/net21_13_ xsel_50_ XI11_5/XI0/XI0_50/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_1 XI11_5/net21_14_ xsel_50_ XI11_5/XI0/XI0_50/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN0_0 XI11_5/net21_15_ xsel_50_ XI11_5/XI0/XI0_50/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_15 XI11_5/XI0/XI0_50/d__15_ xsel_50_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_14 XI11_5/XI0/XI0_50/d__14_ xsel_50_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_13 XI11_5/XI0/XI0_50/d__13_ xsel_50_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_12 XI11_5/XI0/XI0_50/d__12_ xsel_50_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_11 XI11_5/XI0/XI0_50/d__11_ xsel_50_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_10 XI11_5/XI0/XI0_50/d__10_ xsel_50_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_9 XI11_5/XI0/XI0_50/d__9_ xsel_50_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_8 XI11_5/XI0/XI0_50/d__8_ xsel_50_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_7 XI11_5/XI0/XI0_50/d__7_ xsel_50_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_6 XI11_5/XI0/XI0_50/d__6_ xsel_50_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_5 XI11_5/XI0/XI0_50/d__5_ xsel_50_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_4 XI11_5/XI0/XI0_50/d__4_ xsel_50_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_3 XI11_5/XI0/XI0_50/d__3_ xsel_50_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_2 XI11_5/XI0/XI0_50/d__2_ xsel_50_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_1 XI11_5/XI0/XI0_50/d__1_ xsel_50_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_50/MN1_0 XI11_5/XI0/XI0_50/d__0_ xsel_50_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_15 XI11_5/net21_0_ xsel_49_ XI11_5/XI0/XI0_49/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_14 XI11_5/net21_1_ xsel_49_ XI11_5/XI0/XI0_49/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_13 XI11_5/net21_2_ xsel_49_ XI11_5/XI0/XI0_49/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_12 XI11_5/net21_3_ xsel_49_ XI11_5/XI0/XI0_49/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_11 XI11_5/net21_4_ xsel_49_ XI11_5/XI0/XI0_49/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_10 XI11_5/net21_5_ xsel_49_ XI11_5/XI0/XI0_49/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_9 XI11_5/net21_6_ xsel_49_ XI11_5/XI0/XI0_49/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_8 XI11_5/net21_7_ xsel_49_ XI11_5/XI0/XI0_49/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_7 XI11_5/net21_8_ xsel_49_ XI11_5/XI0/XI0_49/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_6 XI11_5/net21_9_ xsel_49_ XI11_5/XI0/XI0_49/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_5 XI11_5/net21_10_ xsel_49_ XI11_5/XI0/XI0_49/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_4 XI11_5/net21_11_ xsel_49_ XI11_5/XI0/XI0_49/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_3 XI11_5/net21_12_ xsel_49_ XI11_5/XI0/XI0_49/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_2 XI11_5/net21_13_ xsel_49_ XI11_5/XI0/XI0_49/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_1 XI11_5/net21_14_ xsel_49_ XI11_5/XI0/XI0_49/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN0_0 XI11_5/net21_15_ xsel_49_ XI11_5/XI0/XI0_49/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_15 XI11_5/XI0/XI0_49/d__15_ xsel_49_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_14 XI11_5/XI0/XI0_49/d__14_ xsel_49_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_13 XI11_5/XI0/XI0_49/d__13_ xsel_49_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_12 XI11_5/XI0/XI0_49/d__12_ xsel_49_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_11 XI11_5/XI0/XI0_49/d__11_ xsel_49_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_10 XI11_5/XI0/XI0_49/d__10_ xsel_49_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_9 XI11_5/XI0/XI0_49/d__9_ xsel_49_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_8 XI11_5/XI0/XI0_49/d__8_ xsel_49_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_7 XI11_5/XI0/XI0_49/d__7_ xsel_49_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_6 XI11_5/XI0/XI0_49/d__6_ xsel_49_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_5 XI11_5/XI0/XI0_49/d__5_ xsel_49_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_4 XI11_5/XI0/XI0_49/d__4_ xsel_49_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_3 XI11_5/XI0/XI0_49/d__3_ xsel_49_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_2 XI11_5/XI0/XI0_49/d__2_ xsel_49_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_1 XI11_5/XI0/XI0_49/d__1_ xsel_49_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_49/MN1_0 XI11_5/XI0/XI0_49/d__0_ xsel_49_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_15 XI11_5/net21_0_ xsel_48_ XI11_5/XI0/XI0_48/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_14 XI11_5/net21_1_ xsel_48_ XI11_5/XI0/XI0_48/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_13 XI11_5/net21_2_ xsel_48_ XI11_5/XI0/XI0_48/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_12 XI11_5/net21_3_ xsel_48_ XI11_5/XI0/XI0_48/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_11 XI11_5/net21_4_ xsel_48_ XI11_5/XI0/XI0_48/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_10 XI11_5/net21_5_ xsel_48_ XI11_5/XI0/XI0_48/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_9 XI11_5/net21_6_ xsel_48_ XI11_5/XI0/XI0_48/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_8 XI11_5/net21_7_ xsel_48_ XI11_5/XI0/XI0_48/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_7 XI11_5/net21_8_ xsel_48_ XI11_5/XI0/XI0_48/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_6 XI11_5/net21_9_ xsel_48_ XI11_5/XI0/XI0_48/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_5 XI11_5/net21_10_ xsel_48_ XI11_5/XI0/XI0_48/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_4 XI11_5/net21_11_ xsel_48_ XI11_5/XI0/XI0_48/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_3 XI11_5/net21_12_ xsel_48_ XI11_5/XI0/XI0_48/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_2 XI11_5/net21_13_ xsel_48_ XI11_5/XI0/XI0_48/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_1 XI11_5/net21_14_ xsel_48_ XI11_5/XI0/XI0_48/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN0_0 XI11_5/net21_15_ xsel_48_ XI11_5/XI0/XI0_48/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_15 XI11_5/XI0/XI0_48/d__15_ xsel_48_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_14 XI11_5/XI0/XI0_48/d__14_ xsel_48_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_13 XI11_5/XI0/XI0_48/d__13_ xsel_48_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_12 XI11_5/XI0/XI0_48/d__12_ xsel_48_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_11 XI11_5/XI0/XI0_48/d__11_ xsel_48_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_10 XI11_5/XI0/XI0_48/d__10_ xsel_48_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_9 XI11_5/XI0/XI0_48/d__9_ xsel_48_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_8 XI11_5/XI0/XI0_48/d__8_ xsel_48_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_7 XI11_5/XI0/XI0_48/d__7_ xsel_48_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_6 XI11_5/XI0/XI0_48/d__6_ xsel_48_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_5 XI11_5/XI0/XI0_48/d__5_ xsel_48_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_4 XI11_5/XI0/XI0_48/d__4_ xsel_48_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_3 XI11_5/XI0/XI0_48/d__3_ xsel_48_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_2 XI11_5/XI0/XI0_48/d__2_ xsel_48_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_1 XI11_5/XI0/XI0_48/d__1_ xsel_48_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_48/MN1_0 XI11_5/XI0/XI0_48/d__0_ xsel_48_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_15 XI11_5/net21_0_ xsel_47_ XI11_5/XI0/XI0_47/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_14 XI11_5/net21_1_ xsel_47_ XI11_5/XI0/XI0_47/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_13 XI11_5/net21_2_ xsel_47_ XI11_5/XI0/XI0_47/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_12 XI11_5/net21_3_ xsel_47_ XI11_5/XI0/XI0_47/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_11 XI11_5/net21_4_ xsel_47_ XI11_5/XI0/XI0_47/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_10 XI11_5/net21_5_ xsel_47_ XI11_5/XI0/XI0_47/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_9 XI11_5/net21_6_ xsel_47_ XI11_5/XI0/XI0_47/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_8 XI11_5/net21_7_ xsel_47_ XI11_5/XI0/XI0_47/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_7 XI11_5/net21_8_ xsel_47_ XI11_5/XI0/XI0_47/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_6 XI11_5/net21_9_ xsel_47_ XI11_5/XI0/XI0_47/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_5 XI11_5/net21_10_ xsel_47_ XI11_5/XI0/XI0_47/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_4 XI11_5/net21_11_ xsel_47_ XI11_5/XI0/XI0_47/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_3 XI11_5/net21_12_ xsel_47_ XI11_5/XI0/XI0_47/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_2 XI11_5/net21_13_ xsel_47_ XI11_5/XI0/XI0_47/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_1 XI11_5/net21_14_ xsel_47_ XI11_5/XI0/XI0_47/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN0_0 XI11_5/net21_15_ xsel_47_ XI11_5/XI0/XI0_47/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_15 XI11_5/XI0/XI0_47/d__15_ xsel_47_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_14 XI11_5/XI0/XI0_47/d__14_ xsel_47_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_13 XI11_5/XI0/XI0_47/d__13_ xsel_47_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_12 XI11_5/XI0/XI0_47/d__12_ xsel_47_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_11 XI11_5/XI0/XI0_47/d__11_ xsel_47_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_10 XI11_5/XI0/XI0_47/d__10_ xsel_47_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_9 XI11_5/XI0/XI0_47/d__9_ xsel_47_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_8 XI11_5/XI0/XI0_47/d__8_ xsel_47_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_7 XI11_5/XI0/XI0_47/d__7_ xsel_47_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_6 XI11_5/XI0/XI0_47/d__6_ xsel_47_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_5 XI11_5/XI0/XI0_47/d__5_ xsel_47_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_4 XI11_5/XI0/XI0_47/d__4_ xsel_47_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_3 XI11_5/XI0/XI0_47/d__3_ xsel_47_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_2 XI11_5/XI0/XI0_47/d__2_ xsel_47_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_1 XI11_5/XI0/XI0_47/d__1_ xsel_47_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_47/MN1_0 XI11_5/XI0/XI0_47/d__0_ xsel_47_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_15 XI11_5/net21_0_ xsel_46_ XI11_5/XI0/XI0_46/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_14 XI11_5/net21_1_ xsel_46_ XI11_5/XI0/XI0_46/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_13 XI11_5/net21_2_ xsel_46_ XI11_5/XI0/XI0_46/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_12 XI11_5/net21_3_ xsel_46_ XI11_5/XI0/XI0_46/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_11 XI11_5/net21_4_ xsel_46_ XI11_5/XI0/XI0_46/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_10 XI11_5/net21_5_ xsel_46_ XI11_5/XI0/XI0_46/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_9 XI11_5/net21_6_ xsel_46_ XI11_5/XI0/XI0_46/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_8 XI11_5/net21_7_ xsel_46_ XI11_5/XI0/XI0_46/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_7 XI11_5/net21_8_ xsel_46_ XI11_5/XI0/XI0_46/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_6 XI11_5/net21_9_ xsel_46_ XI11_5/XI0/XI0_46/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_5 XI11_5/net21_10_ xsel_46_ XI11_5/XI0/XI0_46/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_4 XI11_5/net21_11_ xsel_46_ XI11_5/XI0/XI0_46/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_3 XI11_5/net21_12_ xsel_46_ XI11_5/XI0/XI0_46/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_2 XI11_5/net21_13_ xsel_46_ XI11_5/XI0/XI0_46/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_1 XI11_5/net21_14_ xsel_46_ XI11_5/XI0/XI0_46/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN0_0 XI11_5/net21_15_ xsel_46_ XI11_5/XI0/XI0_46/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_15 XI11_5/XI0/XI0_46/d__15_ xsel_46_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_14 XI11_5/XI0/XI0_46/d__14_ xsel_46_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_13 XI11_5/XI0/XI0_46/d__13_ xsel_46_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_12 XI11_5/XI0/XI0_46/d__12_ xsel_46_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_11 XI11_5/XI0/XI0_46/d__11_ xsel_46_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_10 XI11_5/XI0/XI0_46/d__10_ xsel_46_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_9 XI11_5/XI0/XI0_46/d__9_ xsel_46_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_8 XI11_5/XI0/XI0_46/d__8_ xsel_46_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_7 XI11_5/XI0/XI0_46/d__7_ xsel_46_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_6 XI11_5/XI0/XI0_46/d__6_ xsel_46_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_5 XI11_5/XI0/XI0_46/d__5_ xsel_46_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_4 XI11_5/XI0/XI0_46/d__4_ xsel_46_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_3 XI11_5/XI0/XI0_46/d__3_ xsel_46_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_2 XI11_5/XI0/XI0_46/d__2_ xsel_46_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_1 XI11_5/XI0/XI0_46/d__1_ xsel_46_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_46/MN1_0 XI11_5/XI0/XI0_46/d__0_ xsel_46_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_15 XI11_5/net21_0_ xsel_45_ XI11_5/XI0/XI0_45/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_14 XI11_5/net21_1_ xsel_45_ XI11_5/XI0/XI0_45/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_13 XI11_5/net21_2_ xsel_45_ XI11_5/XI0/XI0_45/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_12 XI11_5/net21_3_ xsel_45_ XI11_5/XI0/XI0_45/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_11 XI11_5/net21_4_ xsel_45_ XI11_5/XI0/XI0_45/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_10 XI11_5/net21_5_ xsel_45_ XI11_5/XI0/XI0_45/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_9 XI11_5/net21_6_ xsel_45_ XI11_5/XI0/XI0_45/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_8 XI11_5/net21_7_ xsel_45_ XI11_5/XI0/XI0_45/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_7 XI11_5/net21_8_ xsel_45_ XI11_5/XI0/XI0_45/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_6 XI11_5/net21_9_ xsel_45_ XI11_5/XI0/XI0_45/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_5 XI11_5/net21_10_ xsel_45_ XI11_5/XI0/XI0_45/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_4 XI11_5/net21_11_ xsel_45_ XI11_5/XI0/XI0_45/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_3 XI11_5/net21_12_ xsel_45_ XI11_5/XI0/XI0_45/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_2 XI11_5/net21_13_ xsel_45_ XI11_5/XI0/XI0_45/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_1 XI11_5/net21_14_ xsel_45_ XI11_5/XI0/XI0_45/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN0_0 XI11_5/net21_15_ xsel_45_ XI11_5/XI0/XI0_45/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_15 XI11_5/XI0/XI0_45/d__15_ xsel_45_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_14 XI11_5/XI0/XI0_45/d__14_ xsel_45_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_13 XI11_5/XI0/XI0_45/d__13_ xsel_45_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_12 XI11_5/XI0/XI0_45/d__12_ xsel_45_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_11 XI11_5/XI0/XI0_45/d__11_ xsel_45_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_10 XI11_5/XI0/XI0_45/d__10_ xsel_45_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_9 XI11_5/XI0/XI0_45/d__9_ xsel_45_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_8 XI11_5/XI0/XI0_45/d__8_ xsel_45_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_7 XI11_5/XI0/XI0_45/d__7_ xsel_45_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_6 XI11_5/XI0/XI0_45/d__6_ xsel_45_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_5 XI11_5/XI0/XI0_45/d__5_ xsel_45_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_4 XI11_5/XI0/XI0_45/d__4_ xsel_45_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_3 XI11_5/XI0/XI0_45/d__3_ xsel_45_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_2 XI11_5/XI0/XI0_45/d__2_ xsel_45_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_1 XI11_5/XI0/XI0_45/d__1_ xsel_45_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_45/MN1_0 XI11_5/XI0/XI0_45/d__0_ xsel_45_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_15 XI11_5/net21_0_ xsel_44_ XI11_5/XI0/XI0_44/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_14 XI11_5/net21_1_ xsel_44_ XI11_5/XI0/XI0_44/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_13 XI11_5/net21_2_ xsel_44_ XI11_5/XI0/XI0_44/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_12 XI11_5/net21_3_ xsel_44_ XI11_5/XI0/XI0_44/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_11 XI11_5/net21_4_ xsel_44_ XI11_5/XI0/XI0_44/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_10 XI11_5/net21_5_ xsel_44_ XI11_5/XI0/XI0_44/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_9 XI11_5/net21_6_ xsel_44_ XI11_5/XI0/XI0_44/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_8 XI11_5/net21_7_ xsel_44_ XI11_5/XI0/XI0_44/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_7 XI11_5/net21_8_ xsel_44_ XI11_5/XI0/XI0_44/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_6 XI11_5/net21_9_ xsel_44_ XI11_5/XI0/XI0_44/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_5 XI11_5/net21_10_ xsel_44_ XI11_5/XI0/XI0_44/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_4 XI11_5/net21_11_ xsel_44_ XI11_5/XI0/XI0_44/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_3 XI11_5/net21_12_ xsel_44_ XI11_5/XI0/XI0_44/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_2 XI11_5/net21_13_ xsel_44_ XI11_5/XI0/XI0_44/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_1 XI11_5/net21_14_ xsel_44_ XI11_5/XI0/XI0_44/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN0_0 XI11_5/net21_15_ xsel_44_ XI11_5/XI0/XI0_44/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_15 XI11_5/XI0/XI0_44/d__15_ xsel_44_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_14 XI11_5/XI0/XI0_44/d__14_ xsel_44_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_13 XI11_5/XI0/XI0_44/d__13_ xsel_44_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_12 XI11_5/XI0/XI0_44/d__12_ xsel_44_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_11 XI11_5/XI0/XI0_44/d__11_ xsel_44_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_10 XI11_5/XI0/XI0_44/d__10_ xsel_44_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_9 XI11_5/XI0/XI0_44/d__9_ xsel_44_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_8 XI11_5/XI0/XI0_44/d__8_ xsel_44_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_7 XI11_5/XI0/XI0_44/d__7_ xsel_44_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_6 XI11_5/XI0/XI0_44/d__6_ xsel_44_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_5 XI11_5/XI0/XI0_44/d__5_ xsel_44_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_4 XI11_5/XI0/XI0_44/d__4_ xsel_44_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_3 XI11_5/XI0/XI0_44/d__3_ xsel_44_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_2 XI11_5/XI0/XI0_44/d__2_ xsel_44_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_1 XI11_5/XI0/XI0_44/d__1_ xsel_44_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_44/MN1_0 XI11_5/XI0/XI0_44/d__0_ xsel_44_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_15 XI11_5/net21_0_ xsel_43_ XI11_5/XI0/XI0_43/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_14 XI11_5/net21_1_ xsel_43_ XI11_5/XI0/XI0_43/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_13 XI11_5/net21_2_ xsel_43_ XI11_5/XI0/XI0_43/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_12 XI11_5/net21_3_ xsel_43_ XI11_5/XI0/XI0_43/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_11 XI11_5/net21_4_ xsel_43_ XI11_5/XI0/XI0_43/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_10 XI11_5/net21_5_ xsel_43_ XI11_5/XI0/XI0_43/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_9 XI11_5/net21_6_ xsel_43_ XI11_5/XI0/XI0_43/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_8 XI11_5/net21_7_ xsel_43_ XI11_5/XI0/XI0_43/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_7 XI11_5/net21_8_ xsel_43_ XI11_5/XI0/XI0_43/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_6 XI11_5/net21_9_ xsel_43_ XI11_5/XI0/XI0_43/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_5 XI11_5/net21_10_ xsel_43_ XI11_5/XI0/XI0_43/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_4 XI11_5/net21_11_ xsel_43_ XI11_5/XI0/XI0_43/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_3 XI11_5/net21_12_ xsel_43_ XI11_5/XI0/XI0_43/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_2 XI11_5/net21_13_ xsel_43_ XI11_5/XI0/XI0_43/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_1 XI11_5/net21_14_ xsel_43_ XI11_5/XI0/XI0_43/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN0_0 XI11_5/net21_15_ xsel_43_ XI11_5/XI0/XI0_43/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_15 XI11_5/XI0/XI0_43/d__15_ xsel_43_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_14 XI11_5/XI0/XI0_43/d__14_ xsel_43_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_13 XI11_5/XI0/XI0_43/d__13_ xsel_43_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_12 XI11_5/XI0/XI0_43/d__12_ xsel_43_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_11 XI11_5/XI0/XI0_43/d__11_ xsel_43_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_10 XI11_5/XI0/XI0_43/d__10_ xsel_43_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_9 XI11_5/XI0/XI0_43/d__9_ xsel_43_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_8 XI11_5/XI0/XI0_43/d__8_ xsel_43_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_7 XI11_5/XI0/XI0_43/d__7_ xsel_43_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_6 XI11_5/XI0/XI0_43/d__6_ xsel_43_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_5 XI11_5/XI0/XI0_43/d__5_ xsel_43_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_4 XI11_5/XI0/XI0_43/d__4_ xsel_43_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_3 XI11_5/XI0/XI0_43/d__3_ xsel_43_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_2 XI11_5/XI0/XI0_43/d__2_ xsel_43_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_1 XI11_5/XI0/XI0_43/d__1_ xsel_43_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_43/MN1_0 XI11_5/XI0/XI0_43/d__0_ xsel_43_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_15 XI11_5/net21_0_ xsel_42_ XI11_5/XI0/XI0_42/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_14 XI11_5/net21_1_ xsel_42_ XI11_5/XI0/XI0_42/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_13 XI11_5/net21_2_ xsel_42_ XI11_5/XI0/XI0_42/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_12 XI11_5/net21_3_ xsel_42_ XI11_5/XI0/XI0_42/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_11 XI11_5/net21_4_ xsel_42_ XI11_5/XI0/XI0_42/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_10 XI11_5/net21_5_ xsel_42_ XI11_5/XI0/XI0_42/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_9 XI11_5/net21_6_ xsel_42_ XI11_5/XI0/XI0_42/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_8 XI11_5/net21_7_ xsel_42_ XI11_5/XI0/XI0_42/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_7 XI11_5/net21_8_ xsel_42_ XI11_5/XI0/XI0_42/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_6 XI11_5/net21_9_ xsel_42_ XI11_5/XI0/XI0_42/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_5 XI11_5/net21_10_ xsel_42_ XI11_5/XI0/XI0_42/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_4 XI11_5/net21_11_ xsel_42_ XI11_5/XI0/XI0_42/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_3 XI11_5/net21_12_ xsel_42_ XI11_5/XI0/XI0_42/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_2 XI11_5/net21_13_ xsel_42_ XI11_5/XI0/XI0_42/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_1 XI11_5/net21_14_ xsel_42_ XI11_5/XI0/XI0_42/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN0_0 XI11_5/net21_15_ xsel_42_ XI11_5/XI0/XI0_42/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_15 XI11_5/XI0/XI0_42/d__15_ xsel_42_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_14 XI11_5/XI0/XI0_42/d__14_ xsel_42_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_13 XI11_5/XI0/XI0_42/d__13_ xsel_42_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_12 XI11_5/XI0/XI0_42/d__12_ xsel_42_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_11 XI11_5/XI0/XI0_42/d__11_ xsel_42_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_10 XI11_5/XI0/XI0_42/d__10_ xsel_42_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_9 XI11_5/XI0/XI0_42/d__9_ xsel_42_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_8 XI11_5/XI0/XI0_42/d__8_ xsel_42_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_7 XI11_5/XI0/XI0_42/d__7_ xsel_42_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_6 XI11_5/XI0/XI0_42/d__6_ xsel_42_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_5 XI11_5/XI0/XI0_42/d__5_ xsel_42_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_4 XI11_5/XI0/XI0_42/d__4_ xsel_42_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_3 XI11_5/XI0/XI0_42/d__3_ xsel_42_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_2 XI11_5/XI0/XI0_42/d__2_ xsel_42_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_1 XI11_5/XI0/XI0_42/d__1_ xsel_42_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_42/MN1_0 XI11_5/XI0/XI0_42/d__0_ xsel_42_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_15 XI11_5/net21_0_ xsel_41_ XI11_5/XI0/XI0_41/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_14 XI11_5/net21_1_ xsel_41_ XI11_5/XI0/XI0_41/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_13 XI11_5/net21_2_ xsel_41_ XI11_5/XI0/XI0_41/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_12 XI11_5/net21_3_ xsel_41_ XI11_5/XI0/XI0_41/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_11 XI11_5/net21_4_ xsel_41_ XI11_5/XI0/XI0_41/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_10 XI11_5/net21_5_ xsel_41_ XI11_5/XI0/XI0_41/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_9 XI11_5/net21_6_ xsel_41_ XI11_5/XI0/XI0_41/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_8 XI11_5/net21_7_ xsel_41_ XI11_5/XI0/XI0_41/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_7 XI11_5/net21_8_ xsel_41_ XI11_5/XI0/XI0_41/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_6 XI11_5/net21_9_ xsel_41_ XI11_5/XI0/XI0_41/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_5 XI11_5/net21_10_ xsel_41_ XI11_5/XI0/XI0_41/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_4 XI11_5/net21_11_ xsel_41_ XI11_5/XI0/XI0_41/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_3 XI11_5/net21_12_ xsel_41_ XI11_5/XI0/XI0_41/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_2 XI11_5/net21_13_ xsel_41_ XI11_5/XI0/XI0_41/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_1 XI11_5/net21_14_ xsel_41_ XI11_5/XI0/XI0_41/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN0_0 XI11_5/net21_15_ xsel_41_ XI11_5/XI0/XI0_41/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_15 XI11_5/XI0/XI0_41/d__15_ xsel_41_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_14 XI11_5/XI0/XI0_41/d__14_ xsel_41_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_13 XI11_5/XI0/XI0_41/d__13_ xsel_41_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_12 XI11_5/XI0/XI0_41/d__12_ xsel_41_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_11 XI11_5/XI0/XI0_41/d__11_ xsel_41_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_10 XI11_5/XI0/XI0_41/d__10_ xsel_41_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_9 XI11_5/XI0/XI0_41/d__9_ xsel_41_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_8 XI11_5/XI0/XI0_41/d__8_ xsel_41_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_7 XI11_5/XI0/XI0_41/d__7_ xsel_41_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_6 XI11_5/XI0/XI0_41/d__6_ xsel_41_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_5 XI11_5/XI0/XI0_41/d__5_ xsel_41_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_4 XI11_5/XI0/XI0_41/d__4_ xsel_41_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_3 XI11_5/XI0/XI0_41/d__3_ xsel_41_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_2 XI11_5/XI0/XI0_41/d__2_ xsel_41_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_1 XI11_5/XI0/XI0_41/d__1_ xsel_41_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_41/MN1_0 XI11_5/XI0/XI0_41/d__0_ xsel_41_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_15 XI11_5/net21_0_ xsel_40_ XI11_5/XI0/XI0_40/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_14 XI11_5/net21_1_ xsel_40_ XI11_5/XI0/XI0_40/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_13 XI11_5/net21_2_ xsel_40_ XI11_5/XI0/XI0_40/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_12 XI11_5/net21_3_ xsel_40_ XI11_5/XI0/XI0_40/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_11 XI11_5/net21_4_ xsel_40_ XI11_5/XI0/XI0_40/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_10 XI11_5/net21_5_ xsel_40_ XI11_5/XI0/XI0_40/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_9 XI11_5/net21_6_ xsel_40_ XI11_5/XI0/XI0_40/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_8 XI11_5/net21_7_ xsel_40_ XI11_5/XI0/XI0_40/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_7 XI11_5/net21_8_ xsel_40_ XI11_5/XI0/XI0_40/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_6 XI11_5/net21_9_ xsel_40_ XI11_5/XI0/XI0_40/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_5 XI11_5/net21_10_ xsel_40_ XI11_5/XI0/XI0_40/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_4 XI11_5/net21_11_ xsel_40_ XI11_5/XI0/XI0_40/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_3 XI11_5/net21_12_ xsel_40_ XI11_5/XI0/XI0_40/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_2 XI11_5/net21_13_ xsel_40_ XI11_5/XI0/XI0_40/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_1 XI11_5/net21_14_ xsel_40_ XI11_5/XI0/XI0_40/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN0_0 XI11_5/net21_15_ xsel_40_ XI11_5/XI0/XI0_40/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_15 XI11_5/XI0/XI0_40/d__15_ xsel_40_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_14 XI11_5/XI0/XI0_40/d__14_ xsel_40_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_13 XI11_5/XI0/XI0_40/d__13_ xsel_40_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_12 XI11_5/XI0/XI0_40/d__12_ xsel_40_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_11 XI11_5/XI0/XI0_40/d__11_ xsel_40_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_10 XI11_5/XI0/XI0_40/d__10_ xsel_40_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_9 XI11_5/XI0/XI0_40/d__9_ xsel_40_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_8 XI11_5/XI0/XI0_40/d__8_ xsel_40_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_7 XI11_5/XI0/XI0_40/d__7_ xsel_40_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_6 XI11_5/XI0/XI0_40/d__6_ xsel_40_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_5 XI11_5/XI0/XI0_40/d__5_ xsel_40_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_4 XI11_5/XI0/XI0_40/d__4_ xsel_40_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_3 XI11_5/XI0/XI0_40/d__3_ xsel_40_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_2 XI11_5/XI0/XI0_40/d__2_ xsel_40_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_1 XI11_5/XI0/XI0_40/d__1_ xsel_40_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_40/MN1_0 XI11_5/XI0/XI0_40/d__0_ xsel_40_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_15 XI11_5/net21_0_ xsel_39_ XI11_5/XI0/XI0_39/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_14 XI11_5/net21_1_ xsel_39_ XI11_5/XI0/XI0_39/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_13 XI11_5/net21_2_ xsel_39_ XI11_5/XI0/XI0_39/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_12 XI11_5/net21_3_ xsel_39_ XI11_5/XI0/XI0_39/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_11 XI11_5/net21_4_ xsel_39_ XI11_5/XI0/XI0_39/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_10 XI11_5/net21_5_ xsel_39_ XI11_5/XI0/XI0_39/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_9 XI11_5/net21_6_ xsel_39_ XI11_5/XI0/XI0_39/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_8 XI11_5/net21_7_ xsel_39_ XI11_5/XI0/XI0_39/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_7 XI11_5/net21_8_ xsel_39_ XI11_5/XI0/XI0_39/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_6 XI11_5/net21_9_ xsel_39_ XI11_5/XI0/XI0_39/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_5 XI11_5/net21_10_ xsel_39_ XI11_5/XI0/XI0_39/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_4 XI11_5/net21_11_ xsel_39_ XI11_5/XI0/XI0_39/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_3 XI11_5/net21_12_ xsel_39_ XI11_5/XI0/XI0_39/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_2 XI11_5/net21_13_ xsel_39_ XI11_5/XI0/XI0_39/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_1 XI11_5/net21_14_ xsel_39_ XI11_5/XI0/XI0_39/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN0_0 XI11_5/net21_15_ xsel_39_ XI11_5/XI0/XI0_39/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_15 XI11_5/XI0/XI0_39/d__15_ xsel_39_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_14 XI11_5/XI0/XI0_39/d__14_ xsel_39_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_13 XI11_5/XI0/XI0_39/d__13_ xsel_39_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_12 XI11_5/XI0/XI0_39/d__12_ xsel_39_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_11 XI11_5/XI0/XI0_39/d__11_ xsel_39_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_10 XI11_5/XI0/XI0_39/d__10_ xsel_39_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_9 XI11_5/XI0/XI0_39/d__9_ xsel_39_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_8 XI11_5/XI0/XI0_39/d__8_ xsel_39_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_7 XI11_5/XI0/XI0_39/d__7_ xsel_39_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_6 XI11_5/XI0/XI0_39/d__6_ xsel_39_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_5 XI11_5/XI0/XI0_39/d__5_ xsel_39_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_4 XI11_5/XI0/XI0_39/d__4_ xsel_39_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_3 XI11_5/XI0/XI0_39/d__3_ xsel_39_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_2 XI11_5/XI0/XI0_39/d__2_ xsel_39_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_1 XI11_5/XI0/XI0_39/d__1_ xsel_39_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_39/MN1_0 XI11_5/XI0/XI0_39/d__0_ xsel_39_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_15 XI11_5/net21_0_ xsel_38_ XI11_5/XI0/XI0_38/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_14 XI11_5/net21_1_ xsel_38_ XI11_5/XI0/XI0_38/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_13 XI11_5/net21_2_ xsel_38_ XI11_5/XI0/XI0_38/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_12 XI11_5/net21_3_ xsel_38_ XI11_5/XI0/XI0_38/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_11 XI11_5/net21_4_ xsel_38_ XI11_5/XI0/XI0_38/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_10 XI11_5/net21_5_ xsel_38_ XI11_5/XI0/XI0_38/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_9 XI11_5/net21_6_ xsel_38_ XI11_5/XI0/XI0_38/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_8 XI11_5/net21_7_ xsel_38_ XI11_5/XI0/XI0_38/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_7 XI11_5/net21_8_ xsel_38_ XI11_5/XI0/XI0_38/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_6 XI11_5/net21_9_ xsel_38_ XI11_5/XI0/XI0_38/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_5 XI11_5/net21_10_ xsel_38_ XI11_5/XI0/XI0_38/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_4 XI11_5/net21_11_ xsel_38_ XI11_5/XI0/XI0_38/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_3 XI11_5/net21_12_ xsel_38_ XI11_5/XI0/XI0_38/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_2 XI11_5/net21_13_ xsel_38_ XI11_5/XI0/XI0_38/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_1 XI11_5/net21_14_ xsel_38_ XI11_5/XI0/XI0_38/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN0_0 XI11_5/net21_15_ xsel_38_ XI11_5/XI0/XI0_38/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_15 XI11_5/XI0/XI0_38/d__15_ xsel_38_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_14 XI11_5/XI0/XI0_38/d__14_ xsel_38_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_13 XI11_5/XI0/XI0_38/d__13_ xsel_38_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_12 XI11_5/XI0/XI0_38/d__12_ xsel_38_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_11 XI11_5/XI0/XI0_38/d__11_ xsel_38_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_10 XI11_5/XI0/XI0_38/d__10_ xsel_38_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_9 XI11_5/XI0/XI0_38/d__9_ xsel_38_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_8 XI11_5/XI0/XI0_38/d__8_ xsel_38_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_7 XI11_5/XI0/XI0_38/d__7_ xsel_38_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_6 XI11_5/XI0/XI0_38/d__6_ xsel_38_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_5 XI11_5/XI0/XI0_38/d__5_ xsel_38_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_4 XI11_5/XI0/XI0_38/d__4_ xsel_38_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_3 XI11_5/XI0/XI0_38/d__3_ xsel_38_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_2 XI11_5/XI0/XI0_38/d__2_ xsel_38_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_1 XI11_5/XI0/XI0_38/d__1_ xsel_38_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_38/MN1_0 XI11_5/XI0/XI0_38/d__0_ xsel_38_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_15 XI11_5/net21_0_ xsel_37_ XI11_5/XI0/XI0_37/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_14 XI11_5/net21_1_ xsel_37_ XI11_5/XI0/XI0_37/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_13 XI11_5/net21_2_ xsel_37_ XI11_5/XI0/XI0_37/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_12 XI11_5/net21_3_ xsel_37_ XI11_5/XI0/XI0_37/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_11 XI11_5/net21_4_ xsel_37_ XI11_5/XI0/XI0_37/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_10 XI11_5/net21_5_ xsel_37_ XI11_5/XI0/XI0_37/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_9 XI11_5/net21_6_ xsel_37_ XI11_5/XI0/XI0_37/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_8 XI11_5/net21_7_ xsel_37_ XI11_5/XI0/XI0_37/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_7 XI11_5/net21_8_ xsel_37_ XI11_5/XI0/XI0_37/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_6 XI11_5/net21_9_ xsel_37_ XI11_5/XI0/XI0_37/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_5 XI11_5/net21_10_ xsel_37_ XI11_5/XI0/XI0_37/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_4 XI11_5/net21_11_ xsel_37_ XI11_5/XI0/XI0_37/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_3 XI11_5/net21_12_ xsel_37_ XI11_5/XI0/XI0_37/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_2 XI11_5/net21_13_ xsel_37_ XI11_5/XI0/XI0_37/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_1 XI11_5/net21_14_ xsel_37_ XI11_5/XI0/XI0_37/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN0_0 XI11_5/net21_15_ xsel_37_ XI11_5/XI0/XI0_37/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_15 XI11_5/XI0/XI0_37/d__15_ xsel_37_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_14 XI11_5/XI0/XI0_37/d__14_ xsel_37_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_13 XI11_5/XI0/XI0_37/d__13_ xsel_37_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_12 XI11_5/XI0/XI0_37/d__12_ xsel_37_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_11 XI11_5/XI0/XI0_37/d__11_ xsel_37_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_10 XI11_5/XI0/XI0_37/d__10_ xsel_37_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_9 XI11_5/XI0/XI0_37/d__9_ xsel_37_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_8 XI11_5/XI0/XI0_37/d__8_ xsel_37_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_7 XI11_5/XI0/XI0_37/d__7_ xsel_37_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_6 XI11_5/XI0/XI0_37/d__6_ xsel_37_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_5 XI11_5/XI0/XI0_37/d__5_ xsel_37_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_4 XI11_5/XI0/XI0_37/d__4_ xsel_37_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_3 XI11_5/XI0/XI0_37/d__3_ xsel_37_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_2 XI11_5/XI0/XI0_37/d__2_ xsel_37_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_1 XI11_5/XI0/XI0_37/d__1_ xsel_37_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_37/MN1_0 XI11_5/XI0/XI0_37/d__0_ xsel_37_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_15 XI11_5/net21_0_ xsel_36_ XI11_5/XI0/XI0_36/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_14 XI11_5/net21_1_ xsel_36_ XI11_5/XI0/XI0_36/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_13 XI11_5/net21_2_ xsel_36_ XI11_5/XI0/XI0_36/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_12 XI11_5/net21_3_ xsel_36_ XI11_5/XI0/XI0_36/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_11 XI11_5/net21_4_ xsel_36_ XI11_5/XI0/XI0_36/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_10 XI11_5/net21_5_ xsel_36_ XI11_5/XI0/XI0_36/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_9 XI11_5/net21_6_ xsel_36_ XI11_5/XI0/XI0_36/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_8 XI11_5/net21_7_ xsel_36_ XI11_5/XI0/XI0_36/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_7 XI11_5/net21_8_ xsel_36_ XI11_5/XI0/XI0_36/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_6 XI11_5/net21_9_ xsel_36_ XI11_5/XI0/XI0_36/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_5 XI11_5/net21_10_ xsel_36_ XI11_5/XI0/XI0_36/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_4 XI11_5/net21_11_ xsel_36_ XI11_5/XI0/XI0_36/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_3 XI11_5/net21_12_ xsel_36_ XI11_5/XI0/XI0_36/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_2 XI11_5/net21_13_ xsel_36_ XI11_5/XI0/XI0_36/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_1 XI11_5/net21_14_ xsel_36_ XI11_5/XI0/XI0_36/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN0_0 XI11_5/net21_15_ xsel_36_ XI11_5/XI0/XI0_36/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_15 XI11_5/XI0/XI0_36/d__15_ xsel_36_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_14 XI11_5/XI0/XI0_36/d__14_ xsel_36_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_13 XI11_5/XI0/XI0_36/d__13_ xsel_36_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_12 XI11_5/XI0/XI0_36/d__12_ xsel_36_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_11 XI11_5/XI0/XI0_36/d__11_ xsel_36_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_10 XI11_5/XI0/XI0_36/d__10_ xsel_36_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_9 XI11_5/XI0/XI0_36/d__9_ xsel_36_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_8 XI11_5/XI0/XI0_36/d__8_ xsel_36_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_7 XI11_5/XI0/XI0_36/d__7_ xsel_36_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_6 XI11_5/XI0/XI0_36/d__6_ xsel_36_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_5 XI11_5/XI0/XI0_36/d__5_ xsel_36_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_4 XI11_5/XI0/XI0_36/d__4_ xsel_36_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_3 XI11_5/XI0/XI0_36/d__3_ xsel_36_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_2 XI11_5/XI0/XI0_36/d__2_ xsel_36_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_1 XI11_5/XI0/XI0_36/d__1_ xsel_36_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_36/MN1_0 XI11_5/XI0/XI0_36/d__0_ xsel_36_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_15 XI11_5/net21_0_ xsel_35_ XI11_5/XI0/XI0_35/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_14 XI11_5/net21_1_ xsel_35_ XI11_5/XI0/XI0_35/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_13 XI11_5/net21_2_ xsel_35_ XI11_5/XI0/XI0_35/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_12 XI11_5/net21_3_ xsel_35_ XI11_5/XI0/XI0_35/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_11 XI11_5/net21_4_ xsel_35_ XI11_5/XI0/XI0_35/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_10 XI11_5/net21_5_ xsel_35_ XI11_5/XI0/XI0_35/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_9 XI11_5/net21_6_ xsel_35_ XI11_5/XI0/XI0_35/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_8 XI11_5/net21_7_ xsel_35_ XI11_5/XI0/XI0_35/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_7 XI11_5/net21_8_ xsel_35_ XI11_5/XI0/XI0_35/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_6 XI11_5/net21_9_ xsel_35_ XI11_5/XI0/XI0_35/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_5 XI11_5/net21_10_ xsel_35_ XI11_5/XI0/XI0_35/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_4 XI11_5/net21_11_ xsel_35_ XI11_5/XI0/XI0_35/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_3 XI11_5/net21_12_ xsel_35_ XI11_5/XI0/XI0_35/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_2 XI11_5/net21_13_ xsel_35_ XI11_5/XI0/XI0_35/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_1 XI11_5/net21_14_ xsel_35_ XI11_5/XI0/XI0_35/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN0_0 XI11_5/net21_15_ xsel_35_ XI11_5/XI0/XI0_35/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_15 XI11_5/XI0/XI0_35/d__15_ xsel_35_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_14 XI11_5/XI0/XI0_35/d__14_ xsel_35_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_13 XI11_5/XI0/XI0_35/d__13_ xsel_35_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_12 XI11_5/XI0/XI0_35/d__12_ xsel_35_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_11 XI11_5/XI0/XI0_35/d__11_ xsel_35_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_10 XI11_5/XI0/XI0_35/d__10_ xsel_35_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_9 XI11_5/XI0/XI0_35/d__9_ xsel_35_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_8 XI11_5/XI0/XI0_35/d__8_ xsel_35_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_7 XI11_5/XI0/XI0_35/d__7_ xsel_35_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_6 XI11_5/XI0/XI0_35/d__6_ xsel_35_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_5 XI11_5/XI0/XI0_35/d__5_ xsel_35_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_4 XI11_5/XI0/XI0_35/d__4_ xsel_35_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_3 XI11_5/XI0/XI0_35/d__3_ xsel_35_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_2 XI11_5/XI0/XI0_35/d__2_ xsel_35_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_1 XI11_5/XI0/XI0_35/d__1_ xsel_35_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_35/MN1_0 XI11_5/XI0/XI0_35/d__0_ xsel_35_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_15 XI11_5/net21_0_ xsel_34_ XI11_5/XI0/XI0_34/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_14 XI11_5/net21_1_ xsel_34_ XI11_5/XI0/XI0_34/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_13 XI11_5/net21_2_ xsel_34_ XI11_5/XI0/XI0_34/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_12 XI11_5/net21_3_ xsel_34_ XI11_5/XI0/XI0_34/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_11 XI11_5/net21_4_ xsel_34_ XI11_5/XI0/XI0_34/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_10 XI11_5/net21_5_ xsel_34_ XI11_5/XI0/XI0_34/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_9 XI11_5/net21_6_ xsel_34_ XI11_5/XI0/XI0_34/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_8 XI11_5/net21_7_ xsel_34_ XI11_5/XI0/XI0_34/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_7 XI11_5/net21_8_ xsel_34_ XI11_5/XI0/XI0_34/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_6 XI11_5/net21_9_ xsel_34_ XI11_5/XI0/XI0_34/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_5 XI11_5/net21_10_ xsel_34_ XI11_5/XI0/XI0_34/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_4 XI11_5/net21_11_ xsel_34_ XI11_5/XI0/XI0_34/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_3 XI11_5/net21_12_ xsel_34_ XI11_5/XI0/XI0_34/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_2 XI11_5/net21_13_ xsel_34_ XI11_5/XI0/XI0_34/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_1 XI11_5/net21_14_ xsel_34_ XI11_5/XI0/XI0_34/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN0_0 XI11_5/net21_15_ xsel_34_ XI11_5/XI0/XI0_34/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_15 XI11_5/XI0/XI0_34/d__15_ xsel_34_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_14 XI11_5/XI0/XI0_34/d__14_ xsel_34_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_13 XI11_5/XI0/XI0_34/d__13_ xsel_34_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_12 XI11_5/XI0/XI0_34/d__12_ xsel_34_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_11 XI11_5/XI0/XI0_34/d__11_ xsel_34_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_10 XI11_5/XI0/XI0_34/d__10_ xsel_34_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_9 XI11_5/XI0/XI0_34/d__9_ xsel_34_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_8 XI11_5/XI0/XI0_34/d__8_ xsel_34_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_7 XI11_5/XI0/XI0_34/d__7_ xsel_34_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_6 XI11_5/XI0/XI0_34/d__6_ xsel_34_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_5 XI11_5/XI0/XI0_34/d__5_ xsel_34_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_4 XI11_5/XI0/XI0_34/d__4_ xsel_34_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_3 XI11_5/XI0/XI0_34/d__3_ xsel_34_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_2 XI11_5/XI0/XI0_34/d__2_ xsel_34_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_1 XI11_5/XI0/XI0_34/d__1_ xsel_34_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_34/MN1_0 XI11_5/XI0/XI0_34/d__0_ xsel_34_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_15 XI11_5/net21_0_ xsel_33_ XI11_5/XI0/XI0_33/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_14 XI11_5/net21_1_ xsel_33_ XI11_5/XI0/XI0_33/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_13 XI11_5/net21_2_ xsel_33_ XI11_5/XI0/XI0_33/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_12 XI11_5/net21_3_ xsel_33_ XI11_5/XI0/XI0_33/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_11 XI11_5/net21_4_ xsel_33_ XI11_5/XI0/XI0_33/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_10 XI11_5/net21_5_ xsel_33_ XI11_5/XI0/XI0_33/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_9 XI11_5/net21_6_ xsel_33_ XI11_5/XI0/XI0_33/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_8 XI11_5/net21_7_ xsel_33_ XI11_5/XI0/XI0_33/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_7 XI11_5/net21_8_ xsel_33_ XI11_5/XI0/XI0_33/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_6 XI11_5/net21_9_ xsel_33_ XI11_5/XI0/XI0_33/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_5 XI11_5/net21_10_ xsel_33_ XI11_5/XI0/XI0_33/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_4 XI11_5/net21_11_ xsel_33_ XI11_5/XI0/XI0_33/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_3 XI11_5/net21_12_ xsel_33_ XI11_5/XI0/XI0_33/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_2 XI11_5/net21_13_ xsel_33_ XI11_5/XI0/XI0_33/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_1 XI11_5/net21_14_ xsel_33_ XI11_5/XI0/XI0_33/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN0_0 XI11_5/net21_15_ xsel_33_ XI11_5/XI0/XI0_33/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_15 XI11_5/XI0/XI0_33/d__15_ xsel_33_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_14 XI11_5/XI0/XI0_33/d__14_ xsel_33_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_13 XI11_5/XI0/XI0_33/d__13_ xsel_33_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_12 XI11_5/XI0/XI0_33/d__12_ xsel_33_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_11 XI11_5/XI0/XI0_33/d__11_ xsel_33_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_10 XI11_5/XI0/XI0_33/d__10_ xsel_33_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_9 XI11_5/XI0/XI0_33/d__9_ xsel_33_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_8 XI11_5/XI0/XI0_33/d__8_ xsel_33_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_7 XI11_5/XI0/XI0_33/d__7_ xsel_33_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_6 XI11_5/XI0/XI0_33/d__6_ xsel_33_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_5 XI11_5/XI0/XI0_33/d__5_ xsel_33_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_4 XI11_5/XI0/XI0_33/d__4_ xsel_33_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_3 XI11_5/XI0/XI0_33/d__3_ xsel_33_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_2 XI11_5/XI0/XI0_33/d__2_ xsel_33_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_1 XI11_5/XI0/XI0_33/d__1_ xsel_33_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_33/MN1_0 XI11_5/XI0/XI0_33/d__0_ xsel_33_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_15 XI11_5/net21_0_ xsel_32_ XI11_5/XI0/XI0_32/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_14 XI11_5/net21_1_ xsel_32_ XI11_5/XI0/XI0_32/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_13 XI11_5/net21_2_ xsel_32_ XI11_5/XI0/XI0_32/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_12 XI11_5/net21_3_ xsel_32_ XI11_5/XI0/XI0_32/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_11 XI11_5/net21_4_ xsel_32_ XI11_5/XI0/XI0_32/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_10 XI11_5/net21_5_ xsel_32_ XI11_5/XI0/XI0_32/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_9 XI11_5/net21_6_ xsel_32_ XI11_5/XI0/XI0_32/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_8 XI11_5/net21_7_ xsel_32_ XI11_5/XI0/XI0_32/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_7 XI11_5/net21_8_ xsel_32_ XI11_5/XI0/XI0_32/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_6 XI11_5/net21_9_ xsel_32_ XI11_5/XI0/XI0_32/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_5 XI11_5/net21_10_ xsel_32_ XI11_5/XI0/XI0_32/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_4 XI11_5/net21_11_ xsel_32_ XI11_5/XI0/XI0_32/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_3 XI11_5/net21_12_ xsel_32_ XI11_5/XI0/XI0_32/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_2 XI11_5/net21_13_ xsel_32_ XI11_5/XI0/XI0_32/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_1 XI11_5/net21_14_ xsel_32_ XI11_5/XI0/XI0_32/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN0_0 XI11_5/net21_15_ xsel_32_ XI11_5/XI0/XI0_32/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_15 XI11_5/XI0/XI0_32/d__15_ xsel_32_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_14 XI11_5/XI0/XI0_32/d__14_ xsel_32_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_13 XI11_5/XI0/XI0_32/d__13_ xsel_32_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_12 XI11_5/XI0/XI0_32/d__12_ xsel_32_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_11 XI11_5/XI0/XI0_32/d__11_ xsel_32_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_10 XI11_5/XI0/XI0_32/d__10_ xsel_32_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_9 XI11_5/XI0/XI0_32/d__9_ xsel_32_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_8 XI11_5/XI0/XI0_32/d__8_ xsel_32_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_7 XI11_5/XI0/XI0_32/d__7_ xsel_32_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_6 XI11_5/XI0/XI0_32/d__6_ xsel_32_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_5 XI11_5/XI0/XI0_32/d__5_ xsel_32_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_4 XI11_5/XI0/XI0_32/d__4_ xsel_32_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_3 XI11_5/XI0/XI0_32/d__3_ xsel_32_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_2 XI11_5/XI0/XI0_32/d__2_ xsel_32_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_1 XI11_5/XI0/XI0_32/d__1_ xsel_32_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_32/MN1_0 XI11_5/XI0/XI0_32/d__0_ xsel_32_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_15 XI11_5/net21_0_ xsel_31_ XI11_5/XI0/XI0_31/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_14 XI11_5/net21_1_ xsel_31_ XI11_5/XI0/XI0_31/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_13 XI11_5/net21_2_ xsel_31_ XI11_5/XI0/XI0_31/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_12 XI11_5/net21_3_ xsel_31_ XI11_5/XI0/XI0_31/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_11 XI11_5/net21_4_ xsel_31_ XI11_5/XI0/XI0_31/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_10 XI11_5/net21_5_ xsel_31_ XI11_5/XI0/XI0_31/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_9 XI11_5/net21_6_ xsel_31_ XI11_5/XI0/XI0_31/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_8 XI11_5/net21_7_ xsel_31_ XI11_5/XI0/XI0_31/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_7 XI11_5/net21_8_ xsel_31_ XI11_5/XI0/XI0_31/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_6 XI11_5/net21_9_ xsel_31_ XI11_5/XI0/XI0_31/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_5 XI11_5/net21_10_ xsel_31_ XI11_5/XI0/XI0_31/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_4 XI11_5/net21_11_ xsel_31_ XI11_5/XI0/XI0_31/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_3 XI11_5/net21_12_ xsel_31_ XI11_5/XI0/XI0_31/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_2 XI11_5/net21_13_ xsel_31_ XI11_5/XI0/XI0_31/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_1 XI11_5/net21_14_ xsel_31_ XI11_5/XI0/XI0_31/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN0_0 XI11_5/net21_15_ xsel_31_ XI11_5/XI0/XI0_31/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_15 XI11_5/XI0/XI0_31/d__15_ xsel_31_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_14 XI11_5/XI0/XI0_31/d__14_ xsel_31_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_13 XI11_5/XI0/XI0_31/d__13_ xsel_31_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_12 XI11_5/XI0/XI0_31/d__12_ xsel_31_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_11 XI11_5/XI0/XI0_31/d__11_ xsel_31_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_10 XI11_5/XI0/XI0_31/d__10_ xsel_31_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_9 XI11_5/XI0/XI0_31/d__9_ xsel_31_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_8 XI11_5/XI0/XI0_31/d__8_ xsel_31_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_7 XI11_5/XI0/XI0_31/d__7_ xsel_31_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_6 XI11_5/XI0/XI0_31/d__6_ xsel_31_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_5 XI11_5/XI0/XI0_31/d__5_ xsel_31_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_4 XI11_5/XI0/XI0_31/d__4_ xsel_31_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_3 XI11_5/XI0/XI0_31/d__3_ xsel_31_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_2 XI11_5/XI0/XI0_31/d__2_ xsel_31_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_1 XI11_5/XI0/XI0_31/d__1_ xsel_31_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_31/MN1_0 XI11_5/XI0/XI0_31/d__0_ xsel_31_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_15 XI11_5/net21_0_ xsel_30_ XI11_5/XI0/XI0_30/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_14 XI11_5/net21_1_ xsel_30_ XI11_5/XI0/XI0_30/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_13 XI11_5/net21_2_ xsel_30_ XI11_5/XI0/XI0_30/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_12 XI11_5/net21_3_ xsel_30_ XI11_5/XI0/XI0_30/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_11 XI11_5/net21_4_ xsel_30_ XI11_5/XI0/XI0_30/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_10 XI11_5/net21_5_ xsel_30_ XI11_5/XI0/XI0_30/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_9 XI11_5/net21_6_ xsel_30_ XI11_5/XI0/XI0_30/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_8 XI11_5/net21_7_ xsel_30_ XI11_5/XI0/XI0_30/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_7 XI11_5/net21_8_ xsel_30_ XI11_5/XI0/XI0_30/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_6 XI11_5/net21_9_ xsel_30_ XI11_5/XI0/XI0_30/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_5 XI11_5/net21_10_ xsel_30_ XI11_5/XI0/XI0_30/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_4 XI11_5/net21_11_ xsel_30_ XI11_5/XI0/XI0_30/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_3 XI11_5/net21_12_ xsel_30_ XI11_5/XI0/XI0_30/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_2 XI11_5/net21_13_ xsel_30_ XI11_5/XI0/XI0_30/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_1 XI11_5/net21_14_ xsel_30_ XI11_5/XI0/XI0_30/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN0_0 XI11_5/net21_15_ xsel_30_ XI11_5/XI0/XI0_30/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_15 XI11_5/XI0/XI0_30/d__15_ xsel_30_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_14 XI11_5/XI0/XI0_30/d__14_ xsel_30_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_13 XI11_5/XI0/XI0_30/d__13_ xsel_30_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_12 XI11_5/XI0/XI0_30/d__12_ xsel_30_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_11 XI11_5/XI0/XI0_30/d__11_ xsel_30_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_10 XI11_5/XI0/XI0_30/d__10_ xsel_30_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_9 XI11_5/XI0/XI0_30/d__9_ xsel_30_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_8 XI11_5/XI0/XI0_30/d__8_ xsel_30_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_7 XI11_5/XI0/XI0_30/d__7_ xsel_30_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_6 XI11_5/XI0/XI0_30/d__6_ xsel_30_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_5 XI11_5/XI0/XI0_30/d__5_ xsel_30_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_4 XI11_5/XI0/XI0_30/d__4_ xsel_30_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_3 XI11_5/XI0/XI0_30/d__3_ xsel_30_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_2 XI11_5/XI0/XI0_30/d__2_ xsel_30_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_1 XI11_5/XI0/XI0_30/d__1_ xsel_30_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_30/MN1_0 XI11_5/XI0/XI0_30/d__0_ xsel_30_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_15 XI11_5/net21_0_ xsel_29_ XI11_5/XI0/XI0_29/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_14 XI11_5/net21_1_ xsel_29_ XI11_5/XI0/XI0_29/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_13 XI11_5/net21_2_ xsel_29_ XI11_5/XI0/XI0_29/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_12 XI11_5/net21_3_ xsel_29_ XI11_5/XI0/XI0_29/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_11 XI11_5/net21_4_ xsel_29_ XI11_5/XI0/XI0_29/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_10 XI11_5/net21_5_ xsel_29_ XI11_5/XI0/XI0_29/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_9 XI11_5/net21_6_ xsel_29_ XI11_5/XI0/XI0_29/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_8 XI11_5/net21_7_ xsel_29_ XI11_5/XI0/XI0_29/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_7 XI11_5/net21_8_ xsel_29_ XI11_5/XI0/XI0_29/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_6 XI11_5/net21_9_ xsel_29_ XI11_5/XI0/XI0_29/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_5 XI11_5/net21_10_ xsel_29_ XI11_5/XI0/XI0_29/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_4 XI11_5/net21_11_ xsel_29_ XI11_5/XI0/XI0_29/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_3 XI11_5/net21_12_ xsel_29_ XI11_5/XI0/XI0_29/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_2 XI11_5/net21_13_ xsel_29_ XI11_5/XI0/XI0_29/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_1 XI11_5/net21_14_ xsel_29_ XI11_5/XI0/XI0_29/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN0_0 XI11_5/net21_15_ xsel_29_ XI11_5/XI0/XI0_29/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_15 XI11_5/XI0/XI0_29/d__15_ xsel_29_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_14 XI11_5/XI0/XI0_29/d__14_ xsel_29_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_13 XI11_5/XI0/XI0_29/d__13_ xsel_29_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_12 XI11_5/XI0/XI0_29/d__12_ xsel_29_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_11 XI11_5/XI0/XI0_29/d__11_ xsel_29_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_10 XI11_5/XI0/XI0_29/d__10_ xsel_29_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_9 XI11_5/XI0/XI0_29/d__9_ xsel_29_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_8 XI11_5/XI0/XI0_29/d__8_ xsel_29_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_7 XI11_5/XI0/XI0_29/d__7_ xsel_29_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_6 XI11_5/XI0/XI0_29/d__6_ xsel_29_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_5 XI11_5/XI0/XI0_29/d__5_ xsel_29_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_4 XI11_5/XI0/XI0_29/d__4_ xsel_29_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_3 XI11_5/XI0/XI0_29/d__3_ xsel_29_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_2 XI11_5/XI0/XI0_29/d__2_ xsel_29_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_1 XI11_5/XI0/XI0_29/d__1_ xsel_29_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_29/MN1_0 XI11_5/XI0/XI0_29/d__0_ xsel_29_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_15 XI11_5/net21_0_ xsel_28_ XI11_5/XI0/XI0_28/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_14 XI11_5/net21_1_ xsel_28_ XI11_5/XI0/XI0_28/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_13 XI11_5/net21_2_ xsel_28_ XI11_5/XI0/XI0_28/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_12 XI11_5/net21_3_ xsel_28_ XI11_5/XI0/XI0_28/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_11 XI11_5/net21_4_ xsel_28_ XI11_5/XI0/XI0_28/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_10 XI11_5/net21_5_ xsel_28_ XI11_5/XI0/XI0_28/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_9 XI11_5/net21_6_ xsel_28_ XI11_5/XI0/XI0_28/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_8 XI11_5/net21_7_ xsel_28_ XI11_5/XI0/XI0_28/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_7 XI11_5/net21_8_ xsel_28_ XI11_5/XI0/XI0_28/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_6 XI11_5/net21_9_ xsel_28_ XI11_5/XI0/XI0_28/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_5 XI11_5/net21_10_ xsel_28_ XI11_5/XI0/XI0_28/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_4 XI11_5/net21_11_ xsel_28_ XI11_5/XI0/XI0_28/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_3 XI11_5/net21_12_ xsel_28_ XI11_5/XI0/XI0_28/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_2 XI11_5/net21_13_ xsel_28_ XI11_5/XI0/XI0_28/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_1 XI11_5/net21_14_ xsel_28_ XI11_5/XI0/XI0_28/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN0_0 XI11_5/net21_15_ xsel_28_ XI11_5/XI0/XI0_28/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_15 XI11_5/XI0/XI0_28/d__15_ xsel_28_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_14 XI11_5/XI0/XI0_28/d__14_ xsel_28_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_13 XI11_5/XI0/XI0_28/d__13_ xsel_28_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_12 XI11_5/XI0/XI0_28/d__12_ xsel_28_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_11 XI11_5/XI0/XI0_28/d__11_ xsel_28_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_10 XI11_5/XI0/XI0_28/d__10_ xsel_28_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_9 XI11_5/XI0/XI0_28/d__9_ xsel_28_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_8 XI11_5/XI0/XI0_28/d__8_ xsel_28_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_7 XI11_5/XI0/XI0_28/d__7_ xsel_28_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_6 XI11_5/XI0/XI0_28/d__6_ xsel_28_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_5 XI11_5/XI0/XI0_28/d__5_ xsel_28_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_4 XI11_5/XI0/XI0_28/d__4_ xsel_28_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_3 XI11_5/XI0/XI0_28/d__3_ xsel_28_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_2 XI11_5/XI0/XI0_28/d__2_ xsel_28_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_1 XI11_5/XI0/XI0_28/d__1_ xsel_28_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_28/MN1_0 XI11_5/XI0/XI0_28/d__0_ xsel_28_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_15 XI11_5/net21_0_ xsel_27_ XI11_5/XI0/XI0_27/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_14 XI11_5/net21_1_ xsel_27_ XI11_5/XI0/XI0_27/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_13 XI11_5/net21_2_ xsel_27_ XI11_5/XI0/XI0_27/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_12 XI11_5/net21_3_ xsel_27_ XI11_5/XI0/XI0_27/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_11 XI11_5/net21_4_ xsel_27_ XI11_5/XI0/XI0_27/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_10 XI11_5/net21_5_ xsel_27_ XI11_5/XI0/XI0_27/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_9 XI11_5/net21_6_ xsel_27_ XI11_5/XI0/XI0_27/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_8 XI11_5/net21_7_ xsel_27_ XI11_5/XI0/XI0_27/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_7 XI11_5/net21_8_ xsel_27_ XI11_5/XI0/XI0_27/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_6 XI11_5/net21_9_ xsel_27_ XI11_5/XI0/XI0_27/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_5 XI11_5/net21_10_ xsel_27_ XI11_5/XI0/XI0_27/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_4 XI11_5/net21_11_ xsel_27_ XI11_5/XI0/XI0_27/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_3 XI11_5/net21_12_ xsel_27_ XI11_5/XI0/XI0_27/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_2 XI11_5/net21_13_ xsel_27_ XI11_5/XI0/XI0_27/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_1 XI11_5/net21_14_ xsel_27_ XI11_5/XI0/XI0_27/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN0_0 XI11_5/net21_15_ xsel_27_ XI11_5/XI0/XI0_27/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_15 XI11_5/XI0/XI0_27/d__15_ xsel_27_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_14 XI11_5/XI0/XI0_27/d__14_ xsel_27_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_13 XI11_5/XI0/XI0_27/d__13_ xsel_27_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_12 XI11_5/XI0/XI0_27/d__12_ xsel_27_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_11 XI11_5/XI0/XI0_27/d__11_ xsel_27_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_10 XI11_5/XI0/XI0_27/d__10_ xsel_27_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_9 XI11_5/XI0/XI0_27/d__9_ xsel_27_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_8 XI11_5/XI0/XI0_27/d__8_ xsel_27_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_7 XI11_5/XI0/XI0_27/d__7_ xsel_27_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_6 XI11_5/XI0/XI0_27/d__6_ xsel_27_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_5 XI11_5/XI0/XI0_27/d__5_ xsel_27_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_4 XI11_5/XI0/XI0_27/d__4_ xsel_27_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_3 XI11_5/XI0/XI0_27/d__3_ xsel_27_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_2 XI11_5/XI0/XI0_27/d__2_ xsel_27_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_1 XI11_5/XI0/XI0_27/d__1_ xsel_27_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_27/MN1_0 XI11_5/XI0/XI0_27/d__0_ xsel_27_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_15 XI11_5/net21_0_ xsel_26_ XI11_5/XI0/XI0_26/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_14 XI11_5/net21_1_ xsel_26_ XI11_5/XI0/XI0_26/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_13 XI11_5/net21_2_ xsel_26_ XI11_5/XI0/XI0_26/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_12 XI11_5/net21_3_ xsel_26_ XI11_5/XI0/XI0_26/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_11 XI11_5/net21_4_ xsel_26_ XI11_5/XI0/XI0_26/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_10 XI11_5/net21_5_ xsel_26_ XI11_5/XI0/XI0_26/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_9 XI11_5/net21_6_ xsel_26_ XI11_5/XI0/XI0_26/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_8 XI11_5/net21_7_ xsel_26_ XI11_5/XI0/XI0_26/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_7 XI11_5/net21_8_ xsel_26_ XI11_5/XI0/XI0_26/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_6 XI11_5/net21_9_ xsel_26_ XI11_5/XI0/XI0_26/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_5 XI11_5/net21_10_ xsel_26_ XI11_5/XI0/XI0_26/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_4 XI11_5/net21_11_ xsel_26_ XI11_5/XI0/XI0_26/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_3 XI11_5/net21_12_ xsel_26_ XI11_5/XI0/XI0_26/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_2 XI11_5/net21_13_ xsel_26_ XI11_5/XI0/XI0_26/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_1 XI11_5/net21_14_ xsel_26_ XI11_5/XI0/XI0_26/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN0_0 XI11_5/net21_15_ xsel_26_ XI11_5/XI0/XI0_26/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_15 XI11_5/XI0/XI0_26/d__15_ xsel_26_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_14 XI11_5/XI0/XI0_26/d__14_ xsel_26_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_13 XI11_5/XI0/XI0_26/d__13_ xsel_26_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_12 XI11_5/XI0/XI0_26/d__12_ xsel_26_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_11 XI11_5/XI0/XI0_26/d__11_ xsel_26_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_10 XI11_5/XI0/XI0_26/d__10_ xsel_26_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_9 XI11_5/XI0/XI0_26/d__9_ xsel_26_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_8 XI11_5/XI0/XI0_26/d__8_ xsel_26_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_7 XI11_5/XI0/XI0_26/d__7_ xsel_26_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_6 XI11_5/XI0/XI0_26/d__6_ xsel_26_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_5 XI11_5/XI0/XI0_26/d__5_ xsel_26_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_4 XI11_5/XI0/XI0_26/d__4_ xsel_26_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_3 XI11_5/XI0/XI0_26/d__3_ xsel_26_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_2 XI11_5/XI0/XI0_26/d__2_ xsel_26_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_1 XI11_5/XI0/XI0_26/d__1_ xsel_26_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_26/MN1_0 XI11_5/XI0/XI0_26/d__0_ xsel_26_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_15 XI11_5/net21_0_ xsel_25_ XI11_5/XI0/XI0_25/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_14 XI11_5/net21_1_ xsel_25_ XI11_5/XI0/XI0_25/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_13 XI11_5/net21_2_ xsel_25_ XI11_5/XI0/XI0_25/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_12 XI11_5/net21_3_ xsel_25_ XI11_5/XI0/XI0_25/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_11 XI11_5/net21_4_ xsel_25_ XI11_5/XI0/XI0_25/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_10 XI11_5/net21_5_ xsel_25_ XI11_5/XI0/XI0_25/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_9 XI11_5/net21_6_ xsel_25_ XI11_5/XI0/XI0_25/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_8 XI11_5/net21_7_ xsel_25_ XI11_5/XI0/XI0_25/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_7 XI11_5/net21_8_ xsel_25_ XI11_5/XI0/XI0_25/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_6 XI11_5/net21_9_ xsel_25_ XI11_5/XI0/XI0_25/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_5 XI11_5/net21_10_ xsel_25_ XI11_5/XI0/XI0_25/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_4 XI11_5/net21_11_ xsel_25_ XI11_5/XI0/XI0_25/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_3 XI11_5/net21_12_ xsel_25_ XI11_5/XI0/XI0_25/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_2 XI11_5/net21_13_ xsel_25_ XI11_5/XI0/XI0_25/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_1 XI11_5/net21_14_ xsel_25_ XI11_5/XI0/XI0_25/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN0_0 XI11_5/net21_15_ xsel_25_ XI11_5/XI0/XI0_25/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_15 XI11_5/XI0/XI0_25/d__15_ xsel_25_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_14 XI11_5/XI0/XI0_25/d__14_ xsel_25_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_13 XI11_5/XI0/XI0_25/d__13_ xsel_25_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_12 XI11_5/XI0/XI0_25/d__12_ xsel_25_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_11 XI11_5/XI0/XI0_25/d__11_ xsel_25_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_10 XI11_5/XI0/XI0_25/d__10_ xsel_25_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_9 XI11_5/XI0/XI0_25/d__9_ xsel_25_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_8 XI11_5/XI0/XI0_25/d__8_ xsel_25_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_7 XI11_5/XI0/XI0_25/d__7_ xsel_25_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_6 XI11_5/XI0/XI0_25/d__6_ xsel_25_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_5 XI11_5/XI0/XI0_25/d__5_ xsel_25_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_4 XI11_5/XI0/XI0_25/d__4_ xsel_25_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_3 XI11_5/XI0/XI0_25/d__3_ xsel_25_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_2 XI11_5/XI0/XI0_25/d__2_ xsel_25_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_1 XI11_5/XI0/XI0_25/d__1_ xsel_25_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_25/MN1_0 XI11_5/XI0/XI0_25/d__0_ xsel_25_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_15 XI11_5/net21_0_ xsel_24_ XI11_5/XI0/XI0_24/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_14 XI11_5/net21_1_ xsel_24_ XI11_5/XI0/XI0_24/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_13 XI11_5/net21_2_ xsel_24_ XI11_5/XI0/XI0_24/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_12 XI11_5/net21_3_ xsel_24_ XI11_5/XI0/XI0_24/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_11 XI11_5/net21_4_ xsel_24_ XI11_5/XI0/XI0_24/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_10 XI11_5/net21_5_ xsel_24_ XI11_5/XI0/XI0_24/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_9 XI11_5/net21_6_ xsel_24_ XI11_5/XI0/XI0_24/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_8 XI11_5/net21_7_ xsel_24_ XI11_5/XI0/XI0_24/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_7 XI11_5/net21_8_ xsel_24_ XI11_5/XI0/XI0_24/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_6 XI11_5/net21_9_ xsel_24_ XI11_5/XI0/XI0_24/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_5 XI11_5/net21_10_ xsel_24_ XI11_5/XI0/XI0_24/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_4 XI11_5/net21_11_ xsel_24_ XI11_5/XI0/XI0_24/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_3 XI11_5/net21_12_ xsel_24_ XI11_5/XI0/XI0_24/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_2 XI11_5/net21_13_ xsel_24_ XI11_5/XI0/XI0_24/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_1 XI11_5/net21_14_ xsel_24_ XI11_5/XI0/XI0_24/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN0_0 XI11_5/net21_15_ xsel_24_ XI11_5/XI0/XI0_24/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_15 XI11_5/XI0/XI0_24/d__15_ xsel_24_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_14 XI11_5/XI0/XI0_24/d__14_ xsel_24_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_13 XI11_5/XI0/XI0_24/d__13_ xsel_24_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_12 XI11_5/XI0/XI0_24/d__12_ xsel_24_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_11 XI11_5/XI0/XI0_24/d__11_ xsel_24_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_10 XI11_5/XI0/XI0_24/d__10_ xsel_24_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_9 XI11_5/XI0/XI0_24/d__9_ xsel_24_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_8 XI11_5/XI0/XI0_24/d__8_ xsel_24_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_7 XI11_5/XI0/XI0_24/d__7_ xsel_24_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_6 XI11_5/XI0/XI0_24/d__6_ xsel_24_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_5 XI11_5/XI0/XI0_24/d__5_ xsel_24_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_4 XI11_5/XI0/XI0_24/d__4_ xsel_24_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_3 XI11_5/XI0/XI0_24/d__3_ xsel_24_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_2 XI11_5/XI0/XI0_24/d__2_ xsel_24_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_1 XI11_5/XI0/XI0_24/d__1_ xsel_24_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_24/MN1_0 XI11_5/XI0/XI0_24/d__0_ xsel_24_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_15 XI11_5/net21_0_ xsel_23_ XI11_5/XI0/XI0_23/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_14 XI11_5/net21_1_ xsel_23_ XI11_5/XI0/XI0_23/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_13 XI11_5/net21_2_ xsel_23_ XI11_5/XI0/XI0_23/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_12 XI11_5/net21_3_ xsel_23_ XI11_5/XI0/XI0_23/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_11 XI11_5/net21_4_ xsel_23_ XI11_5/XI0/XI0_23/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_10 XI11_5/net21_5_ xsel_23_ XI11_5/XI0/XI0_23/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_9 XI11_5/net21_6_ xsel_23_ XI11_5/XI0/XI0_23/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_8 XI11_5/net21_7_ xsel_23_ XI11_5/XI0/XI0_23/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_7 XI11_5/net21_8_ xsel_23_ XI11_5/XI0/XI0_23/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_6 XI11_5/net21_9_ xsel_23_ XI11_5/XI0/XI0_23/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_5 XI11_5/net21_10_ xsel_23_ XI11_5/XI0/XI0_23/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_4 XI11_5/net21_11_ xsel_23_ XI11_5/XI0/XI0_23/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_3 XI11_5/net21_12_ xsel_23_ XI11_5/XI0/XI0_23/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_2 XI11_5/net21_13_ xsel_23_ XI11_5/XI0/XI0_23/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_1 XI11_5/net21_14_ xsel_23_ XI11_5/XI0/XI0_23/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN0_0 XI11_5/net21_15_ xsel_23_ XI11_5/XI0/XI0_23/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_15 XI11_5/XI0/XI0_23/d__15_ xsel_23_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_14 XI11_5/XI0/XI0_23/d__14_ xsel_23_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_13 XI11_5/XI0/XI0_23/d__13_ xsel_23_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_12 XI11_5/XI0/XI0_23/d__12_ xsel_23_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_11 XI11_5/XI0/XI0_23/d__11_ xsel_23_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_10 XI11_5/XI0/XI0_23/d__10_ xsel_23_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_9 XI11_5/XI0/XI0_23/d__9_ xsel_23_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_8 XI11_5/XI0/XI0_23/d__8_ xsel_23_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_7 XI11_5/XI0/XI0_23/d__7_ xsel_23_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_6 XI11_5/XI0/XI0_23/d__6_ xsel_23_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_5 XI11_5/XI0/XI0_23/d__5_ xsel_23_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_4 XI11_5/XI0/XI0_23/d__4_ xsel_23_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_3 XI11_5/XI0/XI0_23/d__3_ xsel_23_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_2 XI11_5/XI0/XI0_23/d__2_ xsel_23_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_1 XI11_5/XI0/XI0_23/d__1_ xsel_23_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_23/MN1_0 XI11_5/XI0/XI0_23/d__0_ xsel_23_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_15 XI11_5/net21_0_ xsel_22_ XI11_5/XI0/XI0_22/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_14 XI11_5/net21_1_ xsel_22_ XI11_5/XI0/XI0_22/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_13 XI11_5/net21_2_ xsel_22_ XI11_5/XI0/XI0_22/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_12 XI11_5/net21_3_ xsel_22_ XI11_5/XI0/XI0_22/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_11 XI11_5/net21_4_ xsel_22_ XI11_5/XI0/XI0_22/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_10 XI11_5/net21_5_ xsel_22_ XI11_5/XI0/XI0_22/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_9 XI11_5/net21_6_ xsel_22_ XI11_5/XI0/XI0_22/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_8 XI11_5/net21_7_ xsel_22_ XI11_5/XI0/XI0_22/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_7 XI11_5/net21_8_ xsel_22_ XI11_5/XI0/XI0_22/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_6 XI11_5/net21_9_ xsel_22_ XI11_5/XI0/XI0_22/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_5 XI11_5/net21_10_ xsel_22_ XI11_5/XI0/XI0_22/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_4 XI11_5/net21_11_ xsel_22_ XI11_5/XI0/XI0_22/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_3 XI11_5/net21_12_ xsel_22_ XI11_5/XI0/XI0_22/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_2 XI11_5/net21_13_ xsel_22_ XI11_5/XI0/XI0_22/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_1 XI11_5/net21_14_ xsel_22_ XI11_5/XI0/XI0_22/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN0_0 XI11_5/net21_15_ xsel_22_ XI11_5/XI0/XI0_22/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_15 XI11_5/XI0/XI0_22/d__15_ xsel_22_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_14 XI11_5/XI0/XI0_22/d__14_ xsel_22_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_13 XI11_5/XI0/XI0_22/d__13_ xsel_22_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_12 XI11_5/XI0/XI0_22/d__12_ xsel_22_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_11 XI11_5/XI0/XI0_22/d__11_ xsel_22_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_10 XI11_5/XI0/XI0_22/d__10_ xsel_22_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_9 XI11_5/XI0/XI0_22/d__9_ xsel_22_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_8 XI11_5/XI0/XI0_22/d__8_ xsel_22_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_7 XI11_5/XI0/XI0_22/d__7_ xsel_22_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_6 XI11_5/XI0/XI0_22/d__6_ xsel_22_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_5 XI11_5/XI0/XI0_22/d__5_ xsel_22_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_4 XI11_5/XI0/XI0_22/d__4_ xsel_22_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_3 XI11_5/XI0/XI0_22/d__3_ xsel_22_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_2 XI11_5/XI0/XI0_22/d__2_ xsel_22_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_1 XI11_5/XI0/XI0_22/d__1_ xsel_22_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_22/MN1_0 XI11_5/XI0/XI0_22/d__0_ xsel_22_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_15 XI11_5/net21_0_ xsel_21_ XI11_5/XI0/XI0_21/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_14 XI11_5/net21_1_ xsel_21_ XI11_5/XI0/XI0_21/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_13 XI11_5/net21_2_ xsel_21_ XI11_5/XI0/XI0_21/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_12 XI11_5/net21_3_ xsel_21_ XI11_5/XI0/XI0_21/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_11 XI11_5/net21_4_ xsel_21_ XI11_5/XI0/XI0_21/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_10 XI11_5/net21_5_ xsel_21_ XI11_5/XI0/XI0_21/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_9 XI11_5/net21_6_ xsel_21_ XI11_5/XI0/XI0_21/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_8 XI11_5/net21_7_ xsel_21_ XI11_5/XI0/XI0_21/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_7 XI11_5/net21_8_ xsel_21_ XI11_5/XI0/XI0_21/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_6 XI11_5/net21_9_ xsel_21_ XI11_5/XI0/XI0_21/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_5 XI11_5/net21_10_ xsel_21_ XI11_5/XI0/XI0_21/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_4 XI11_5/net21_11_ xsel_21_ XI11_5/XI0/XI0_21/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_3 XI11_5/net21_12_ xsel_21_ XI11_5/XI0/XI0_21/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_2 XI11_5/net21_13_ xsel_21_ XI11_5/XI0/XI0_21/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_1 XI11_5/net21_14_ xsel_21_ XI11_5/XI0/XI0_21/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN0_0 XI11_5/net21_15_ xsel_21_ XI11_5/XI0/XI0_21/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_15 XI11_5/XI0/XI0_21/d__15_ xsel_21_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_14 XI11_5/XI0/XI0_21/d__14_ xsel_21_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_13 XI11_5/XI0/XI0_21/d__13_ xsel_21_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_12 XI11_5/XI0/XI0_21/d__12_ xsel_21_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_11 XI11_5/XI0/XI0_21/d__11_ xsel_21_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_10 XI11_5/XI0/XI0_21/d__10_ xsel_21_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_9 XI11_5/XI0/XI0_21/d__9_ xsel_21_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_8 XI11_5/XI0/XI0_21/d__8_ xsel_21_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_7 XI11_5/XI0/XI0_21/d__7_ xsel_21_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_6 XI11_5/XI0/XI0_21/d__6_ xsel_21_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_5 XI11_5/XI0/XI0_21/d__5_ xsel_21_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_4 XI11_5/XI0/XI0_21/d__4_ xsel_21_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_3 XI11_5/XI0/XI0_21/d__3_ xsel_21_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_2 XI11_5/XI0/XI0_21/d__2_ xsel_21_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_1 XI11_5/XI0/XI0_21/d__1_ xsel_21_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_21/MN1_0 XI11_5/XI0/XI0_21/d__0_ xsel_21_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_15 XI11_5/net21_0_ xsel_20_ XI11_5/XI0/XI0_20/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_14 XI11_5/net21_1_ xsel_20_ XI11_5/XI0/XI0_20/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_13 XI11_5/net21_2_ xsel_20_ XI11_5/XI0/XI0_20/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_12 XI11_5/net21_3_ xsel_20_ XI11_5/XI0/XI0_20/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_11 XI11_5/net21_4_ xsel_20_ XI11_5/XI0/XI0_20/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_10 XI11_5/net21_5_ xsel_20_ XI11_5/XI0/XI0_20/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_9 XI11_5/net21_6_ xsel_20_ XI11_5/XI0/XI0_20/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_8 XI11_5/net21_7_ xsel_20_ XI11_5/XI0/XI0_20/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_7 XI11_5/net21_8_ xsel_20_ XI11_5/XI0/XI0_20/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_6 XI11_5/net21_9_ xsel_20_ XI11_5/XI0/XI0_20/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_5 XI11_5/net21_10_ xsel_20_ XI11_5/XI0/XI0_20/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_4 XI11_5/net21_11_ xsel_20_ XI11_5/XI0/XI0_20/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_3 XI11_5/net21_12_ xsel_20_ XI11_5/XI0/XI0_20/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_2 XI11_5/net21_13_ xsel_20_ XI11_5/XI0/XI0_20/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_1 XI11_5/net21_14_ xsel_20_ XI11_5/XI0/XI0_20/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN0_0 XI11_5/net21_15_ xsel_20_ XI11_5/XI0/XI0_20/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_15 XI11_5/XI0/XI0_20/d__15_ xsel_20_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_14 XI11_5/XI0/XI0_20/d__14_ xsel_20_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_13 XI11_5/XI0/XI0_20/d__13_ xsel_20_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_12 XI11_5/XI0/XI0_20/d__12_ xsel_20_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_11 XI11_5/XI0/XI0_20/d__11_ xsel_20_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_10 XI11_5/XI0/XI0_20/d__10_ xsel_20_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_9 XI11_5/XI0/XI0_20/d__9_ xsel_20_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_8 XI11_5/XI0/XI0_20/d__8_ xsel_20_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_7 XI11_5/XI0/XI0_20/d__7_ xsel_20_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_6 XI11_5/XI0/XI0_20/d__6_ xsel_20_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_5 XI11_5/XI0/XI0_20/d__5_ xsel_20_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_4 XI11_5/XI0/XI0_20/d__4_ xsel_20_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_3 XI11_5/XI0/XI0_20/d__3_ xsel_20_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_2 XI11_5/XI0/XI0_20/d__2_ xsel_20_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_1 XI11_5/XI0/XI0_20/d__1_ xsel_20_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_20/MN1_0 XI11_5/XI0/XI0_20/d__0_ xsel_20_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_15 XI11_5/net21_0_ xsel_19_ XI11_5/XI0/XI0_19/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_14 XI11_5/net21_1_ xsel_19_ XI11_5/XI0/XI0_19/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_13 XI11_5/net21_2_ xsel_19_ XI11_5/XI0/XI0_19/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_12 XI11_5/net21_3_ xsel_19_ XI11_5/XI0/XI0_19/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_11 XI11_5/net21_4_ xsel_19_ XI11_5/XI0/XI0_19/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_10 XI11_5/net21_5_ xsel_19_ XI11_5/XI0/XI0_19/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_9 XI11_5/net21_6_ xsel_19_ XI11_5/XI0/XI0_19/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_8 XI11_5/net21_7_ xsel_19_ XI11_5/XI0/XI0_19/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_7 XI11_5/net21_8_ xsel_19_ XI11_5/XI0/XI0_19/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_6 XI11_5/net21_9_ xsel_19_ XI11_5/XI0/XI0_19/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_5 XI11_5/net21_10_ xsel_19_ XI11_5/XI0/XI0_19/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_4 XI11_5/net21_11_ xsel_19_ XI11_5/XI0/XI0_19/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_3 XI11_5/net21_12_ xsel_19_ XI11_5/XI0/XI0_19/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_2 XI11_5/net21_13_ xsel_19_ XI11_5/XI0/XI0_19/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_1 XI11_5/net21_14_ xsel_19_ XI11_5/XI0/XI0_19/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN0_0 XI11_5/net21_15_ xsel_19_ XI11_5/XI0/XI0_19/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_15 XI11_5/XI0/XI0_19/d__15_ xsel_19_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_14 XI11_5/XI0/XI0_19/d__14_ xsel_19_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_13 XI11_5/XI0/XI0_19/d__13_ xsel_19_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_12 XI11_5/XI0/XI0_19/d__12_ xsel_19_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_11 XI11_5/XI0/XI0_19/d__11_ xsel_19_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_10 XI11_5/XI0/XI0_19/d__10_ xsel_19_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_9 XI11_5/XI0/XI0_19/d__9_ xsel_19_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_8 XI11_5/XI0/XI0_19/d__8_ xsel_19_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_7 XI11_5/XI0/XI0_19/d__7_ xsel_19_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_6 XI11_5/XI0/XI0_19/d__6_ xsel_19_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_5 XI11_5/XI0/XI0_19/d__5_ xsel_19_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_4 XI11_5/XI0/XI0_19/d__4_ xsel_19_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_3 XI11_5/XI0/XI0_19/d__3_ xsel_19_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_2 XI11_5/XI0/XI0_19/d__2_ xsel_19_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_1 XI11_5/XI0/XI0_19/d__1_ xsel_19_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_19/MN1_0 XI11_5/XI0/XI0_19/d__0_ xsel_19_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_15 XI11_5/net21_0_ xsel_18_ XI11_5/XI0/XI0_18/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_14 XI11_5/net21_1_ xsel_18_ XI11_5/XI0/XI0_18/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_13 XI11_5/net21_2_ xsel_18_ XI11_5/XI0/XI0_18/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_12 XI11_5/net21_3_ xsel_18_ XI11_5/XI0/XI0_18/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_11 XI11_5/net21_4_ xsel_18_ XI11_5/XI0/XI0_18/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_10 XI11_5/net21_5_ xsel_18_ XI11_5/XI0/XI0_18/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_9 XI11_5/net21_6_ xsel_18_ XI11_5/XI0/XI0_18/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_8 XI11_5/net21_7_ xsel_18_ XI11_5/XI0/XI0_18/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_7 XI11_5/net21_8_ xsel_18_ XI11_5/XI0/XI0_18/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_6 XI11_5/net21_9_ xsel_18_ XI11_5/XI0/XI0_18/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_5 XI11_5/net21_10_ xsel_18_ XI11_5/XI0/XI0_18/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_4 XI11_5/net21_11_ xsel_18_ XI11_5/XI0/XI0_18/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_3 XI11_5/net21_12_ xsel_18_ XI11_5/XI0/XI0_18/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_2 XI11_5/net21_13_ xsel_18_ XI11_5/XI0/XI0_18/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_1 XI11_5/net21_14_ xsel_18_ XI11_5/XI0/XI0_18/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN0_0 XI11_5/net21_15_ xsel_18_ XI11_5/XI0/XI0_18/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_15 XI11_5/XI0/XI0_18/d__15_ xsel_18_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_14 XI11_5/XI0/XI0_18/d__14_ xsel_18_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_13 XI11_5/XI0/XI0_18/d__13_ xsel_18_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_12 XI11_5/XI0/XI0_18/d__12_ xsel_18_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_11 XI11_5/XI0/XI0_18/d__11_ xsel_18_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_10 XI11_5/XI0/XI0_18/d__10_ xsel_18_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_9 XI11_5/XI0/XI0_18/d__9_ xsel_18_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_8 XI11_5/XI0/XI0_18/d__8_ xsel_18_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_7 XI11_5/XI0/XI0_18/d__7_ xsel_18_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_6 XI11_5/XI0/XI0_18/d__6_ xsel_18_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_5 XI11_5/XI0/XI0_18/d__5_ xsel_18_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_4 XI11_5/XI0/XI0_18/d__4_ xsel_18_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_3 XI11_5/XI0/XI0_18/d__3_ xsel_18_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_2 XI11_5/XI0/XI0_18/d__2_ xsel_18_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_1 XI11_5/XI0/XI0_18/d__1_ xsel_18_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_18/MN1_0 XI11_5/XI0/XI0_18/d__0_ xsel_18_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_15 XI11_5/net21_0_ xsel_17_ XI11_5/XI0/XI0_17/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_14 XI11_5/net21_1_ xsel_17_ XI11_5/XI0/XI0_17/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_13 XI11_5/net21_2_ xsel_17_ XI11_5/XI0/XI0_17/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_12 XI11_5/net21_3_ xsel_17_ XI11_5/XI0/XI0_17/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_11 XI11_5/net21_4_ xsel_17_ XI11_5/XI0/XI0_17/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_10 XI11_5/net21_5_ xsel_17_ XI11_5/XI0/XI0_17/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_9 XI11_5/net21_6_ xsel_17_ XI11_5/XI0/XI0_17/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_8 XI11_5/net21_7_ xsel_17_ XI11_5/XI0/XI0_17/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_7 XI11_5/net21_8_ xsel_17_ XI11_5/XI0/XI0_17/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_6 XI11_5/net21_9_ xsel_17_ XI11_5/XI0/XI0_17/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_5 XI11_5/net21_10_ xsel_17_ XI11_5/XI0/XI0_17/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_4 XI11_5/net21_11_ xsel_17_ XI11_5/XI0/XI0_17/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_3 XI11_5/net21_12_ xsel_17_ XI11_5/XI0/XI0_17/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_2 XI11_5/net21_13_ xsel_17_ XI11_5/XI0/XI0_17/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_1 XI11_5/net21_14_ xsel_17_ XI11_5/XI0/XI0_17/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN0_0 XI11_5/net21_15_ xsel_17_ XI11_5/XI0/XI0_17/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_15 XI11_5/XI0/XI0_17/d__15_ xsel_17_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_14 XI11_5/XI0/XI0_17/d__14_ xsel_17_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_13 XI11_5/XI0/XI0_17/d__13_ xsel_17_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_12 XI11_5/XI0/XI0_17/d__12_ xsel_17_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_11 XI11_5/XI0/XI0_17/d__11_ xsel_17_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_10 XI11_5/XI0/XI0_17/d__10_ xsel_17_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_9 XI11_5/XI0/XI0_17/d__9_ xsel_17_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_8 XI11_5/XI0/XI0_17/d__8_ xsel_17_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_7 XI11_5/XI0/XI0_17/d__7_ xsel_17_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_6 XI11_5/XI0/XI0_17/d__6_ xsel_17_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_5 XI11_5/XI0/XI0_17/d__5_ xsel_17_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_4 XI11_5/XI0/XI0_17/d__4_ xsel_17_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_3 XI11_5/XI0/XI0_17/d__3_ xsel_17_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_2 XI11_5/XI0/XI0_17/d__2_ xsel_17_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_1 XI11_5/XI0/XI0_17/d__1_ xsel_17_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_17/MN1_0 XI11_5/XI0/XI0_17/d__0_ xsel_17_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_15 XI11_5/net21_0_ xsel_16_ XI11_5/XI0/XI0_16/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_14 XI11_5/net21_1_ xsel_16_ XI11_5/XI0/XI0_16/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_13 XI11_5/net21_2_ xsel_16_ XI11_5/XI0/XI0_16/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_12 XI11_5/net21_3_ xsel_16_ XI11_5/XI0/XI0_16/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_11 XI11_5/net21_4_ xsel_16_ XI11_5/XI0/XI0_16/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_10 XI11_5/net21_5_ xsel_16_ XI11_5/XI0/XI0_16/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_9 XI11_5/net21_6_ xsel_16_ XI11_5/XI0/XI0_16/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_8 XI11_5/net21_7_ xsel_16_ XI11_5/XI0/XI0_16/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_7 XI11_5/net21_8_ xsel_16_ XI11_5/XI0/XI0_16/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_6 XI11_5/net21_9_ xsel_16_ XI11_5/XI0/XI0_16/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_5 XI11_5/net21_10_ xsel_16_ XI11_5/XI0/XI0_16/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_4 XI11_5/net21_11_ xsel_16_ XI11_5/XI0/XI0_16/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_3 XI11_5/net21_12_ xsel_16_ XI11_5/XI0/XI0_16/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_2 XI11_5/net21_13_ xsel_16_ XI11_5/XI0/XI0_16/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_1 XI11_5/net21_14_ xsel_16_ XI11_5/XI0/XI0_16/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN0_0 XI11_5/net21_15_ xsel_16_ XI11_5/XI0/XI0_16/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_15 XI11_5/XI0/XI0_16/d__15_ xsel_16_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_14 XI11_5/XI0/XI0_16/d__14_ xsel_16_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_13 XI11_5/XI0/XI0_16/d__13_ xsel_16_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_12 XI11_5/XI0/XI0_16/d__12_ xsel_16_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_11 XI11_5/XI0/XI0_16/d__11_ xsel_16_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_10 XI11_5/XI0/XI0_16/d__10_ xsel_16_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_9 XI11_5/XI0/XI0_16/d__9_ xsel_16_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_8 XI11_5/XI0/XI0_16/d__8_ xsel_16_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_7 XI11_5/XI0/XI0_16/d__7_ xsel_16_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_6 XI11_5/XI0/XI0_16/d__6_ xsel_16_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_5 XI11_5/XI0/XI0_16/d__5_ xsel_16_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_4 XI11_5/XI0/XI0_16/d__4_ xsel_16_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_3 XI11_5/XI0/XI0_16/d__3_ xsel_16_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_2 XI11_5/XI0/XI0_16/d__2_ xsel_16_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_1 XI11_5/XI0/XI0_16/d__1_ xsel_16_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_16/MN1_0 XI11_5/XI0/XI0_16/d__0_ xsel_16_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_15 XI11_5/net21_0_ xsel_15_ XI11_5/XI0/XI0_15/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_14 XI11_5/net21_1_ xsel_15_ XI11_5/XI0/XI0_15/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_13 XI11_5/net21_2_ xsel_15_ XI11_5/XI0/XI0_15/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_12 XI11_5/net21_3_ xsel_15_ XI11_5/XI0/XI0_15/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_11 XI11_5/net21_4_ xsel_15_ XI11_5/XI0/XI0_15/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_10 XI11_5/net21_5_ xsel_15_ XI11_5/XI0/XI0_15/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_9 XI11_5/net21_6_ xsel_15_ XI11_5/XI0/XI0_15/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_8 XI11_5/net21_7_ xsel_15_ XI11_5/XI0/XI0_15/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_7 XI11_5/net21_8_ xsel_15_ XI11_5/XI0/XI0_15/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_6 XI11_5/net21_9_ xsel_15_ XI11_5/XI0/XI0_15/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_5 XI11_5/net21_10_ xsel_15_ XI11_5/XI0/XI0_15/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_4 XI11_5/net21_11_ xsel_15_ XI11_5/XI0/XI0_15/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_3 XI11_5/net21_12_ xsel_15_ XI11_5/XI0/XI0_15/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_2 XI11_5/net21_13_ xsel_15_ XI11_5/XI0/XI0_15/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_1 XI11_5/net21_14_ xsel_15_ XI11_5/XI0/XI0_15/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN0_0 XI11_5/net21_15_ xsel_15_ XI11_5/XI0/XI0_15/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_15 XI11_5/XI0/XI0_15/d__15_ xsel_15_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_14 XI11_5/XI0/XI0_15/d__14_ xsel_15_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_13 XI11_5/XI0/XI0_15/d__13_ xsel_15_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_12 XI11_5/XI0/XI0_15/d__12_ xsel_15_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_11 XI11_5/XI0/XI0_15/d__11_ xsel_15_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_10 XI11_5/XI0/XI0_15/d__10_ xsel_15_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_9 XI11_5/XI0/XI0_15/d__9_ xsel_15_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_8 XI11_5/XI0/XI0_15/d__8_ xsel_15_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_7 XI11_5/XI0/XI0_15/d__7_ xsel_15_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_6 XI11_5/XI0/XI0_15/d__6_ xsel_15_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_5 XI11_5/XI0/XI0_15/d__5_ xsel_15_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_4 XI11_5/XI0/XI0_15/d__4_ xsel_15_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_3 XI11_5/XI0/XI0_15/d__3_ xsel_15_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_2 XI11_5/XI0/XI0_15/d__2_ xsel_15_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_1 XI11_5/XI0/XI0_15/d__1_ xsel_15_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_15/MN1_0 XI11_5/XI0/XI0_15/d__0_ xsel_15_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_15 XI11_5/net21_0_ xsel_14_ XI11_5/XI0/XI0_14/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_14 XI11_5/net21_1_ xsel_14_ XI11_5/XI0/XI0_14/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_13 XI11_5/net21_2_ xsel_14_ XI11_5/XI0/XI0_14/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_12 XI11_5/net21_3_ xsel_14_ XI11_5/XI0/XI0_14/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_11 XI11_5/net21_4_ xsel_14_ XI11_5/XI0/XI0_14/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_10 XI11_5/net21_5_ xsel_14_ XI11_5/XI0/XI0_14/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_9 XI11_5/net21_6_ xsel_14_ XI11_5/XI0/XI0_14/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_8 XI11_5/net21_7_ xsel_14_ XI11_5/XI0/XI0_14/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_7 XI11_5/net21_8_ xsel_14_ XI11_5/XI0/XI0_14/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_6 XI11_5/net21_9_ xsel_14_ XI11_5/XI0/XI0_14/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_5 XI11_5/net21_10_ xsel_14_ XI11_5/XI0/XI0_14/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_4 XI11_5/net21_11_ xsel_14_ XI11_5/XI0/XI0_14/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_3 XI11_5/net21_12_ xsel_14_ XI11_5/XI0/XI0_14/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_2 XI11_5/net21_13_ xsel_14_ XI11_5/XI0/XI0_14/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_1 XI11_5/net21_14_ xsel_14_ XI11_5/XI0/XI0_14/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN0_0 XI11_5/net21_15_ xsel_14_ XI11_5/XI0/XI0_14/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_15 XI11_5/XI0/XI0_14/d__15_ xsel_14_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_14 XI11_5/XI0/XI0_14/d__14_ xsel_14_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_13 XI11_5/XI0/XI0_14/d__13_ xsel_14_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_12 XI11_5/XI0/XI0_14/d__12_ xsel_14_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_11 XI11_5/XI0/XI0_14/d__11_ xsel_14_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_10 XI11_5/XI0/XI0_14/d__10_ xsel_14_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_9 XI11_5/XI0/XI0_14/d__9_ xsel_14_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_8 XI11_5/XI0/XI0_14/d__8_ xsel_14_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_7 XI11_5/XI0/XI0_14/d__7_ xsel_14_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_6 XI11_5/XI0/XI0_14/d__6_ xsel_14_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_5 XI11_5/XI0/XI0_14/d__5_ xsel_14_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_4 XI11_5/XI0/XI0_14/d__4_ xsel_14_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_3 XI11_5/XI0/XI0_14/d__3_ xsel_14_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_2 XI11_5/XI0/XI0_14/d__2_ xsel_14_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_1 XI11_5/XI0/XI0_14/d__1_ xsel_14_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_14/MN1_0 XI11_5/XI0/XI0_14/d__0_ xsel_14_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_15 XI11_5/net21_0_ xsel_13_ XI11_5/XI0/XI0_13/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_14 XI11_5/net21_1_ xsel_13_ XI11_5/XI0/XI0_13/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_13 XI11_5/net21_2_ xsel_13_ XI11_5/XI0/XI0_13/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_12 XI11_5/net21_3_ xsel_13_ XI11_5/XI0/XI0_13/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_11 XI11_5/net21_4_ xsel_13_ XI11_5/XI0/XI0_13/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_10 XI11_5/net21_5_ xsel_13_ XI11_5/XI0/XI0_13/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_9 XI11_5/net21_6_ xsel_13_ XI11_5/XI0/XI0_13/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_8 XI11_5/net21_7_ xsel_13_ XI11_5/XI0/XI0_13/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_7 XI11_5/net21_8_ xsel_13_ XI11_5/XI0/XI0_13/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_6 XI11_5/net21_9_ xsel_13_ XI11_5/XI0/XI0_13/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_5 XI11_5/net21_10_ xsel_13_ XI11_5/XI0/XI0_13/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_4 XI11_5/net21_11_ xsel_13_ XI11_5/XI0/XI0_13/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_3 XI11_5/net21_12_ xsel_13_ XI11_5/XI0/XI0_13/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_2 XI11_5/net21_13_ xsel_13_ XI11_5/XI0/XI0_13/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_1 XI11_5/net21_14_ xsel_13_ XI11_5/XI0/XI0_13/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN0_0 XI11_5/net21_15_ xsel_13_ XI11_5/XI0/XI0_13/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_15 XI11_5/XI0/XI0_13/d__15_ xsel_13_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_14 XI11_5/XI0/XI0_13/d__14_ xsel_13_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_13 XI11_5/XI0/XI0_13/d__13_ xsel_13_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_12 XI11_5/XI0/XI0_13/d__12_ xsel_13_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_11 XI11_5/XI0/XI0_13/d__11_ xsel_13_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_10 XI11_5/XI0/XI0_13/d__10_ xsel_13_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_9 XI11_5/XI0/XI0_13/d__9_ xsel_13_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_8 XI11_5/XI0/XI0_13/d__8_ xsel_13_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_7 XI11_5/XI0/XI0_13/d__7_ xsel_13_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_6 XI11_5/XI0/XI0_13/d__6_ xsel_13_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_5 XI11_5/XI0/XI0_13/d__5_ xsel_13_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_4 XI11_5/XI0/XI0_13/d__4_ xsel_13_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_3 XI11_5/XI0/XI0_13/d__3_ xsel_13_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_2 XI11_5/XI0/XI0_13/d__2_ xsel_13_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_1 XI11_5/XI0/XI0_13/d__1_ xsel_13_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_13/MN1_0 XI11_5/XI0/XI0_13/d__0_ xsel_13_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_15 XI11_5/net21_0_ xsel_12_ XI11_5/XI0/XI0_12/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_14 XI11_5/net21_1_ xsel_12_ XI11_5/XI0/XI0_12/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_13 XI11_5/net21_2_ xsel_12_ XI11_5/XI0/XI0_12/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_12 XI11_5/net21_3_ xsel_12_ XI11_5/XI0/XI0_12/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_11 XI11_5/net21_4_ xsel_12_ XI11_5/XI0/XI0_12/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_10 XI11_5/net21_5_ xsel_12_ XI11_5/XI0/XI0_12/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_9 XI11_5/net21_6_ xsel_12_ XI11_5/XI0/XI0_12/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_8 XI11_5/net21_7_ xsel_12_ XI11_5/XI0/XI0_12/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_7 XI11_5/net21_8_ xsel_12_ XI11_5/XI0/XI0_12/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_6 XI11_5/net21_9_ xsel_12_ XI11_5/XI0/XI0_12/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_5 XI11_5/net21_10_ xsel_12_ XI11_5/XI0/XI0_12/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_4 XI11_5/net21_11_ xsel_12_ XI11_5/XI0/XI0_12/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_3 XI11_5/net21_12_ xsel_12_ XI11_5/XI0/XI0_12/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_2 XI11_5/net21_13_ xsel_12_ XI11_5/XI0/XI0_12/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_1 XI11_5/net21_14_ xsel_12_ XI11_5/XI0/XI0_12/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN0_0 XI11_5/net21_15_ xsel_12_ XI11_5/XI0/XI0_12/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_15 XI11_5/XI0/XI0_12/d__15_ xsel_12_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_14 XI11_5/XI0/XI0_12/d__14_ xsel_12_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_13 XI11_5/XI0/XI0_12/d__13_ xsel_12_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_12 XI11_5/XI0/XI0_12/d__12_ xsel_12_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_11 XI11_5/XI0/XI0_12/d__11_ xsel_12_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_10 XI11_5/XI0/XI0_12/d__10_ xsel_12_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_9 XI11_5/XI0/XI0_12/d__9_ xsel_12_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_8 XI11_5/XI0/XI0_12/d__8_ xsel_12_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_7 XI11_5/XI0/XI0_12/d__7_ xsel_12_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_6 XI11_5/XI0/XI0_12/d__6_ xsel_12_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_5 XI11_5/XI0/XI0_12/d__5_ xsel_12_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_4 XI11_5/XI0/XI0_12/d__4_ xsel_12_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_3 XI11_5/XI0/XI0_12/d__3_ xsel_12_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_2 XI11_5/XI0/XI0_12/d__2_ xsel_12_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_1 XI11_5/XI0/XI0_12/d__1_ xsel_12_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_12/MN1_0 XI11_5/XI0/XI0_12/d__0_ xsel_12_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_15 XI11_5/net21_0_ xsel_11_ XI11_5/XI0/XI0_11/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_14 XI11_5/net21_1_ xsel_11_ XI11_5/XI0/XI0_11/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_13 XI11_5/net21_2_ xsel_11_ XI11_5/XI0/XI0_11/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_12 XI11_5/net21_3_ xsel_11_ XI11_5/XI0/XI0_11/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_11 XI11_5/net21_4_ xsel_11_ XI11_5/XI0/XI0_11/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_10 XI11_5/net21_5_ xsel_11_ XI11_5/XI0/XI0_11/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_9 XI11_5/net21_6_ xsel_11_ XI11_5/XI0/XI0_11/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_8 XI11_5/net21_7_ xsel_11_ XI11_5/XI0/XI0_11/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_7 XI11_5/net21_8_ xsel_11_ XI11_5/XI0/XI0_11/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_6 XI11_5/net21_9_ xsel_11_ XI11_5/XI0/XI0_11/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_5 XI11_5/net21_10_ xsel_11_ XI11_5/XI0/XI0_11/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_4 XI11_5/net21_11_ xsel_11_ XI11_5/XI0/XI0_11/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_3 XI11_5/net21_12_ xsel_11_ XI11_5/XI0/XI0_11/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_2 XI11_5/net21_13_ xsel_11_ XI11_5/XI0/XI0_11/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_1 XI11_5/net21_14_ xsel_11_ XI11_5/XI0/XI0_11/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN0_0 XI11_5/net21_15_ xsel_11_ XI11_5/XI0/XI0_11/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_15 XI11_5/XI0/XI0_11/d__15_ xsel_11_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_14 XI11_5/XI0/XI0_11/d__14_ xsel_11_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_13 XI11_5/XI0/XI0_11/d__13_ xsel_11_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_12 XI11_5/XI0/XI0_11/d__12_ xsel_11_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_11 XI11_5/XI0/XI0_11/d__11_ xsel_11_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_10 XI11_5/XI0/XI0_11/d__10_ xsel_11_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_9 XI11_5/XI0/XI0_11/d__9_ xsel_11_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_8 XI11_5/XI0/XI0_11/d__8_ xsel_11_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_7 XI11_5/XI0/XI0_11/d__7_ xsel_11_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_6 XI11_5/XI0/XI0_11/d__6_ xsel_11_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_5 XI11_5/XI0/XI0_11/d__5_ xsel_11_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_4 XI11_5/XI0/XI0_11/d__4_ xsel_11_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_3 XI11_5/XI0/XI0_11/d__3_ xsel_11_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_2 XI11_5/XI0/XI0_11/d__2_ xsel_11_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_1 XI11_5/XI0/XI0_11/d__1_ xsel_11_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_11/MN1_0 XI11_5/XI0/XI0_11/d__0_ xsel_11_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_15 XI11_5/net21_0_ xsel_10_ XI11_5/XI0/XI0_10/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_14 XI11_5/net21_1_ xsel_10_ XI11_5/XI0/XI0_10/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_13 XI11_5/net21_2_ xsel_10_ XI11_5/XI0/XI0_10/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_12 XI11_5/net21_3_ xsel_10_ XI11_5/XI0/XI0_10/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_11 XI11_5/net21_4_ xsel_10_ XI11_5/XI0/XI0_10/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_10 XI11_5/net21_5_ xsel_10_ XI11_5/XI0/XI0_10/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_9 XI11_5/net21_6_ xsel_10_ XI11_5/XI0/XI0_10/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_8 XI11_5/net21_7_ xsel_10_ XI11_5/XI0/XI0_10/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_7 XI11_5/net21_8_ xsel_10_ XI11_5/XI0/XI0_10/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_6 XI11_5/net21_9_ xsel_10_ XI11_5/XI0/XI0_10/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_5 XI11_5/net21_10_ xsel_10_ XI11_5/XI0/XI0_10/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_4 XI11_5/net21_11_ xsel_10_ XI11_5/XI0/XI0_10/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_3 XI11_5/net21_12_ xsel_10_ XI11_5/XI0/XI0_10/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_2 XI11_5/net21_13_ xsel_10_ XI11_5/XI0/XI0_10/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_1 XI11_5/net21_14_ xsel_10_ XI11_5/XI0/XI0_10/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN0_0 XI11_5/net21_15_ xsel_10_ XI11_5/XI0/XI0_10/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_15 XI11_5/XI0/XI0_10/d__15_ xsel_10_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_14 XI11_5/XI0/XI0_10/d__14_ xsel_10_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_13 XI11_5/XI0/XI0_10/d__13_ xsel_10_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_12 XI11_5/XI0/XI0_10/d__12_ xsel_10_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_11 XI11_5/XI0/XI0_10/d__11_ xsel_10_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_10 XI11_5/XI0/XI0_10/d__10_ xsel_10_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_9 XI11_5/XI0/XI0_10/d__9_ xsel_10_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_8 XI11_5/XI0/XI0_10/d__8_ xsel_10_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_7 XI11_5/XI0/XI0_10/d__7_ xsel_10_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_6 XI11_5/XI0/XI0_10/d__6_ xsel_10_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_5 XI11_5/XI0/XI0_10/d__5_ xsel_10_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_4 XI11_5/XI0/XI0_10/d__4_ xsel_10_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_3 XI11_5/XI0/XI0_10/d__3_ xsel_10_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_2 XI11_5/XI0/XI0_10/d__2_ xsel_10_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_1 XI11_5/XI0/XI0_10/d__1_ xsel_10_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_10/MN1_0 XI11_5/XI0/XI0_10/d__0_ xsel_10_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_15 XI11_5/net21_0_ xsel_9_ XI11_5/XI0/XI0_9/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_14 XI11_5/net21_1_ xsel_9_ XI11_5/XI0/XI0_9/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_13 XI11_5/net21_2_ xsel_9_ XI11_5/XI0/XI0_9/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_12 XI11_5/net21_3_ xsel_9_ XI11_5/XI0/XI0_9/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_11 XI11_5/net21_4_ xsel_9_ XI11_5/XI0/XI0_9/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_10 XI11_5/net21_5_ xsel_9_ XI11_5/XI0/XI0_9/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_9 XI11_5/net21_6_ xsel_9_ XI11_5/XI0/XI0_9/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_8 XI11_5/net21_7_ xsel_9_ XI11_5/XI0/XI0_9/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_7 XI11_5/net21_8_ xsel_9_ XI11_5/XI0/XI0_9/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_6 XI11_5/net21_9_ xsel_9_ XI11_5/XI0/XI0_9/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_5 XI11_5/net21_10_ xsel_9_ XI11_5/XI0/XI0_9/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_4 XI11_5/net21_11_ xsel_9_ XI11_5/XI0/XI0_9/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_3 XI11_5/net21_12_ xsel_9_ XI11_5/XI0/XI0_9/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_2 XI11_5/net21_13_ xsel_9_ XI11_5/XI0/XI0_9/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_1 XI11_5/net21_14_ xsel_9_ XI11_5/XI0/XI0_9/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN0_0 XI11_5/net21_15_ xsel_9_ XI11_5/XI0/XI0_9/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_15 XI11_5/XI0/XI0_9/d__15_ xsel_9_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_14 XI11_5/XI0/XI0_9/d__14_ xsel_9_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_13 XI11_5/XI0/XI0_9/d__13_ xsel_9_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_12 XI11_5/XI0/XI0_9/d__12_ xsel_9_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_11 XI11_5/XI0/XI0_9/d__11_ xsel_9_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_10 XI11_5/XI0/XI0_9/d__10_ xsel_9_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_9 XI11_5/XI0/XI0_9/d__9_ xsel_9_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_8 XI11_5/XI0/XI0_9/d__8_ xsel_9_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_7 XI11_5/XI0/XI0_9/d__7_ xsel_9_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_6 XI11_5/XI0/XI0_9/d__6_ xsel_9_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_5 XI11_5/XI0/XI0_9/d__5_ xsel_9_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_4 XI11_5/XI0/XI0_9/d__4_ xsel_9_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_3 XI11_5/XI0/XI0_9/d__3_ xsel_9_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_2 XI11_5/XI0/XI0_9/d__2_ xsel_9_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_1 XI11_5/XI0/XI0_9/d__1_ xsel_9_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_9/MN1_0 XI11_5/XI0/XI0_9/d__0_ xsel_9_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_15 XI11_5/net21_0_ xsel_8_ XI11_5/XI0/XI0_8/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_14 XI11_5/net21_1_ xsel_8_ XI11_5/XI0/XI0_8/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_13 XI11_5/net21_2_ xsel_8_ XI11_5/XI0/XI0_8/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_12 XI11_5/net21_3_ xsel_8_ XI11_5/XI0/XI0_8/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_11 XI11_5/net21_4_ xsel_8_ XI11_5/XI0/XI0_8/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_10 XI11_5/net21_5_ xsel_8_ XI11_5/XI0/XI0_8/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_9 XI11_5/net21_6_ xsel_8_ XI11_5/XI0/XI0_8/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_8 XI11_5/net21_7_ xsel_8_ XI11_5/XI0/XI0_8/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_7 XI11_5/net21_8_ xsel_8_ XI11_5/XI0/XI0_8/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_6 XI11_5/net21_9_ xsel_8_ XI11_5/XI0/XI0_8/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_5 XI11_5/net21_10_ xsel_8_ XI11_5/XI0/XI0_8/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_4 XI11_5/net21_11_ xsel_8_ XI11_5/XI0/XI0_8/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_3 XI11_5/net21_12_ xsel_8_ XI11_5/XI0/XI0_8/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_2 XI11_5/net21_13_ xsel_8_ XI11_5/XI0/XI0_8/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_1 XI11_5/net21_14_ xsel_8_ XI11_5/XI0/XI0_8/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN0_0 XI11_5/net21_15_ xsel_8_ XI11_5/XI0/XI0_8/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_15 XI11_5/XI0/XI0_8/d__15_ xsel_8_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_14 XI11_5/XI0/XI0_8/d__14_ xsel_8_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_13 XI11_5/XI0/XI0_8/d__13_ xsel_8_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_12 XI11_5/XI0/XI0_8/d__12_ xsel_8_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_11 XI11_5/XI0/XI0_8/d__11_ xsel_8_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_10 XI11_5/XI0/XI0_8/d__10_ xsel_8_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_9 XI11_5/XI0/XI0_8/d__9_ xsel_8_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_8 XI11_5/XI0/XI0_8/d__8_ xsel_8_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_7 XI11_5/XI0/XI0_8/d__7_ xsel_8_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_6 XI11_5/XI0/XI0_8/d__6_ xsel_8_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_5 XI11_5/XI0/XI0_8/d__5_ xsel_8_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_4 XI11_5/XI0/XI0_8/d__4_ xsel_8_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_3 XI11_5/XI0/XI0_8/d__3_ xsel_8_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_2 XI11_5/XI0/XI0_8/d__2_ xsel_8_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_1 XI11_5/XI0/XI0_8/d__1_ xsel_8_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_8/MN1_0 XI11_5/XI0/XI0_8/d__0_ xsel_8_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_15 XI11_5/net21_0_ xsel_7_ XI11_5/XI0/XI0_7/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_14 XI11_5/net21_1_ xsel_7_ XI11_5/XI0/XI0_7/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_13 XI11_5/net21_2_ xsel_7_ XI11_5/XI0/XI0_7/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_12 XI11_5/net21_3_ xsel_7_ XI11_5/XI0/XI0_7/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_11 XI11_5/net21_4_ xsel_7_ XI11_5/XI0/XI0_7/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_10 XI11_5/net21_5_ xsel_7_ XI11_5/XI0/XI0_7/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_9 XI11_5/net21_6_ xsel_7_ XI11_5/XI0/XI0_7/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_8 XI11_5/net21_7_ xsel_7_ XI11_5/XI0/XI0_7/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_7 XI11_5/net21_8_ xsel_7_ XI11_5/XI0/XI0_7/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_6 XI11_5/net21_9_ xsel_7_ XI11_5/XI0/XI0_7/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_5 XI11_5/net21_10_ xsel_7_ XI11_5/XI0/XI0_7/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_4 XI11_5/net21_11_ xsel_7_ XI11_5/XI0/XI0_7/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_3 XI11_5/net21_12_ xsel_7_ XI11_5/XI0/XI0_7/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_2 XI11_5/net21_13_ xsel_7_ XI11_5/XI0/XI0_7/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_1 XI11_5/net21_14_ xsel_7_ XI11_5/XI0/XI0_7/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN0_0 XI11_5/net21_15_ xsel_7_ XI11_5/XI0/XI0_7/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_15 XI11_5/XI0/XI0_7/d__15_ xsel_7_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_14 XI11_5/XI0/XI0_7/d__14_ xsel_7_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_13 XI11_5/XI0/XI0_7/d__13_ xsel_7_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_12 XI11_5/XI0/XI0_7/d__12_ xsel_7_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_11 XI11_5/XI0/XI0_7/d__11_ xsel_7_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_10 XI11_5/XI0/XI0_7/d__10_ xsel_7_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_9 XI11_5/XI0/XI0_7/d__9_ xsel_7_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_8 XI11_5/XI0/XI0_7/d__8_ xsel_7_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_7 XI11_5/XI0/XI0_7/d__7_ xsel_7_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_6 XI11_5/XI0/XI0_7/d__6_ xsel_7_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_5 XI11_5/XI0/XI0_7/d__5_ xsel_7_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_4 XI11_5/XI0/XI0_7/d__4_ xsel_7_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_3 XI11_5/XI0/XI0_7/d__3_ xsel_7_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_2 XI11_5/XI0/XI0_7/d__2_ xsel_7_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_1 XI11_5/XI0/XI0_7/d__1_ xsel_7_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_7/MN1_0 XI11_5/XI0/XI0_7/d__0_ xsel_7_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_15 XI11_5/net21_0_ xsel_6_ XI11_5/XI0/XI0_6/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_14 XI11_5/net21_1_ xsel_6_ XI11_5/XI0/XI0_6/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_13 XI11_5/net21_2_ xsel_6_ XI11_5/XI0/XI0_6/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_12 XI11_5/net21_3_ xsel_6_ XI11_5/XI0/XI0_6/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_11 XI11_5/net21_4_ xsel_6_ XI11_5/XI0/XI0_6/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_10 XI11_5/net21_5_ xsel_6_ XI11_5/XI0/XI0_6/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_9 XI11_5/net21_6_ xsel_6_ XI11_5/XI0/XI0_6/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_8 XI11_5/net21_7_ xsel_6_ XI11_5/XI0/XI0_6/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_7 XI11_5/net21_8_ xsel_6_ XI11_5/XI0/XI0_6/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_6 XI11_5/net21_9_ xsel_6_ XI11_5/XI0/XI0_6/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_5 XI11_5/net21_10_ xsel_6_ XI11_5/XI0/XI0_6/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_4 XI11_5/net21_11_ xsel_6_ XI11_5/XI0/XI0_6/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_3 XI11_5/net21_12_ xsel_6_ XI11_5/XI0/XI0_6/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_2 XI11_5/net21_13_ xsel_6_ XI11_5/XI0/XI0_6/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_1 XI11_5/net21_14_ xsel_6_ XI11_5/XI0/XI0_6/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN0_0 XI11_5/net21_15_ xsel_6_ XI11_5/XI0/XI0_6/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_15 XI11_5/XI0/XI0_6/d__15_ xsel_6_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_14 XI11_5/XI0/XI0_6/d__14_ xsel_6_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_13 XI11_5/XI0/XI0_6/d__13_ xsel_6_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_12 XI11_5/XI0/XI0_6/d__12_ xsel_6_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_11 XI11_5/XI0/XI0_6/d__11_ xsel_6_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_10 XI11_5/XI0/XI0_6/d__10_ xsel_6_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_9 XI11_5/XI0/XI0_6/d__9_ xsel_6_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_8 XI11_5/XI0/XI0_6/d__8_ xsel_6_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_7 XI11_5/XI0/XI0_6/d__7_ xsel_6_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_6 XI11_5/XI0/XI0_6/d__6_ xsel_6_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_5 XI11_5/XI0/XI0_6/d__5_ xsel_6_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_4 XI11_5/XI0/XI0_6/d__4_ xsel_6_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_3 XI11_5/XI0/XI0_6/d__3_ xsel_6_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_2 XI11_5/XI0/XI0_6/d__2_ xsel_6_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_1 XI11_5/XI0/XI0_6/d__1_ xsel_6_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_6/MN1_0 XI11_5/XI0/XI0_6/d__0_ xsel_6_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_15 XI11_5/net21_0_ xsel_5_ XI11_5/XI0/XI0_5/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_14 XI11_5/net21_1_ xsel_5_ XI11_5/XI0/XI0_5/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_13 XI11_5/net21_2_ xsel_5_ XI11_5/XI0/XI0_5/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_12 XI11_5/net21_3_ xsel_5_ XI11_5/XI0/XI0_5/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_11 XI11_5/net21_4_ xsel_5_ XI11_5/XI0/XI0_5/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_10 XI11_5/net21_5_ xsel_5_ XI11_5/XI0/XI0_5/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_9 XI11_5/net21_6_ xsel_5_ XI11_5/XI0/XI0_5/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_8 XI11_5/net21_7_ xsel_5_ XI11_5/XI0/XI0_5/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_7 XI11_5/net21_8_ xsel_5_ XI11_5/XI0/XI0_5/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_6 XI11_5/net21_9_ xsel_5_ XI11_5/XI0/XI0_5/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_5 XI11_5/net21_10_ xsel_5_ XI11_5/XI0/XI0_5/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_4 XI11_5/net21_11_ xsel_5_ XI11_5/XI0/XI0_5/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_3 XI11_5/net21_12_ xsel_5_ XI11_5/XI0/XI0_5/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_2 XI11_5/net21_13_ xsel_5_ XI11_5/XI0/XI0_5/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_1 XI11_5/net21_14_ xsel_5_ XI11_5/XI0/XI0_5/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN0_0 XI11_5/net21_15_ xsel_5_ XI11_5/XI0/XI0_5/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_15 XI11_5/XI0/XI0_5/d__15_ xsel_5_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_14 XI11_5/XI0/XI0_5/d__14_ xsel_5_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_13 XI11_5/XI0/XI0_5/d__13_ xsel_5_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_12 XI11_5/XI0/XI0_5/d__12_ xsel_5_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_11 XI11_5/XI0/XI0_5/d__11_ xsel_5_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_10 XI11_5/XI0/XI0_5/d__10_ xsel_5_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_9 XI11_5/XI0/XI0_5/d__9_ xsel_5_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_8 XI11_5/XI0/XI0_5/d__8_ xsel_5_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_7 XI11_5/XI0/XI0_5/d__7_ xsel_5_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_6 XI11_5/XI0/XI0_5/d__6_ xsel_5_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_5 XI11_5/XI0/XI0_5/d__5_ xsel_5_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_4 XI11_5/XI0/XI0_5/d__4_ xsel_5_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_3 XI11_5/XI0/XI0_5/d__3_ xsel_5_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_2 XI11_5/XI0/XI0_5/d__2_ xsel_5_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_1 XI11_5/XI0/XI0_5/d__1_ xsel_5_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_5/MN1_0 XI11_5/XI0/XI0_5/d__0_ xsel_5_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_15 XI11_5/net21_0_ xsel_4_ XI11_5/XI0/XI0_4/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_14 XI11_5/net21_1_ xsel_4_ XI11_5/XI0/XI0_4/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_13 XI11_5/net21_2_ xsel_4_ XI11_5/XI0/XI0_4/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_12 XI11_5/net21_3_ xsel_4_ XI11_5/XI0/XI0_4/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_11 XI11_5/net21_4_ xsel_4_ XI11_5/XI0/XI0_4/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_10 XI11_5/net21_5_ xsel_4_ XI11_5/XI0/XI0_4/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_9 XI11_5/net21_6_ xsel_4_ XI11_5/XI0/XI0_4/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_8 XI11_5/net21_7_ xsel_4_ XI11_5/XI0/XI0_4/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_7 XI11_5/net21_8_ xsel_4_ XI11_5/XI0/XI0_4/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_6 XI11_5/net21_9_ xsel_4_ XI11_5/XI0/XI0_4/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_5 XI11_5/net21_10_ xsel_4_ XI11_5/XI0/XI0_4/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_4 XI11_5/net21_11_ xsel_4_ XI11_5/XI0/XI0_4/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_3 XI11_5/net21_12_ xsel_4_ XI11_5/XI0/XI0_4/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_2 XI11_5/net21_13_ xsel_4_ XI11_5/XI0/XI0_4/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_1 XI11_5/net21_14_ xsel_4_ XI11_5/XI0/XI0_4/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN0_0 XI11_5/net21_15_ xsel_4_ XI11_5/XI0/XI0_4/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_15 XI11_5/XI0/XI0_4/d__15_ xsel_4_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_14 XI11_5/XI0/XI0_4/d__14_ xsel_4_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_13 XI11_5/XI0/XI0_4/d__13_ xsel_4_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_12 XI11_5/XI0/XI0_4/d__12_ xsel_4_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_11 XI11_5/XI0/XI0_4/d__11_ xsel_4_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_10 XI11_5/XI0/XI0_4/d__10_ xsel_4_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_9 XI11_5/XI0/XI0_4/d__9_ xsel_4_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_8 XI11_5/XI0/XI0_4/d__8_ xsel_4_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_7 XI11_5/XI0/XI0_4/d__7_ xsel_4_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_6 XI11_5/XI0/XI0_4/d__6_ xsel_4_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_5 XI11_5/XI0/XI0_4/d__5_ xsel_4_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_4 XI11_5/XI0/XI0_4/d__4_ xsel_4_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_3 XI11_5/XI0/XI0_4/d__3_ xsel_4_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_2 XI11_5/XI0/XI0_4/d__2_ xsel_4_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_1 XI11_5/XI0/XI0_4/d__1_ xsel_4_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_4/MN1_0 XI11_5/XI0/XI0_4/d__0_ xsel_4_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_15 XI11_5/net21_0_ xsel_3_ XI11_5/XI0/XI0_3/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_14 XI11_5/net21_1_ xsel_3_ XI11_5/XI0/XI0_3/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_13 XI11_5/net21_2_ xsel_3_ XI11_5/XI0/XI0_3/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_12 XI11_5/net21_3_ xsel_3_ XI11_5/XI0/XI0_3/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_11 XI11_5/net21_4_ xsel_3_ XI11_5/XI0/XI0_3/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_10 XI11_5/net21_5_ xsel_3_ XI11_5/XI0/XI0_3/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_9 XI11_5/net21_6_ xsel_3_ XI11_5/XI0/XI0_3/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_8 XI11_5/net21_7_ xsel_3_ XI11_5/XI0/XI0_3/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_7 XI11_5/net21_8_ xsel_3_ XI11_5/XI0/XI0_3/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_6 XI11_5/net21_9_ xsel_3_ XI11_5/XI0/XI0_3/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_5 XI11_5/net21_10_ xsel_3_ XI11_5/XI0/XI0_3/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_4 XI11_5/net21_11_ xsel_3_ XI11_5/XI0/XI0_3/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_3 XI11_5/net21_12_ xsel_3_ XI11_5/XI0/XI0_3/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_2 XI11_5/net21_13_ xsel_3_ XI11_5/XI0/XI0_3/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_1 XI11_5/net21_14_ xsel_3_ XI11_5/XI0/XI0_3/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN0_0 XI11_5/net21_15_ xsel_3_ XI11_5/XI0/XI0_3/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_15 XI11_5/XI0/XI0_3/d__15_ xsel_3_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_14 XI11_5/XI0/XI0_3/d__14_ xsel_3_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_13 XI11_5/XI0/XI0_3/d__13_ xsel_3_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_12 XI11_5/XI0/XI0_3/d__12_ xsel_3_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_11 XI11_5/XI0/XI0_3/d__11_ xsel_3_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_10 XI11_5/XI0/XI0_3/d__10_ xsel_3_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_9 XI11_5/XI0/XI0_3/d__9_ xsel_3_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_8 XI11_5/XI0/XI0_3/d__8_ xsel_3_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_7 XI11_5/XI0/XI0_3/d__7_ xsel_3_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_6 XI11_5/XI0/XI0_3/d__6_ xsel_3_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_5 XI11_5/XI0/XI0_3/d__5_ xsel_3_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_4 XI11_5/XI0/XI0_3/d__4_ xsel_3_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_3 XI11_5/XI0/XI0_3/d__3_ xsel_3_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_2 XI11_5/XI0/XI0_3/d__2_ xsel_3_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_1 XI11_5/XI0/XI0_3/d__1_ xsel_3_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_3/MN1_0 XI11_5/XI0/XI0_3/d__0_ xsel_3_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_15 XI11_5/net21_0_ xsel_2_ XI11_5/XI0/XI0_2/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_14 XI11_5/net21_1_ xsel_2_ XI11_5/XI0/XI0_2/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_13 XI11_5/net21_2_ xsel_2_ XI11_5/XI0/XI0_2/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_12 XI11_5/net21_3_ xsel_2_ XI11_5/XI0/XI0_2/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_11 XI11_5/net21_4_ xsel_2_ XI11_5/XI0/XI0_2/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_10 XI11_5/net21_5_ xsel_2_ XI11_5/XI0/XI0_2/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_9 XI11_5/net21_6_ xsel_2_ XI11_5/XI0/XI0_2/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_8 XI11_5/net21_7_ xsel_2_ XI11_5/XI0/XI0_2/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_7 XI11_5/net21_8_ xsel_2_ XI11_5/XI0/XI0_2/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_6 XI11_5/net21_9_ xsel_2_ XI11_5/XI0/XI0_2/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_5 XI11_5/net21_10_ xsel_2_ XI11_5/XI0/XI0_2/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_4 XI11_5/net21_11_ xsel_2_ XI11_5/XI0/XI0_2/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_3 XI11_5/net21_12_ xsel_2_ XI11_5/XI0/XI0_2/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_2 XI11_5/net21_13_ xsel_2_ XI11_5/XI0/XI0_2/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_1 XI11_5/net21_14_ xsel_2_ XI11_5/XI0/XI0_2/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN0_0 XI11_5/net21_15_ xsel_2_ XI11_5/XI0/XI0_2/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_15 XI11_5/XI0/XI0_2/d__15_ xsel_2_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_14 XI11_5/XI0/XI0_2/d__14_ xsel_2_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_13 XI11_5/XI0/XI0_2/d__13_ xsel_2_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_12 XI11_5/XI0/XI0_2/d__12_ xsel_2_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_11 XI11_5/XI0/XI0_2/d__11_ xsel_2_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_10 XI11_5/XI0/XI0_2/d__10_ xsel_2_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_9 XI11_5/XI0/XI0_2/d__9_ xsel_2_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_8 XI11_5/XI0/XI0_2/d__8_ xsel_2_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_7 XI11_5/XI0/XI0_2/d__7_ xsel_2_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_6 XI11_5/XI0/XI0_2/d__6_ xsel_2_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_5 XI11_5/XI0/XI0_2/d__5_ xsel_2_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_4 XI11_5/XI0/XI0_2/d__4_ xsel_2_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_3 XI11_5/XI0/XI0_2/d__3_ xsel_2_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_2 XI11_5/XI0/XI0_2/d__2_ xsel_2_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_1 XI11_5/XI0/XI0_2/d__1_ xsel_2_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_2/MN1_0 XI11_5/XI0/XI0_2/d__0_ xsel_2_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_15 XI11_5/net21_0_ xsel_1_ XI11_5/XI0/XI0_1/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_14 XI11_5/net21_1_ xsel_1_ XI11_5/XI0/XI0_1/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_13 XI11_5/net21_2_ xsel_1_ XI11_5/XI0/XI0_1/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_12 XI11_5/net21_3_ xsel_1_ XI11_5/XI0/XI0_1/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_11 XI11_5/net21_4_ xsel_1_ XI11_5/XI0/XI0_1/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_10 XI11_5/net21_5_ xsel_1_ XI11_5/XI0/XI0_1/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_9 XI11_5/net21_6_ xsel_1_ XI11_5/XI0/XI0_1/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_8 XI11_5/net21_7_ xsel_1_ XI11_5/XI0/XI0_1/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_7 XI11_5/net21_8_ xsel_1_ XI11_5/XI0/XI0_1/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_6 XI11_5/net21_9_ xsel_1_ XI11_5/XI0/XI0_1/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_5 XI11_5/net21_10_ xsel_1_ XI11_5/XI0/XI0_1/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_4 XI11_5/net21_11_ xsel_1_ XI11_5/XI0/XI0_1/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_3 XI11_5/net21_12_ xsel_1_ XI11_5/XI0/XI0_1/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_2 XI11_5/net21_13_ xsel_1_ XI11_5/XI0/XI0_1/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_1 XI11_5/net21_14_ xsel_1_ XI11_5/XI0/XI0_1/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN0_0 XI11_5/net21_15_ xsel_1_ XI11_5/XI0/XI0_1/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_15 XI11_5/XI0/XI0_1/d__15_ xsel_1_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_14 XI11_5/XI0/XI0_1/d__14_ xsel_1_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_13 XI11_5/XI0/XI0_1/d__13_ xsel_1_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_12 XI11_5/XI0/XI0_1/d__12_ xsel_1_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_11 XI11_5/XI0/XI0_1/d__11_ xsel_1_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_10 XI11_5/XI0/XI0_1/d__10_ xsel_1_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_9 XI11_5/XI0/XI0_1/d__9_ xsel_1_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_8 XI11_5/XI0/XI0_1/d__8_ xsel_1_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_7 XI11_5/XI0/XI0_1/d__7_ xsel_1_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_6 XI11_5/XI0/XI0_1/d__6_ xsel_1_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_5 XI11_5/XI0/XI0_1/d__5_ xsel_1_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_4 XI11_5/XI0/XI0_1/d__4_ xsel_1_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_3 XI11_5/XI0/XI0_1/d__3_ xsel_1_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_2 XI11_5/XI0/XI0_1/d__2_ xsel_1_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_1 XI11_5/XI0/XI0_1/d__1_ xsel_1_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_1/MN1_0 XI11_5/XI0/XI0_1/d__0_ xsel_1_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_15 XI11_5/net21_0_ xsel_0_ XI11_5/XI0/XI0_0/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_14 XI11_5/net21_1_ xsel_0_ XI11_5/XI0/XI0_0/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_13 XI11_5/net21_2_ xsel_0_ XI11_5/XI0/XI0_0/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_12 XI11_5/net21_3_ xsel_0_ XI11_5/XI0/XI0_0/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_11 XI11_5/net21_4_ xsel_0_ XI11_5/XI0/XI0_0/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_10 XI11_5/net21_5_ xsel_0_ XI11_5/XI0/XI0_0/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_9 XI11_5/net21_6_ xsel_0_ XI11_5/XI0/XI0_0/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_8 XI11_5/net21_7_ xsel_0_ XI11_5/XI0/XI0_0/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_7 XI11_5/net21_8_ xsel_0_ XI11_5/XI0/XI0_0/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_6 XI11_5/net21_9_ xsel_0_ XI11_5/XI0/XI0_0/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_5 XI11_5/net21_10_ xsel_0_ XI11_5/XI0/XI0_0/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_4 XI11_5/net21_11_ xsel_0_ XI11_5/XI0/XI0_0/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_3 XI11_5/net21_12_ xsel_0_ XI11_5/XI0/XI0_0/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_2 XI11_5/net21_13_ xsel_0_ XI11_5/XI0/XI0_0/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_1 XI11_5/net21_14_ xsel_0_ XI11_5/XI0/XI0_0/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN0_0 XI11_5/net21_15_ xsel_0_ XI11_5/XI0/XI0_0/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_15 XI11_5/XI0/XI0_0/d__15_ xsel_0_ XI11_5/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_14 XI11_5/XI0/XI0_0/d__14_ xsel_0_ XI11_5/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_13 XI11_5/XI0/XI0_0/d__13_ xsel_0_ XI11_5/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_12 XI11_5/XI0/XI0_0/d__12_ xsel_0_ XI11_5/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_11 XI11_5/XI0/XI0_0/d__11_ xsel_0_ XI11_5/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_10 XI11_5/XI0/XI0_0/d__10_ xsel_0_ XI11_5/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_9 XI11_5/XI0/XI0_0/d__9_ xsel_0_ XI11_5/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_8 XI11_5/XI0/XI0_0/d__8_ xsel_0_ XI11_5/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_7 XI11_5/XI0/XI0_0/d__7_ xsel_0_ XI11_5/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_6 XI11_5/XI0/XI0_0/d__6_ xsel_0_ XI11_5/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_5 XI11_5/XI0/XI0_0/d__5_ xsel_0_ XI11_5/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_4 XI11_5/XI0/XI0_0/d__4_ xsel_0_ XI11_5/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_3 XI11_5/XI0/XI0_0/d__3_ xsel_0_ XI11_5/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_2 XI11_5/XI0/XI0_0/d__2_ xsel_0_ XI11_5/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_1 XI11_5/XI0/XI0_0/d__1_ xsel_0_ XI11_5/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_5/XI0/XI0_0/MN1_0 XI11_5/XI0/XI0_0/d__0_ xsel_0_ XI11_5/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI2/MN0_15 XI11_4/net21_0_ ysel_15_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_14 XI11_4/net21_1_ ysel_14_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_13 XI11_4/net21_2_ ysel_13_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_12 XI11_4/net21_3_ ysel_12_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_11 XI11_4/net21_4_ ysel_11_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_10 XI11_4/net21_5_ ysel_10_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_9 XI11_4/net21_6_ ysel_9_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_8 XI11_4/net21_7_ ysel_8_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_7 XI11_4/net21_8_ ysel_7_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_6 XI11_4/net21_9_ ysel_6_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_5 XI11_4/net21_10_ ysel_5_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_4 XI11_4/net21_11_ ysel_4_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_3 XI11_4/net21_12_ ysel_3_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_2 XI11_4/net21_13_ ysel_2_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_1 XI11_4/net21_14_ ysel_1_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN0_0 XI11_4/net21_15_ ysel_0_ XI11_4/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_15 XI11_4/net20_0_ ysel_15_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_14 XI11_4/net20_1_ ysel_14_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_13 XI11_4/net20_2_ ysel_13_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_12 XI11_4/net20_3_ ysel_12_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_11 XI11_4/net20_4_ ysel_11_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_10 XI11_4/net20_5_ ysel_10_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_9 XI11_4/net20_6_ ysel_9_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_8 XI11_4/net20_7_ ysel_8_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_7 XI11_4/net20_8_ ysel_7_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_6 XI11_4/net20_9_ ysel_6_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_5 XI11_4/net20_10_ ysel_5_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_4 XI11_4/net20_11_ ysel_4_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_3 XI11_4/net20_12_ ysel_3_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_2 XI11_4/net20_13_ ysel_2_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_1 XI11_4/net20_14_ ysel_1_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI2/MN1_0 XI11_4/net20_15_ ysel_0_ XI11_4/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_4/XI4/MN8 vdd XI11_4/XI4/net8 XI11_4/net12 vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_4/XI4/MP0 XI11_4/net9 XI11_4/XI4/net23 vdd vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_4/XI4/MP4 XI11_4/net12 XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI4/MP1 XI11_4/net9 XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI4/MP5 XI11_4/net12 XI11_4/preck XI11_4/net9 vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI4/MN7 vdd XI11_4/XI4/net090 DOUT_4_ vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_4/XI4/MP3 gnd XI11_4/XI4/net089 XI11_4/net12 gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_4/XI4/MN5 XI11_4/net9 XI11_4/XI4/net0103 gnd gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_4/XI4/MN4 XI11_4/XI4/data_out_ XI11_4/XI4/net32 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_4/XI4/MN0 XI11_4/XI4/data_out XI11_4/XI4/net52 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_4/XI4/MN9 gnd XI11_4/XI4/net0112 DOUT_4_ gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_4/XI1_15/MP2 XI11_4/net20_0_ XI11_4/preck XI11_4/net21_0_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_15/MP1 XI11_4/net20_0_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_15/MP0 XI11_4/net21_0_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_14/MP2 XI11_4/net20_1_ XI11_4/preck XI11_4/net21_1_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_14/MP1 XI11_4/net20_1_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_14/MP0 XI11_4/net21_1_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_13/MP2 XI11_4/net20_2_ XI11_4/preck XI11_4/net21_2_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_13/MP1 XI11_4/net20_2_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_13/MP0 XI11_4/net21_2_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_12/MP2 XI11_4/net20_3_ XI11_4/preck XI11_4/net21_3_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_12/MP1 XI11_4/net20_3_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_12/MP0 XI11_4/net21_3_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_11/MP2 XI11_4/net20_4_ XI11_4/preck XI11_4/net21_4_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_11/MP1 XI11_4/net20_4_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_11/MP0 XI11_4/net21_4_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_10/MP2 XI11_4/net20_5_ XI11_4/preck XI11_4/net21_5_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_10/MP1 XI11_4/net20_5_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_10/MP0 XI11_4/net21_5_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_9/MP2 XI11_4/net20_6_ XI11_4/preck XI11_4/net21_6_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_9/MP1 XI11_4/net20_6_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_9/MP0 XI11_4/net21_6_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_8/MP2 XI11_4/net20_7_ XI11_4/preck XI11_4/net21_7_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_8/MP1 XI11_4/net20_7_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_8/MP0 XI11_4/net21_7_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_7/MP2 XI11_4/net20_8_ XI11_4/preck XI11_4/net21_8_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_7/MP1 XI11_4/net20_8_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_7/MP0 XI11_4/net21_8_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_6/MP2 XI11_4/net20_9_ XI11_4/preck XI11_4/net21_9_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_6/MP1 XI11_4/net20_9_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_6/MP0 XI11_4/net21_9_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_5/MP2 XI11_4/net20_10_ XI11_4/preck XI11_4/net21_10_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_5/MP1 XI11_4/net20_10_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_5/MP0 XI11_4/net21_10_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_4/MP2 XI11_4/net20_11_ XI11_4/preck XI11_4/net21_11_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_4/MP1 XI11_4/net20_11_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_4/MP0 XI11_4/net21_11_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_3/MP2 XI11_4/net20_12_ XI11_4/preck XI11_4/net21_12_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_3/MP1 XI11_4/net20_12_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_3/MP0 XI11_4/net21_12_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_2/MP2 XI11_4/net20_13_ XI11_4/preck XI11_4/net21_13_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_2/MP1 XI11_4/net20_13_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_2/MP0 XI11_4/net21_13_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_1/MP2 XI11_4/net20_14_ XI11_4/preck XI11_4/net21_14_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_1/MP1 XI11_4/net20_14_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_1/MP0 XI11_4/net21_14_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_0/MP2 XI11_4/net20_15_ XI11_4/preck XI11_4/net21_15_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_4/XI1_0/MP1 XI11_4/net20_15_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI1_0/MP0 XI11_4/net21_15_ XI11_4/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_4/XI0/MN0_15 gnd gnd XI11_4/net21_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_14 gnd gnd XI11_4/net21_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_13 gnd gnd XI11_4/net21_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_12 gnd gnd XI11_4/net21_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_11 gnd gnd XI11_4/net21_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_10 gnd gnd XI11_4/net21_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_9 gnd gnd XI11_4/net21_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_8 gnd gnd XI11_4/net21_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_7 gnd gnd XI11_4/net21_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_6 gnd gnd XI11_4/net21_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_5 gnd gnd XI11_4/net21_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_4 gnd gnd XI11_4/net21_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_3 gnd gnd XI11_4/net21_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_2 gnd gnd XI11_4/net21_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_1 gnd gnd XI11_4/net21_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN0_0 gnd gnd XI11_4/net21_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_15 gnd gnd XI11_4/net20_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_14 gnd gnd XI11_4/net20_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_13 gnd gnd XI11_4/net20_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_12 gnd gnd XI11_4/net20_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_11 gnd gnd XI11_4/net20_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_10 gnd gnd XI11_4/net20_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_9 gnd gnd XI11_4/net20_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_8 gnd gnd XI11_4/net20_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_7 gnd gnd XI11_4/net20_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_6 gnd gnd XI11_4/net20_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_5 gnd gnd XI11_4/net20_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_4 gnd gnd XI11_4/net20_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_3 gnd gnd XI11_4/net20_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_2 gnd gnd XI11_4/net20_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_1 gnd gnd XI11_4/net20_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/MN1_0 gnd gnd XI11_4/net20_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_15 XI11_4/net21_0_ xsel_63_ XI11_4/XI0/XI0_63/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_14 XI11_4/net21_1_ xsel_63_ XI11_4/XI0/XI0_63/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_13 XI11_4/net21_2_ xsel_63_ XI11_4/XI0/XI0_63/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_12 XI11_4/net21_3_ xsel_63_ XI11_4/XI0/XI0_63/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_11 XI11_4/net21_4_ xsel_63_ XI11_4/XI0/XI0_63/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_10 XI11_4/net21_5_ xsel_63_ XI11_4/XI0/XI0_63/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_9 XI11_4/net21_6_ xsel_63_ XI11_4/XI0/XI0_63/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_8 XI11_4/net21_7_ xsel_63_ XI11_4/XI0/XI0_63/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_7 XI11_4/net21_8_ xsel_63_ XI11_4/XI0/XI0_63/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_6 XI11_4/net21_9_ xsel_63_ XI11_4/XI0/XI0_63/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_5 XI11_4/net21_10_ xsel_63_ XI11_4/XI0/XI0_63/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_4 XI11_4/net21_11_ xsel_63_ XI11_4/XI0/XI0_63/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_3 XI11_4/net21_12_ xsel_63_ XI11_4/XI0/XI0_63/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_2 XI11_4/net21_13_ xsel_63_ XI11_4/XI0/XI0_63/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_1 XI11_4/net21_14_ xsel_63_ XI11_4/XI0/XI0_63/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN0_0 XI11_4/net21_15_ xsel_63_ XI11_4/XI0/XI0_63/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_15 XI11_4/XI0/XI0_63/d__15_ xsel_63_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_14 XI11_4/XI0/XI0_63/d__14_ xsel_63_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_13 XI11_4/XI0/XI0_63/d__13_ xsel_63_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_12 XI11_4/XI0/XI0_63/d__12_ xsel_63_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_11 XI11_4/XI0/XI0_63/d__11_ xsel_63_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_10 XI11_4/XI0/XI0_63/d__10_ xsel_63_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_9 XI11_4/XI0/XI0_63/d__9_ xsel_63_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_8 XI11_4/XI0/XI0_63/d__8_ xsel_63_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_7 XI11_4/XI0/XI0_63/d__7_ xsel_63_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_6 XI11_4/XI0/XI0_63/d__6_ xsel_63_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_5 XI11_4/XI0/XI0_63/d__5_ xsel_63_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_4 XI11_4/XI0/XI0_63/d__4_ xsel_63_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_3 XI11_4/XI0/XI0_63/d__3_ xsel_63_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_2 XI11_4/XI0/XI0_63/d__2_ xsel_63_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_1 XI11_4/XI0/XI0_63/d__1_ xsel_63_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_63/MN1_0 XI11_4/XI0/XI0_63/d__0_ xsel_63_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_15 XI11_4/net21_0_ xsel_62_ XI11_4/XI0/XI0_62/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_14 XI11_4/net21_1_ xsel_62_ XI11_4/XI0/XI0_62/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_13 XI11_4/net21_2_ xsel_62_ XI11_4/XI0/XI0_62/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_12 XI11_4/net21_3_ xsel_62_ XI11_4/XI0/XI0_62/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_11 XI11_4/net21_4_ xsel_62_ XI11_4/XI0/XI0_62/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_10 XI11_4/net21_5_ xsel_62_ XI11_4/XI0/XI0_62/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_9 XI11_4/net21_6_ xsel_62_ XI11_4/XI0/XI0_62/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_8 XI11_4/net21_7_ xsel_62_ XI11_4/XI0/XI0_62/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_7 XI11_4/net21_8_ xsel_62_ XI11_4/XI0/XI0_62/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_6 XI11_4/net21_9_ xsel_62_ XI11_4/XI0/XI0_62/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_5 XI11_4/net21_10_ xsel_62_ XI11_4/XI0/XI0_62/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_4 XI11_4/net21_11_ xsel_62_ XI11_4/XI0/XI0_62/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_3 XI11_4/net21_12_ xsel_62_ XI11_4/XI0/XI0_62/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_2 XI11_4/net21_13_ xsel_62_ XI11_4/XI0/XI0_62/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_1 XI11_4/net21_14_ xsel_62_ XI11_4/XI0/XI0_62/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN0_0 XI11_4/net21_15_ xsel_62_ XI11_4/XI0/XI0_62/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_15 XI11_4/XI0/XI0_62/d__15_ xsel_62_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_14 XI11_4/XI0/XI0_62/d__14_ xsel_62_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_13 XI11_4/XI0/XI0_62/d__13_ xsel_62_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_12 XI11_4/XI0/XI0_62/d__12_ xsel_62_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_11 XI11_4/XI0/XI0_62/d__11_ xsel_62_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_10 XI11_4/XI0/XI0_62/d__10_ xsel_62_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_9 XI11_4/XI0/XI0_62/d__9_ xsel_62_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_8 XI11_4/XI0/XI0_62/d__8_ xsel_62_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_7 XI11_4/XI0/XI0_62/d__7_ xsel_62_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_6 XI11_4/XI0/XI0_62/d__6_ xsel_62_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_5 XI11_4/XI0/XI0_62/d__5_ xsel_62_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_4 XI11_4/XI0/XI0_62/d__4_ xsel_62_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_3 XI11_4/XI0/XI0_62/d__3_ xsel_62_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_2 XI11_4/XI0/XI0_62/d__2_ xsel_62_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_1 XI11_4/XI0/XI0_62/d__1_ xsel_62_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_62/MN1_0 XI11_4/XI0/XI0_62/d__0_ xsel_62_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_15 XI11_4/net21_0_ xsel_61_ XI11_4/XI0/XI0_61/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_14 XI11_4/net21_1_ xsel_61_ XI11_4/XI0/XI0_61/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_13 XI11_4/net21_2_ xsel_61_ XI11_4/XI0/XI0_61/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_12 XI11_4/net21_3_ xsel_61_ XI11_4/XI0/XI0_61/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_11 XI11_4/net21_4_ xsel_61_ XI11_4/XI0/XI0_61/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_10 XI11_4/net21_5_ xsel_61_ XI11_4/XI0/XI0_61/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_9 XI11_4/net21_6_ xsel_61_ XI11_4/XI0/XI0_61/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_8 XI11_4/net21_7_ xsel_61_ XI11_4/XI0/XI0_61/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_7 XI11_4/net21_8_ xsel_61_ XI11_4/XI0/XI0_61/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_6 XI11_4/net21_9_ xsel_61_ XI11_4/XI0/XI0_61/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_5 XI11_4/net21_10_ xsel_61_ XI11_4/XI0/XI0_61/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_4 XI11_4/net21_11_ xsel_61_ XI11_4/XI0/XI0_61/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_3 XI11_4/net21_12_ xsel_61_ XI11_4/XI0/XI0_61/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_2 XI11_4/net21_13_ xsel_61_ XI11_4/XI0/XI0_61/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_1 XI11_4/net21_14_ xsel_61_ XI11_4/XI0/XI0_61/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN0_0 XI11_4/net21_15_ xsel_61_ XI11_4/XI0/XI0_61/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_15 XI11_4/XI0/XI0_61/d__15_ xsel_61_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_14 XI11_4/XI0/XI0_61/d__14_ xsel_61_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_13 XI11_4/XI0/XI0_61/d__13_ xsel_61_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_12 XI11_4/XI0/XI0_61/d__12_ xsel_61_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_11 XI11_4/XI0/XI0_61/d__11_ xsel_61_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_10 XI11_4/XI0/XI0_61/d__10_ xsel_61_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_9 XI11_4/XI0/XI0_61/d__9_ xsel_61_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_8 XI11_4/XI0/XI0_61/d__8_ xsel_61_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_7 XI11_4/XI0/XI0_61/d__7_ xsel_61_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_6 XI11_4/XI0/XI0_61/d__6_ xsel_61_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_5 XI11_4/XI0/XI0_61/d__5_ xsel_61_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_4 XI11_4/XI0/XI0_61/d__4_ xsel_61_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_3 XI11_4/XI0/XI0_61/d__3_ xsel_61_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_2 XI11_4/XI0/XI0_61/d__2_ xsel_61_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_1 XI11_4/XI0/XI0_61/d__1_ xsel_61_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_61/MN1_0 XI11_4/XI0/XI0_61/d__0_ xsel_61_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_15 XI11_4/net21_0_ xsel_60_ XI11_4/XI0/XI0_60/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_14 XI11_4/net21_1_ xsel_60_ XI11_4/XI0/XI0_60/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_13 XI11_4/net21_2_ xsel_60_ XI11_4/XI0/XI0_60/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_12 XI11_4/net21_3_ xsel_60_ XI11_4/XI0/XI0_60/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_11 XI11_4/net21_4_ xsel_60_ XI11_4/XI0/XI0_60/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_10 XI11_4/net21_5_ xsel_60_ XI11_4/XI0/XI0_60/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_9 XI11_4/net21_6_ xsel_60_ XI11_4/XI0/XI0_60/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_8 XI11_4/net21_7_ xsel_60_ XI11_4/XI0/XI0_60/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_7 XI11_4/net21_8_ xsel_60_ XI11_4/XI0/XI0_60/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_6 XI11_4/net21_9_ xsel_60_ XI11_4/XI0/XI0_60/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_5 XI11_4/net21_10_ xsel_60_ XI11_4/XI0/XI0_60/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_4 XI11_4/net21_11_ xsel_60_ XI11_4/XI0/XI0_60/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_3 XI11_4/net21_12_ xsel_60_ XI11_4/XI0/XI0_60/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_2 XI11_4/net21_13_ xsel_60_ XI11_4/XI0/XI0_60/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_1 XI11_4/net21_14_ xsel_60_ XI11_4/XI0/XI0_60/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN0_0 XI11_4/net21_15_ xsel_60_ XI11_4/XI0/XI0_60/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_15 XI11_4/XI0/XI0_60/d__15_ xsel_60_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_14 XI11_4/XI0/XI0_60/d__14_ xsel_60_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_13 XI11_4/XI0/XI0_60/d__13_ xsel_60_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_12 XI11_4/XI0/XI0_60/d__12_ xsel_60_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_11 XI11_4/XI0/XI0_60/d__11_ xsel_60_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_10 XI11_4/XI0/XI0_60/d__10_ xsel_60_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_9 XI11_4/XI0/XI0_60/d__9_ xsel_60_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_8 XI11_4/XI0/XI0_60/d__8_ xsel_60_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_7 XI11_4/XI0/XI0_60/d__7_ xsel_60_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_6 XI11_4/XI0/XI0_60/d__6_ xsel_60_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_5 XI11_4/XI0/XI0_60/d__5_ xsel_60_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_4 XI11_4/XI0/XI0_60/d__4_ xsel_60_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_3 XI11_4/XI0/XI0_60/d__3_ xsel_60_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_2 XI11_4/XI0/XI0_60/d__2_ xsel_60_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_1 XI11_4/XI0/XI0_60/d__1_ xsel_60_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_60/MN1_0 XI11_4/XI0/XI0_60/d__0_ xsel_60_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_15 XI11_4/net21_0_ xsel_59_ XI11_4/XI0/XI0_59/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_14 XI11_4/net21_1_ xsel_59_ XI11_4/XI0/XI0_59/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_13 XI11_4/net21_2_ xsel_59_ XI11_4/XI0/XI0_59/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_12 XI11_4/net21_3_ xsel_59_ XI11_4/XI0/XI0_59/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_11 XI11_4/net21_4_ xsel_59_ XI11_4/XI0/XI0_59/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_10 XI11_4/net21_5_ xsel_59_ XI11_4/XI0/XI0_59/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_9 XI11_4/net21_6_ xsel_59_ XI11_4/XI0/XI0_59/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_8 XI11_4/net21_7_ xsel_59_ XI11_4/XI0/XI0_59/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_7 XI11_4/net21_8_ xsel_59_ XI11_4/XI0/XI0_59/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_6 XI11_4/net21_9_ xsel_59_ XI11_4/XI0/XI0_59/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_5 XI11_4/net21_10_ xsel_59_ XI11_4/XI0/XI0_59/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_4 XI11_4/net21_11_ xsel_59_ XI11_4/XI0/XI0_59/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_3 XI11_4/net21_12_ xsel_59_ XI11_4/XI0/XI0_59/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_2 XI11_4/net21_13_ xsel_59_ XI11_4/XI0/XI0_59/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_1 XI11_4/net21_14_ xsel_59_ XI11_4/XI0/XI0_59/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN0_0 XI11_4/net21_15_ xsel_59_ XI11_4/XI0/XI0_59/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_15 XI11_4/XI0/XI0_59/d__15_ xsel_59_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_14 XI11_4/XI0/XI0_59/d__14_ xsel_59_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_13 XI11_4/XI0/XI0_59/d__13_ xsel_59_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_12 XI11_4/XI0/XI0_59/d__12_ xsel_59_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_11 XI11_4/XI0/XI0_59/d__11_ xsel_59_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_10 XI11_4/XI0/XI0_59/d__10_ xsel_59_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_9 XI11_4/XI0/XI0_59/d__9_ xsel_59_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_8 XI11_4/XI0/XI0_59/d__8_ xsel_59_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_7 XI11_4/XI0/XI0_59/d__7_ xsel_59_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_6 XI11_4/XI0/XI0_59/d__6_ xsel_59_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_5 XI11_4/XI0/XI0_59/d__5_ xsel_59_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_4 XI11_4/XI0/XI0_59/d__4_ xsel_59_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_3 XI11_4/XI0/XI0_59/d__3_ xsel_59_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_2 XI11_4/XI0/XI0_59/d__2_ xsel_59_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_1 XI11_4/XI0/XI0_59/d__1_ xsel_59_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_59/MN1_0 XI11_4/XI0/XI0_59/d__0_ xsel_59_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_15 XI11_4/net21_0_ xsel_58_ XI11_4/XI0/XI0_58/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_14 XI11_4/net21_1_ xsel_58_ XI11_4/XI0/XI0_58/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_13 XI11_4/net21_2_ xsel_58_ XI11_4/XI0/XI0_58/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_12 XI11_4/net21_3_ xsel_58_ XI11_4/XI0/XI0_58/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_11 XI11_4/net21_4_ xsel_58_ XI11_4/XI0/XI0_58/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_10 XI11_4/net21_5_ xsel_58_ XI11_4/XI0/XI0_58/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_9 XI11_4/net21_6_ xsel_58_ XI11_4/XI0/XI0_58/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_8 XI11_4/net21_7_ xsel_58_ XI11_4/XI0/XI0_58/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_7 XI11_4/net21_8_ xsel_58_ XI11_4/XI0/XI0_58/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_6 XI11_4/net21_9_ xsel_58_ XI11_4/XI0/XI0_58/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_5 XI11_4/net21_10_ xsel_58_ XI11_4/XI0/XI0_58/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_4 XI11_4/net21_11_ xsel_58_ XI11_4/XI0/XI0_58/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_3 XI11_4/net21_12_ xsel_58_ XI11_4/XI0/XI0_58/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_2 XI11_4/net21_13_ xsel_58_ XI11_4/XI0/XI0_58/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_1 XI11_4/net21_14_ xsel_58_ XI11_4/XI0/XI0_58/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN0_0 XI11_4/net21_15_ xsel_58_ XI11_4/XI0/XI0_58/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_15 XI11_4/XI0/XI0_58/d__15_ xsel_58_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_14 XI11_4/XI0/XI0_58/d__14_ xsel_58_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_13 XI11_4/XI0/XI0_58/d__13_ xsel_58_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_12 XI11_4/XI0/XI0_58/d__12_ xsel_58_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_11 XI11_4/XI0/XI0_58/d__11_ xsel_58_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_10 XI11_4/XI0/XI0_58/d__10_ xsel_58_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_9 XI11_4/XI0/XI0_58/d__9_ xsel_58_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_8 XI11_4/XI0/XI0_58/d__8_ xsel_58_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_7 XI11_4/XI0/XI0_58/d__7_ xsel_58_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_6 XI11_4/XI0/XI0_58/d__6_ xsel_58_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_5 XI11_4/XI0/XI0_58/d__5_ xsel_58_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_4 XI11_4/XI0/XI0_58/d__4_ xsel_58_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_3 XI11_4/XI0/XI0_58/d__3_ xsel_58_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_2 XI11_4/XI0/XI0_58/d__2_ xsel_58_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_1 XI11_4/XI0/XI0_58/d__1_ xsel_58_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_58/MN1_0 XI11_4/XI0/XI0_58/d__0_ xsel_58_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_15 XI11_4/net21_0_ xsel_57_ XI11_4/XI0/XI0_57/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_14 XI11_4/net21_1_ xsel_57_ XI11_4/XI0/XI0_57/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_13 XI11_4/net21_2_ xsel_57_ XI11_4/XI0/XI0_57/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_12 XI11_4/net21_3_ xsel_57_ XI11_4/XI0/XI0_57/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_11 XI11_4/net21_4_ xsel_57_ XI11_4/XI0/XI0_57/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_10 XI11_4/net21_5_ xsel_57_ XI11_4/XI0/XI0_57/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_9 XI11_4/net21_6_ xsel_57_ XI11_4/XI0/XI0_57/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_8 XI11_4/net21_7_ xsel_57_ XI11_4/XI0/XI0_57/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_7 XI11_4/net21_8_ xsel_57_ XI11_4/XI0/XI0_57/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_6 XI11_4/net21_9_ xsel_57_ XI11_4/XI0/XI0_57/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_5 XI11_4/net21_10_ xsel_57_ XI11_4/XI0/XI0_57/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_4 XI11_4/net21_11_ xsel_57_ XI11_4/XI0/XI0_57/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_3 XI11_4/net21_12_ xsel_57_ XI11_4/XI0/XI0_57/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_2 XI11_4/net21_13_ xsel_57_ XI11_4/XI0/XI0_57/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_1 XI11_4/net21_14_ xsel_57_ XI11_4/XI0/XI0_57/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN0_0 XI11_4/net21_15_ xsel_57_ XI11_4/XI0/XI0_57/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_15 XI11_4/XI0/XI0_57/d__15_ xsel_57_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_14 XI11_4/XI0/XI0_57/d__14_ xsel_57_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_13 XI11_4/XI0/XI0_57/d__13_ xsel_57_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_12 XI11_4/XI0/XI0_57/d__12_ xsel_57_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_11 XI11_4/XI0/XI0_57/d__11_ xsel_57_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_10 XI11_4/XI0/XI0_57/d__10_ xsel_57_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_9 XI11_4/XI0/XI0_57/d__9_ xsel_57_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_8 XI11_4/XI0/XI0_57/d__8_ xsel_57_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_7 XI11_4/XI0/XI0_57/d__7_ xsel_57_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_6 XI11_4/XI0/XI0_57/d__6_ xsel_57_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_5 XI11_4/XI0/XI0_57/d__5_ xsel_57_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_4 XI11_4/XI0/XI0_57/d__4_ xsel_57_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_3 XI11_4/XI0/XI0_57/d__3_ xsel_57_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_2 XI11_4/XI0/XI0_57/d__2_ xsel_57_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_1 XI11_4/XI0/XI0_57/d__1_ xsel_57_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_57/MN1_0 XI11_4/XI0/XI0_57/d__0_ xsel_57_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_15 XI11_4/net21_0_ xsel_56_ XI11_4/XI0/XI0_56/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_14 XI11_4/net21_1_ xsel_56_ XI11_4/XI0/XI0_56/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_13 XI11_4/net21_2_ xsel_56_ XI11_4/XI0/XI0_56/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_12 XI11_4/net21_3_ xsel_56_ XI11_4/XI0/XI0_56/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_11 XI11_4/net21_4_ xsel_56_ XI11_4/XI0/XI0_56/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_10 XI11_4/net21_5_ xsel_56_ XI11_4/XI0/XI0_56/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_9 XI11_4/net21_6_ xsel_56_ XI11_4/XI0/XI0_56/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_8 XI11_4/net21_7_ xsel_56_ XI11_4/XI0/XI0_56/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_7 XI11_4/net21_8_ xsel_56_ XI11_4/XI0/XI0_56/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_6 XI11_4/net21_9_ xsel_56_ XI11_4/XI0/XI0_56/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_5 XI11_4/net21_10_ xsel_56_ XI11_4/XI0/XI0_56/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_4 XI11_4/net21_11_ xsel_56_ XI11_4/XI0/XI0_56/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_3 XI11_4/net21_12_ xsel_56_ XI11_4/XI0/XI0_56/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_2 XI11_4/net21_13_ xsel_56_ XI11_4/XI0/XI0_56/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_1 XI11_4/net21_14_ xsel_56_ XI11_4/XI0/XI0_56/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN0_0 XI11_4/net21_15_ xsel_56_ XI11_4/XI0/XI0_56/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_15 XI11_4/XI0/XI0_56/d__15_ xsel_56_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_14 XI11_4/XI0/XI0_56/d__14_ xsel_56_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_13 XI11_4/XI0/XI0_56/d__13_ xsel_56_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_12 XI11_4/XI0/XI0_56/d__12_ xsel_56_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_11 XI11_4/XI0/XI0_56/d__11_ xsel_56_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_10 XI11_4/XI0/XI0_56/d__10_ xsel_56_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_9 XI11_4/XI0/XI0_56/d__9_ xsel_56_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_8 XI11_4/XI0/XI0_56/d__8_ xsel_56_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_7 XI11_4/XI0/XI0_56/d__7_ xsel_56_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_6 XI11_4/XI0/XI0_56/d__6_ xsel_56_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_5 XI11_4/XI0/XI0_56/d__5_ xsel_56_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_4 XI11_4/XI0/XI0_56/d__4_ xsel_56_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_3 XI11_4/XI0/XI0_56/d__3_ xsel_56_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_2 XI11_4/XI0/XI0_56/d__2_ xsel_56_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_1 XI11_4/XI0/XI0_56/d__1_ xsel_56_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_56/MN1_0 XI11_4/XI0/XI0_56/d__0_ xsel_56_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_15 XI11_4/net21_0_ xsel_55_ XI11_4/XI0/XI0_55/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_14 XI11_4/net21_1_ xsel_55_ XI11_4/XI0/XI0_55/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_13 XI11_4/net21_2_ xsel_55_ XI11_4/XI0/XI0_55/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_12 XI11_4/net21_3_ xsel_55_ XI11_4/XI0/XI0_55/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_11 XI11_4/net21_4_ xsel_55_ XI11_4/XI0/XI0_55/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_10 XI11_4/net21_5_ xsel_55_ XI11_4/XI0/XI0_55/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_9 XI11_4/net21_6_ xsel_55_ XI11_4/XI0/XI0_55/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_8 XI11_4/net21_7_ xsel_55_ XI11_4/XI0/XI0_55/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_7 XI11_4/net21_8_ xsel_55_ XI11_4/XI0/XI0_55/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_6 XI11_4/net21_9_ xsel_55_ XI11_4/XI0/XI0_55/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_5 XI11_4/net21_10_ xsel_55_ XI11_4/XI0/XI0_55/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_4 XI11_4/net21_11_ xsel_55_ XI11_4/XI0/XI0_55/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_3 XI11_4/net21_12_ xsel_55_ XI11_4/XI0/XI0_55/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_2 XI11_4/net21_13_ xsel_55_ XI11_4/XI0/XI0_55/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_1 XI11_4/net21_14_ xsel_55_ XI11_4/XI0/XI0_55/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN0_0 XI11_4/net21_15_ xsel_55_ XI11_4/XI0/XI0_55/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_15 XI11_4/XI0/XI0_55/d__15_ xsel_55_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_14 XI11_4/XI0/XI0_55/d__14_ xsel_55_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_13 XI11_4/XI0/XI0_55/d__13_ xsel_55_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_12 XI11_4/XI0/XI0_55/d__12_ xsel_55_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_11 XI11_4/XI0/XI0_55/d__11_ xsel_55_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_10 XI11_4/XI0/XI0_55/d__10_ xsel_55_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_9 XI11_4/XI0/XI0_55/d__9_ xsel_55_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_8 XI11_4/XI0/XI0_55/d__8_ xsel_55_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_7 XI11_4/XI0/XI0_55/d__7_ xsel_55_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_6 XI11_4/XI0/XI0_55/d__6_ xsel_55_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_5 XI11_4/XI0/XI0_55/d__5_ xsel_55_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_4 XI11_4/XI0/XI0_55/d__4_ xsel_55_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_3 XI11_4/XI0/XI0_55/d__3_ xsel_55_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_2 XI11_4/XI0/XI0_55/d__2_ xsel_55_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_1 XI11_4/XI0/XI0_55/d__1_ xsel_55_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_55/MN1_0 XI11_4/XI0/XI0_55/d__0_ xsel_55_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_15 XI11_4/net21_0_ xsel_54_ XI11_4/XI0/XI0_54/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_14 XI11_4/net21_1_ xsel_54_ XI11_4/XI0/XI0_54/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_13 XI11_4/net21_2_ xsel_54_ XI11_4/XI0/XI0_54/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_12 XI11_4/net21_3_ xsel_54_ XI11_4/XI0/XI0_54/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_11 XI11_4/net21_4_ xsel_54_ XI11_4/XI0/XI0_54/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_10 XI11_4/net21_5_ xsel_54_ XI11_4/XI0/XI0_54/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_9 XI11_4/net21_6_ xsel_54_ XI11_4/XI0/XI0_54/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_8 XI11_4/net21_7_ xsel_54_ XI11_4/XI0/XI0_54/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_7 XI11_4/net21_8_ xsel_54_ XI11_4/XI0/XI0_54/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_6 XI11_4/net21_9_ xsel_54_ XI11_4/XI0/XI0_54/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_5 XI11_4/net21_10_ xsel_54_ XI11_4/XI0/XI0_54/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_4 XI11_4/net21_11_ xsel_54_ XI11_4/XI0/XI0_54/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_3 XI11_4/net21_12_ xsel_54_ XI11_4/XI0/XI0_54/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_2 XI11_4/net21_13_ xsel_54_ XI11_4/XI0/XI0_54/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_1 XI11_4/net21_14_ xsel_54_ XI11_4/XI0/XI0_54/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN0_0 XI11_4/net21_15_ xsel_54_ XI11_4/XI0/XI0_54/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_15 XI11_4/XI0/XI0_54/d__15_ xsel_54_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_14 XI11_4/XI0/XI0_54/d__14_ xsel_54_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_13 XI11_4/XI0/XI0_54/d__13_ xsel_54_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_12 XI11_4/XI0/XI0_54/d__12_ xsel_54_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_11 XI11_4/XI0/XI0_54/d__11_ xsel_54_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_10 XI11_4/XI0/XI0_54/d__10_ xsel_54_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_9 XI11_4/XI0/XI0_54/d__9_ xsel_54_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_8 XI11_4/XI0/XI0_54/d__8_ xsel_54_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_7 XI11_4/XI0/XI0_54/d__7_ xsel_54_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_6 XI11_4/XI0/XI0_54/d__6_ xsel_54_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_5 XI11_4/XI0/XI0_54/d__5_ xsel_54_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_4 XI11_4/XI0/XI0_54/d__4_ xsel_54_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_3 XI11_4/XI0/XI0_54/d__3_ xsel_54_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_2 XI11_4/XI0/XI0_54/d__2_ xsel_54_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_1 XI11_4/XI0/XI0_54/d__1_ xsel_54_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_54/MN1_0 XI11_4/XI0/XI0_54/d__0_ xsel_54_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_15 XI11_4/net21_0_ xsel_53_ XI11_4/XI0/XI0_53/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_14 XI11_4/net21_1_ xsel_53_ XI11_4/XI0/XI0_53/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_13 XI11_4/net21_2_ xsel_53_ XI11_4/XI0/XI0_53/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_12 XI11_4/net21_3_ xsel_53_ XI11_4/XI0/XI0_53/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_11 XI11_4/net21_4_ xsel_53_ XI11_4/XI0/XI0_53/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_10 XI11_4/net21_5_ xsel_53_ XI11_4/XI0/XI0_53/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_9 XI11_4/net21_6_ xsel_53_ XI11_4/XI0/XI0_53/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_8 XI11_4/net21_7_ xsel_53_ XI11_4/XI0/XI0_53/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_7 XI11_4/net21_8_ xsel_53_ XI11_4/XI0/XI0_53/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_6 XI11_4/net21_9_ xsel_53_ XI11_4/XI0/XI0_53/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_5 XI11_4/net21_10_ xsel_53_ XI11_4/XI0/XI0_53/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_4 XI11_4/net21_11_ xsel_53_ XI11_4/XI0/XI0_53/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_3 XI11_4/net21_12_ xsel_53_ XI11_4/XI0/XI0_53/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_2 XI11_4/net21_13_ xsel_53_ XI11_4/XI0/XI0_53/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_1 XI11_4/net21_14_ xsel_53_ XI11_4/XI0/XI0_53/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN0_0 XI11_4/net21_15_ xsel_53_ XI11_4/XI0/XI0_53/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_15 XI11_4/XI0/XI0_53/d__15_ xsel_53_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_14 XI11_4/XI0/XI0_53/d__14_ xsel_53_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_13 XI11_4/XI0/XI0_53/d__13_ xsel_53_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_12 XI11_4/XI0/XI0_53/d__12_ xsel_53_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_11 XI11_4/XI0/XI0_53/d__11_ xsel_53_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_10 XI11_4/XI0/XI0_53/d__10_ xsel_53_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_9 XI11_4/XI0/XI0_53/d__9_ xsel_53_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_8 XI11_4/XI0/XI0_53/d__8_ xsel_53_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_7 XI11_4/XI0/XI0_53/d__7_ xsel_53_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_6 XI11_4/XI0/XI0_53/d__6_ xsel_53_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_5 XI11_4/XI0/XI0_53/d__5_ xsel_53_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_4 XI11_4/XI0/XI0_53/d__4_ xsel_53_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_3 XI11_4/XI0/XI0_53/d__3_ xsel_53_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_2 XI11_4/XI0/XI0_53/d__2_ xsel_53_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_1 XI11_4/XI0/XI0_53/d__1_ xsel_53_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_53/MN1_0 XI11_4/XI0/XI0_53/d__0_ xsel_53_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_15 XI11_4/net21_0_ xsel_52_ XI11_4/XI0/XI0_52/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_14 XI11_4/net21_1_ xsel_52_ XI11_4/XI0/XI0_52/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_13 XI11_4/net21_2_ xsel_52_ XI11_4/XI0/XI0_52/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_12 XI11_4/net21_3_ xsel_52_ XI11_4/XI0/XI0_52/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_11 XI11_4/net21_4_ xsel_52_ XI11_4/XI0/XI0_52/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_10 XI11_4/net21_5_ xsel_52_ XI11_4/XI0/XI0_52/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_9 XI11_4/net21_6_ xsel_52_ XI11_4/XI0/XI0_52/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_8 XI11_4/net21_7_ xsel_52_ XI11_4/XI0/XI0_52/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_7 XI11_4/net21_8_ xsel_52_ XI11_4/XI0/XI0_52/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_6 XI11_4/net21_9_ xsel_52_ XI11_4/XI0/XI0_52/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_5 XI11_4/net21_10_ xsel_52_ XI11_4/XI0/XI0_52/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_4 XI11_4/net21_11_ xsel_52_ XI11_4/XI0/XI0_52/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_3 XI11_4/net21_12_ xsel_52_ XI11_4/XI0/XI0_52/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_2 XI11_4/net21_13_ xsel_52_ XI11_4/XI0/XI0_52/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_1 XI11_4/net21_14_ xsel_52_ XI11_4/XI0/XI0_52/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN0_0 XI11_4/net21_15_ xsel_52_ XI11_4/XI0/XI0_52/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_15 XI11_4/XI0/XI0_52/d__15_ xsel_52_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_14 XI11_4/XI0/XI0_52/d__14_ xsel_52_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_13 XI11_4/XI0/XI0_52/d__13_ xsel_52_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_12 XI11_4/XI0/XI0_52/d__12_ xsel_52_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_11 XI11_4/XI0/XI0_52/d__11_ xsel_52_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_10 XI11_4/XI0/XI0_52/d__10_ xsel_52_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_9 XI11_4/XI0/XI0_52/d__9_ xsel_52_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_8 XI11_4/XI0/XI0_52/d__8_ xsel_52_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_7 XI11_4/XI0/XI0_52/d__7_ xsel_52_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_6 XI11_4/XI0/XI0_52/d__6_ xsel_52_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_5 XI11_4/XI0/XI0_52/d__5_ xsel_52_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_4 XI11_4/XI0/XI0_52/d__4_ xsel_52_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_3 XI11_4/XI0/XI0_52/d__3_ xsel_52_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_2 XI11_4/XI0/XI0_52/d__2_ xsel_52_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_1 XI11_4/XI0/XI0_52/d__1_ xsel_52_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_52/MN1_0 XI11_4/XI0/XI0_52/d__0_ xsel_52_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_15 XI11_4/net21_0_ xsel_51_ XI11_4/XI0/XI0_51/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_14 XI11_4/net21_1_ xsel_51_ XI11_4/XI0/XI0_51/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_13 XI11_4/net21_2_ xsel_51_ XI11_4/XI0/XI0_51/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_12 XI11_4/net21_3_ xsel_51_ XI11_4/XI0/XI0_51/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_11 XI11_4/net21_4_ xsel_51_ XI11_4/XI0/XI0_51/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_10 XI11_4/net21_5_ xsel_51_ XI11_4/XI0/XI0_51/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_9 XI11_4/net21_6_ xsel_51_ XI11_4/XI0/XI0_51/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_8 XI11_4/net21_7_ xsel_51_ XI11_4/XI0/XI0_51/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_7 XI11_4/net21_8_ xsel_51_ XI11_4/XI0/XI0_51/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_6 XI11_4/net21_9_ xsel_51_ XI11_4/XI0/XI0_51/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_5 XI11_4/net21_10_ xsel_51_ XI11_4/XI0/XI0_51/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_4 XI11_4/net21_11_ xsel_51_ XI11_4/XI0/XI0_51/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_3 XI11_4/net21_12_ xsel_51_ XI11_4/XI0/XI0_51/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_2 XI11_4/net21_13_ xsel_51_ XI11_4/XI0/XI0_51/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_1 XI11_4/net21_14_ xsel_51_ XI11_4/XI0/XI0_51/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN0_0 XI11_4/net21_15_ xsel_51_ XI11_4/XI0/XI0_51/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_15 XI11_4/XI0/XI0_51/d__15_ xsel_51_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_14 XI11_4/XI0/XI0_51/d__14_ xsel_51_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_13 XI11_4/XI0/XI0_51/d__13_ xsel_51_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_12 XI11_4/XI0/XI0_51/d__12_ xsel_51_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_11 XI11_4/XI0/XI0_51/d__11_ xsel_51_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_10 XI11_4/XI0/XI0_51/d__10_ xsel_51_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_9 XI11_4/XI0/XI0_51/d__9_ xsel_51_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_8 XI11_4/XI0/XI0_51/d__8_ xsel_51_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_7 XI11_4/XI0/XI0_51/d__7_ xsel_51_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_6 XI11_4/XI0/XI0_51/d__6_ xsel_51_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_5 XI11_4/XI0/XI0_51/d__5_ xsel_51_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_4 XI11_4/XI0/XI0_51/d__4_ xsel_51_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_3 XI11_4/XI0/XI0_51/d__3_ xsel_51_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_2 XI11_4/XI0/XI0_51/d__2_ xsel_51_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_1 XI11_4/XI0/XI0_51/d__1_ xsel_51_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_51/MN1_0 XI11_4/XI0/XI0_51/d__0_ xsel_51_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_15 XI11_4/net21_0_ xsel_50_ XI11_4/XI0/XI0_50/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_14 XI11_4/net21_1_ xsel_50_ XI11_4/XI0/XI0_50/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_13 XI11_4/net21_2_ xsel_50_ XI11_4/XI0/XI0_50/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_12 XI11_4/net21_3_ xsel_50_ XI11_4/XI0/XI0_50/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_11 XI11_4/net21_4_ xsel_50_ XI11_4/XI0/XI0_50/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_10 XI11_4/net21_5_ xsel_50_ XI11_4/XI0/XI0_50/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_9 XI11_4/net21_6_ xsel_50_ XI11_4/XI0/XI0_50/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_8 XI11_4/net21_7_ xsel_50_ XI11_4/XI0/XI0_50/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_7 XI11_4/net21_8_ xsel_50_ XI11_4/XI0/XI0_50/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_6 XI11_4/net21_9_ xsel_50_ XI11_4/XI0/XI0_50/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_5 XI11_4/net21_10_ xsel_50_ XI11_4/XI0/XI0_50/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_4 XI11_4/net21_11_ xsel_50_ XI11_4/XI0/XI0_50/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_3 XI11_4/net21_12_ xsel_50_ XI11_4/XI0/XI0_50/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_2 XI11_4/net21_13_ xsel_50_ XI11_4/XI0/XI0_50/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_1 XI11_4/net21_14_ xsel_50_ XI11_4/XI0/XI0_50/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN0_0 XI11_4/net21_15_ xsel_50_ XI11_4/XI0/XI0_50/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_15 XI11_4/XI0/XI0_50/d__15_ xsel_50_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_14 XI11_4/XI0/XI0_50/d__14_ xsel_50_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_13 XI11_4/XI0/XI0_50/d__13_ xsel_50_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_12 XI11_4/XI0/XI0_50/d__12_ xsel_50_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_11 XI11_4/XI0/XI0_50/d__11_ xsel_50_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_10 XI11_4/XI0/XI0_50/d__10_ xsel_50_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_9 XI11_4/XI0/XI0_50/d__9_ xsel_50_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_8 XI11_4/XI0/XI0_50/d__8_ xsel_50_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_7 XI11_4/XI0/XI0_50/d__7_ xsel_50_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_6 XI11_4/XI0/XI0_50/d__6_ xsel_50_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_5 XI11_4/XI0/XI0_50/d__5_ xsel_50_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_4 XI11_4/XI0/XI0_50/d__4_ xsel_50_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_3 XI11_4/XI0/XI0_50/d__3_ xsel_50_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_2 XI11_4/XI0/XI0_50/d__2_ xsel_50_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_1 XI11_4/XI0/XI0_50/d__1_ xsel_50_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_50/MN1_0 XI11_4/XI0/XI0_50/d__0_ xsel_50_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_15 XI11_4/net21_0_ xsel_49_ XI11_4/XI0/XI0_49/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_14 XI11_4/net21_1_ xsel_49_ XI11_4/XI0/XI0_49/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_13 XI11_4/net21_2_ xsel_49_ XI11_4/XI0/XI0_49/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_12 XI11_4/net21_3_ xsel_49_ XI11_4/XI0/XI0_49/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_11 XI11_4/net21_4_ xsel_49_ XI11_4/XI0/XI0_49/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_10 XI11_4/net21_5_ xsel_49_ XI11_4/XI0/XI0_49/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_9 XI11_4/net21_6_ xsel_49_ XI11_4/XI0/XI0_49/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_8 XI11_4/net21_7_ xsel_49_ XI11_4/XI0/XI0_49/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_7 XI11_4/net21_8_ xsel_49_ XI11_4/XI0/XI0_49/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_6 XI11_4/net21_9_ xsel_49_ XI11_4/XI0/XI0_49/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_5 XI11_4/net21_10_ xsel_49_ XI11_4/XI0/XI0_49/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_4 XI11_4/net21_11_ xsel_49_ XI11_4/XI0/XI0_49/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_3 XI11_4/net21_12_ xsel_49_ XI11_4/XI0/XI0_49/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_2 XI11_4/net21_13_ xsel_49_ XI11_4/XI0/XI0_49/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_1 XI11_4/net21_14_ xsel_49_ XI11_4/XI0/XI0_49/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN0_0 XI11_4/net21_15_ xsel_49_ XI11_4/XI0/XI0_49/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_15 XI11_4/XI0/XI0_49/d__15_ xsel_49_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_14 XI11_4/XI0/XI0_49/d__14_ xsel_49_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_13 XI11_4/XI0/XI0_49/d__13_ xsel_49_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_12 XI11_4/XI0/XI0_49/d__12_ xsel_49_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_11 XI11_4/XI0/XI0_49/d__11_ xsel_49_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_10 XI11_4/XI0/XI0_49/d__10_ xsel_49_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_9 XI11_4/XI0/XI0_49/d__9_ xsel_49_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_8 XI11_4/XI0/XI0_49/d__8_ xsel_49_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_7 XI11_4/XI0/XI0_49/d__7_ xsel_49_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_6 XI11_4/XI0/XI0_49/d__6_ xsel_49_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_5 XI11_4/XI0/XI0_49/d__5_ xsel_49_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_4 XI11_4/XI0/XI0_49/d__4_ xsel_49_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_3 XI11_4/XI0/XI0_49/d__3_ xsel_49_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_2 XI11_4/XI0/XI0_49/d__2_ xsel_49_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_1 XI11_4/XI0/XI0_49/d__1_ xsel_49_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_49/MN1_0 XI11_4/XI0/XI0_49/d__0_ xsel_49_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_15 XI11_4/net21_0_ xsel_48_ XI11_4/XI0/XI0_48/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_14 XI11_4/net21_1_ xsel_48_ XI11_4/XI0/XI0_48/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_13 XI11_4/net21_2_ xsel_48_ XI11_4/XI0/XI0_48/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_12 XI11_4/net21_3_ xsel_48_ XI11_4/XI0/XI0_48/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_11 XI11_4/net21_4_ xsel_48_ XI11_4/XI0/XI0_48/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_10 XI11_4/net21_5_ xsel_48_ XI11_4/XI0/XI0_48/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_9 XI11_4/net21_6_ xsel_48_ XI11_4/XI0/XI0_48/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_8 XI11_4/net21_7_ xsel_48_ XI11_4/XI0/XI0_48/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_7 XI11_4/net21_8_ xsel_48_ XI11_4/XI0/XI0_48/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_6 XI11_4/net21_9_ xsel_48_ XI11_4/XI0/XI0_48/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_5 XI11_4/net21_10_ xsel_48_ XI11_4/XI0/XI0_48/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_4 XI11_4/net21_11_ xsel_48_ XI11_4/XI0/XI0_48/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_3 XI11_4/net21_12_ xsel_48_ XI11_4/XI0/XI0_48/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_2 XI11_4/net21_13_ xsel_48_ XI11_4/XI0/XI0_48/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_1 XI11_4/net21_14_ xsel_48_ XI11_4/XI0/XI0_48/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN0_0 XI11_4/net21_15_ xsel_48_ XI11_4/XI0/XI0_48/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_15 XI11_4/XI0/XI0_48/d__15_ xsel_48_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_14 XI11_4/XI0/XI0_48/d__14_ xsel_48_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_13 XI11_4/XI0/XI0_48/d__13_ xsel_48_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_12 XI11_4/XI0/XI0_48/d__12_ xsel_48_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_11 XI11_4/XI0/XI0_48/d__11_ xsel_48_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_10 XI11_4/XI0/XI0_48/d__10_ xsel_48_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_9 XI11_4/XI0/XI0_48/d__9_ xsel_48_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_8 XI11_4/XI0/XI0_48/d__8_ xsel_48_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_7 XI11_4/XI0/XI0_48/d__7_ xsel_48_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_6 XI11_4/XI0/XI0_48/d__6_ xsel_48_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_5 XI11_4/XI0/XI0_48/d__5_ xsel_48_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_4 XI11_4/XI0/XI0_48/d__4_ xsel_48_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_3 XI11_4/XI0/XI0_48/d__3_ xsel_48_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_2 XI11_4/XI0/XI0_48/d__2_ xsel_48_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_1 XI11_4/XI0/XI0_48/d__1_ xsel_48_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_48/MN1_0 XI11_4/XI0/XI0_48/d__0_ xsel_48_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_15 XI11_4/net21_0_ xsel_47_ XI11_4/XI0/XI0_47/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_14 XI11_4/net21_1_ xsel_47_ XI11_4/XI0/XI0_47/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_13 XI11_4/net21_2_ xsel_47_ XI11_4/XI0/XI0_47/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_12 XI11_4/net21_3_ xsel_47_ XI11_4/XI0/XI0_47/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_11 XI11_4/net21_4_ xsel_47_ XI11_4/XI0/XI0_47/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_10 XI11_4/net21_5_ xsel_47_ XI11_4/XI0/XI0_47/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_9 XI11_4/net21_6_ xsel_47_ XI11_4/XI0/XI0_47/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_8 XI11_4/net21_7_ xsel_47_ XI11_4/XI0/XI0_47/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_7 XI11_4/net21_8_ xsel_47_ XI11_4/XI0/XI0_47/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_6 XI11_4/net21_9_ xsel_47_ XI11_4/XI0/XI0_47/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_5 XI11_4/net21_10_ xsel_47_ XI11_4/XI0/XI0_47/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_4 XI11_4/net21_11_ xsel_47_ XI11_4/XI0/XI0_47/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_3 XI11_4/net21_12_ xsel_47_ XI11_4/XI0/XI0_47/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_2 XI11_4/net21_13_ xsel_47_ XI11_4/XI0/XI0_47/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_1 XI11_4/net21_14_ xsel_47_ XI11_4/XI0/XI0_47/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN0_0 XI11_4/net21_15_ xsel_47_ XI11_4/XI0/XI0_47/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_15 XI11_4/XI0/XI0_47/d__15_ xsel_47_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_14 XI11_4/XI0/XI0_47/d__14_ xsel_47_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_13 XI11_4/XI0/XI0_47/d__13_ xsel_47_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_12 XI11_4/XI0/XI0_47/d__12_ xsel_47_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_11 XI11_4/XI0/XI0_47/d__11_ xsel_47_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_10 XI11_4/XI0/XI0_47/d__10_ xsel_47_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_9 XI11_4/XI0/XI0_47/d__9_ xsel_47_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_8 XI11_4/XI0/XI0_47/d__8_ xsel_47_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_7 XI11_4/XI0/XI0_47/d__7_ xsel_47_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_6 XI11_4/XI0/XI0_47/d__6_ xsel_47_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_5 XI11_4/XI0/XI0_47/d__5_ xsel_47_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_4 XI11_4/XI0/XI0_47/d__4_ xsel_47_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_3 XI11_4/XI0/XI0_47/d__3_ xsel_47_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_2 XI11_4/XI0/XI0_47/d__2_ xsel_47_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_1 XI11_4/XI0/XI0_47/d__1_ xsel_47_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_47/MN1_0 XI11_4/XI0/XI0_47/d__0_ xsel_47_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_15 XI11_4/net21_0_ xsel_46_ XI11_4/XI0/XI0_46/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_14 XI11_4/net21_1_ xsel_46_ XI11_4/XI0/XI0_46/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_13 XI11_4/net21_2_ xsel_46_ XI11_4/XI0/XI0_46/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_12 XI11_4/net21_3_ xsel_46_ XI11_4/XI0/XI0_46/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_11 XI11_4/net21_4_ xsel_46_ XI11_4/XI0/XI0_46/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_10 XI11_4/net21_5_ xsel_46_ XI11_4/XI0/XI0_46/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_9 XI11_4/net21_6_ xsel_46_ XI11_4/XI0/XI0_46/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_8 XI11_4/net21_7_ xsel_46_ XI11_4/XI0/XI0_46/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_7 XI11_4/net21_8_ xsel_46_ XI11_4/XI0/XI0_46/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_6 XI11_4/net21_9_ xsel_46_ XI11_4/XI0/XI0_46/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_5 XI11_4/net21_10_ xsel_46_ XI11_4/XI0/XI0_46/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_4 XI11_4/net21_11_ xsel_46_ XI11_4/XI0/XI0_46/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_3 XI11_4/net21_12_ xsel_46_ XI11_4/XI0/XI0_46/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_2 XI11_4/net21_13_ xsel_46_ XI11_4/XI0/XI0_46/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_1 XI11_4/net21_14_ xsel_46_ XI11_4/XI0/XI0_46/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN0_0 XI11_4/net21_15_ xsel_46_ XI11_4/XI0/XI0_46/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_15 XI11_4/XI0/XI0_46/d__15_ xsel_46_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_14 XI11_4/XI0/XI0_46/d__14_ xsel_46_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_13 XI11_4/XI0/XI0_46/d__13_ xsel_46_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_12 XI11_4/XI0/XI0_46/d__12_ xsel_46_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_11 XI11_4/XI0/XI0_46/d__11_ xsel_46_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_10 XI11_4/XI0/XI0_46/d__10_ xsel_46_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_9 XI11_4/XI0/XI0_46/d__9_ xsel_46_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_8 XI11_4/XI0/XI0_46/d__8_ xsel_46_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_7 XI11_4/XI0/XI0_46/d__7_ xsel_46_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_6 XI11_4/XI0/XI0_46/d__6_ xsel_46_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_5 XI11_4/XI0/XI0_46/d__5_ xsel_46_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_4 XI11_4/XI0/XI0_46/d__4_ xsel_46_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_3 XI11_4/XI0/XI0_46/d__3_ xsel_46_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_2 XI11_4/XI0/XI0_46/d__2_ xsel_46_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_1 XI11_4/XI0/XI0_46/d__1_ xsel_46_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_46/MN1_0 XI11_4/XI0/XI0_46/d__0_ xsel_46_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_15 XI11_4/net21_0_ xsel_45_ XI11_4/XI0/XI0_45/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_14 XI11_4/net21_1_ xsel_45_ XI11_4/XI0/XI0_45/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_13 XI11_4/net21_2_ xsel_45_ XI11_4/XI0/XI0_45/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_12 XI11_4/net21_3_ xsel_45_ XI11_4/XI0/XI0_45/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_11 XI11_4/net21_4_ xsel_45_ XI11_4/XI0/XI0_45/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_10 XI11_4/net21_5_ xsel_45_ XI11_4/XI0/XI0_45/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_9 XI11_4/net21_6_ xsel_45_ XI11_4/XI0/XI0_45/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_8 XI11_4/net21_7_ xsel_45_ XI11_4/XI0/XI0_45/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_7 XI11_4/net21_8_ xsel_45_ XI11_4/XI0/XI0_45/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_6 XI11_4/net21_9_ xsel_45_ XI11_4/XI0/XI0_45/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_5 XI11_4/net21_10_ xsel_45_ XI11_4/XI0/XI0_45/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_4 XI11_4/net21_11_ xsel_45_ XI11_4/XI0/XI0_45/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_3 XI11_4/net21_12_ xsel_45_ XI11_4/XI0/XI0_45/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_2 XI11_4/net21_13_ xsel_45_ XI11_4/XI0/XI0_45/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_1 XI11_4/net21_14_ xsel_45_ XI11_4/XI0/XI0_45/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN0_0 XI11_4/net21_15_ xsel_45_ XI11_4/XI0/XI0_45/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_15 XI11_4/XI0/XI0_45/d__15_ xsel_45_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_14 XI11_4/XI0/XI0_45/d__14_ xsel_45_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_13 XI11_4/XI0/XI0_45/d__13_ xsel_45_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_12 XI11_4/XI0/XI0_45/d__12_ xsel_45_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_11 XI11_4/XI0/XI0_45/d__11_ xsel_45_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_10 XI11_4/XI0/XI0_45/d__10_ xsel_45_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_9 XI11_4/XI0/XI0_45/d__9_ xsel_45_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_8 XI11_4/XI0/XI0_45/d__8_ xsel_45_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_7 XI11_4/XI0/XI0_45/d__7_ xsel_45_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_6 XI11_4/XI0/XI0_45/d__6_ xsel_45_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_5 XI11_4/XI0/XI0_45/d__5_ xsel_45_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_4 XI11_4/XI0/XI0_45/d__4_ xsel_45_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_3 XI11_4/XI0/XI0_45/d__3_ xsel_45_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_2 XI11_4/XI0/XI0_45/d__2_ xsel_45_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_1 XI11_4/XI0/XI0_45/d__1_ xsel_45_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_45/MN1_0 XI11_4/XI0/XI0_45/d__0_ xsel_45_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_15 XI11_4/net21_0_ xsel_44_ XI11_4/XI0/XI0_44/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_14 XI11_4/net21_1_ xsel_44_ XI11_4/XI0/XI0_44/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_13 XI11_4/net21_2_ xsel_44_ XI11_4/XI0/XI0_44/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_12 XI11_4/net21_3_ xsel_44_ XI11_4/XI0/XI0_44/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_11 XI11_4/net21_4_ xsel_44_ XI11_4/XI0/XI0_44/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_10 XI11_4/net21_5_ xsel_44_ XI11_4/XI0/XI0_44/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_9 XI11_4/net21_6_ xsel_44_ XI11_4/XI0/XI0_44/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_8 XI11_4/net21_7_ xsel_44_ XI11_4/XI0/XI0_44/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_7 XI11_4/net21_8_ xsel_44_ XI11_4/XI0/XI0_44/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_6 XI11_4/net21_9_ xsel_44_ XI11_4/XI0/XI0_44/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_5 XI11_4/net21_10_ xsel_44_ XI11_4/XI0/XI0_44/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_4 XI11_4/net21_11_ xsel_44_ XI11_4/XI0/XI0_44/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_3 XI11_4/net21_12_ xsel_44_ XI11_4/XI0/XI0_44/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_2 XI11_4/net21_13_ xsel_44_ XI11_4/XI0/XI0_44/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_1 XI11_4/net21_14_ xsel_44_ XI11_4/XI0/XI0_44/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN0_0 XI11_4/net21_15_ xsel_44_ XI11_4/XI0/XI0_44/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_15 XI11_4/XI0/XI0_44/d__15_ xsel_44_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_14 XI11_4/XI0/XI0_44/d__14_ xsel_44_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_13 XI11_4/XI0/XI0_44/d__13_ xsel_44_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_12 XI11_4/XI0/XI0_44/d__12_ xsel_44_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_11 XI11_4/XI0/XI0_44/d__11_ xsel_44_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_10 XI11_4/XI0/XI0_44/d__10_ xsel_44_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_9 XI11_4/XI0/XI0_44/d__9_ xsel_44_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_8 XI11_4/XI0/XI0_44/d__8_ xsel_44_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_7 XI11_4/XI0/XI0_44/d__7_ xsel_44_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_6 XI11_4/XI0/XI0_44/d__6_ xsel_44_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_5 XI11_4/XI0/XI0_44/d__5_ xsel_44_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_4 XI11_4/XI0/XI0_44/d__4_ xsel_44_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_3 XI11_4/XI0/XI0_44/d__3_ xsel_44_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_2 XI11_4/XI0/XI0_44/d__2_ xsel_44_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_1 XI11_4/XI0/XI0_44/d__1_ xsel_44_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_44/MN1_0 XI11_4/XI0/XI0_44/d__0_ xsel_44_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_15 XI11_4/net21_0_ xsel_43_ XI11_4/XI0/XI0_43/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_14 XI11_4/net21_1_ xsel_43_ XI11_4/XI0/XI0_43/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_13 XI11_4/net21_2_ xsel_43_ XI11_4/XI0/XI0_43/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_12 XI11_4/net21_3_ xsel_43_ XI11_4/XI0/XI0_43/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_11 XI11_4/net21_4_ xsel_43_ XI11_4/XI0/XI0_43/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_10 XI11_4/net21_5_ xsel_43_ XI11_4/XI0/XI0_43/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_9 XI11_4/net21_6_ xsel_43_ XI11_4/XI0/XI0_43/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_8 XI11_4/net21_7_ xsel_43_ XI11_4/XI0/XI0_43/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_7 XI11_4/net21_8_ xsel_43_ XI11_4/XI0/XI0_43/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_6 XI11_4/net21_9_ xsel_43_ XI11_4/XI0/XI0_43/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_5 XI11_4/net21_10_ xsel_43_ XI11_4/XI0/XI0_43/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_4 XI11_4/net21_11_ xsel_43_ XI11_4/XI0/XI0_43/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_3 XI11_4/net21_12_ xsel_43_ XI11_4/XI0/XI0_43/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_2 XI11_4/net21_13_ xsel_43_ XI11_4/XI0/XI0_43/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_1 XI11_4/net21_14_ xsel_43_ XI11_4/XI0/XI0_43/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN0_0 XI11_4/net21_15_ xsel_43_ XI11_4/XI0/XI0_43/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_15 XI11_4/XI0/XI0_43/d__15_ xsel_43_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_14 XI11_4/XI0/XI0_43/d__14_ xsel_43_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_13 XI11_4/XI0/XI0_43/d__13_ xsel_43_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_12 XI11_4/XI0/XI0_43/d__12_ xsel_43_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_11 XI11_4/XI0/XI0_43/d__11_ xsel_43_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_10 XI11_4/XI0/XI0_43/d__10_ xsel_43_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_9 XI11_4/XI0/XI0_43/d__9_ xsel_43_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_8 XI11_4/XI0/XI0_43/d__8_ xsel_43_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_7 XI11_4/XI0/XI0_43/d__7_ xsel_43_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_6 XI11_4/XI0/XI0_43/d__6_ xsel_43_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_5 XI11_4/XI0/XI0_43/d__5_ xsel_43_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_4 XI11_4/XI0/XI0_43/d__4_ xsel_43_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_3 XI11_4/XI0/XI0_43/d__3_ xsel_43_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_2 XI11_4/XI0/XI0_43/d__2_ xsel_43_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_1 XI11_4/XI0/XI0_43/d__1_ xsel_43_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_43/MN1_0 XI11_4/XI0/XI0_43/d__0_ xsel_43_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_15 XI11_4/net21_0_ xsel_42_ XI11_4/XI0/XI0_42/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_14 XI11_4/net21_1_ xsel_42_ XI11_4/XI0/XI0_42/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_13 XI11_4/net21_2_ xsel_42_ XI11_4/XI0/XI0_42/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_12 XI11_4/net21_3_ xsel_42_ XI11_4/XI0/XI0_42/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_11 XI11_4/net21_4_ xsel_42_ XI11_4/XI0/XI0_42/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_10 XI11_4/net21_5_ xsel_42_ XI11_4/XI0/XI0_42/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_9 XI11_4/net21_6_ xsel_42_ XI11_4/XI0/XI0_42/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_8 XI11_4/net21_7_ xsel_42_ XI11_4/XI0/XI0_42/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_7 XI11_4/net21_8_ xsel_42_ XI11_4/XI0/XI0_42/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_6 XI11_4/net21_9_ xsel_42_ XI11_4/XI0/XI0_42/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_5 XI11_4/net21_10_ xsel_42_ XI11_4/XI0/XI0_42/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_4 XI11_4/net21_11_ xsel_42_ XI11_4/XI0/XI0_42/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_3 XI11_4/net21_12_ xsel_42_ XI11_4/XI0/XI0_42/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_2 XI11_4/net21_13_ xsel_42_ XI11_4/XI0/XI0_42/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_1 XI11_4/net21_14_ xsel_42_ XI11_4/XI0/XI0_42/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN0_0 XI11_4/net21_15_ xsel_42_ XI11_4/XI0/XI0_42/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_15 XI11_4/XI0/XI0_42/d__15_ xsel_42_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_14 XI11_4/XI0/XI0_42/d__14_ xsel_42_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_13 XI11_4/XI0/XI0_42/d__13_ xsel_42_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_12 XI11_4/XI0/XI0_42/d__12_ xsel_42_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_11 XI11_4/XI0/XI0_42/d__11_ xsel_42_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_10 XI11_4/XI0/XI0_42/d__10_ xsel_42_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_9 XI11_4/XI0/XI0_42/d__9_ xsel_42_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_8 XI11_4/XI0/XI0_42/d__8_ xsel_42_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_7 XI11_4/XI0/XI0_42/d__7_ xsel_42_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_6 XI11_4/XI0/XI0_42/d__6_ xsel_42_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_5 XI11_4/XI0/XI0_42/d__5_ xsel_42_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_4 XI11_4/XI0/XI0_42/d__4_ xsel_42_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_3 XI11_4/XI0/XI0_42/d__3_ xsel_42_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_2 XI11_4/XI0/XI0_42/d__2_ xsel_42_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_1 XI11_4/XI0/XI0_42/d__1_ xsel_42_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_42/MN1_0 XI11_4/XI0/XI0_42/d__0_ xsel_42_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_15 XI11_4/net21_0_ xsel_41_ XI11_4/XI0/XI0_41/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_14 XI11_4/net21_1_ xsel_41_ XI11_4/XI0/XI0_41/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_13 XI11_4/net21_2_ xsel_41_ XI11_4/XI0/XI0_41/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_12 XI11_4/net21_3_ xsel_41_ XI11_4/XI0/XI0_41/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_11 XI11_4/net21_4_ xsel_41_ XI11_4/XI0/XI0_41/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_10 XI11_4/net21_5_ xsel_41_ XI11_4/XI0/XI0_41/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_9 XI11_4/net21_6_ xsel_41_ XI11_4/XI0/XI0_41/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_8 XI11_4/net21_7_ xsel_41_ XI11_4/XI0/XI0_41/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_7 XI11_4/net21_8_ xsel_41_ XI11_4/XI0/XI0_41/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_6 XI11_4/net21_9_ xsel_41_ XI11_4/XI0/XI0_41/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_5 XI11_4/net21_10_ xsel_41_ XI11_4/XI0/XI0_41/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_4 XI11_4/net21_11_ xsel_41_ XI11_4/XI0/XI0_41/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_3 XI11_4/net21_12_ xsel_41_ XI11_4/XI0/XI0_41/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_2 XI11_4/net21_13_ xsel_41_ XI11_4/XI0/XI0_41/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_1 XI11_4/net21_14_ xsel_41_ XI11_4/XI0/XI0_41/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN0_0 XI11_4/net21_15_ xsel_41_ XI11_4/XI0/XI0_41/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_15 XI11_4/XI0/XI0_41/d__15_ xsel_41_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_14 XI11_4/XI0/XI0_41/d__14_ xsel_41_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_13 XI11_4/XI0/XI0_41/d__13_ xsel_41_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_12 XI11_4/XI0/XI0_41/d__12_ xsel_41_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_11 XI11_4/XI0/XI0_41/d__11_ xsel_41_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_10 XI11_4/XI0/XI0_41/d__10_ xsel_41_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_9 XI11_4/XI0/XI0_41/d__9_ xsel_41_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_8 XI11_4/XI0/XI0_41/d__8_ xsel_41_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_7 XI11_4/XI0/XI0_41/d__7_ xsel_41_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_6 XI11_4/XI0/XI0_41/d__6_ xsel_41_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_5 XI11_4/XI0/XI0_41/d__5_ xsel_41_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_4 XI11_4/XI0/XI0_41/d__4_ xsel_41_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_3 XI11_4/XI0/XI0_41/d__3_ xsel_41_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_2 XI11_4/XI0/XI0_41/d__2_ xsel_41_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_1 XI11_4/XI0/XI0_41/d__1_ xsel_41_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_41/MN1_0 XI11_4/XI0/XI0_41/d__0_ xsel_41_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_15 XI11_4/net21_0_ xsel_40_ XI11_4/XI0/XI0_40/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_14 XI11_4/net21_1_ xsel_40_ XI11_4/XI0/XI0_40/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_13 XI11_4/net21_2_ xsel_40_ XI11_4/XI0/XI0_40/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_12 XI11_4/net21_3_ xsel_40_ XI11_4/XI0/XI0_40/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_11 XI11_4/net21_4_ xsel_40_ XI11_4/XI0/XI0_40/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_10 XI11_4/net21_5_ xsel_40_ XI11_4/XI0/XI0_40/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_9 XI11_4/net21_6_ xsel_40_ XI11_4/XI0/XI0_40/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_8 XI11_4/net21_7_ xsel_40_ XI11_4/XI0/XI0_40/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_7 XI11_4/net21_8_ xsel_40_ XI11_4/XI0/XI0_40/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_6 XI11_4/net21_9_ xsel_40_ XI11_4/XI0/XI0_40/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_5 XI11_4/net21_10_ xsel_40_ XI11_4/XI0/XI0_40/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_4 XI11_4/net21_11_ xsel_40_ XI11_4/XI0/XI0_40/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_3 XI11_4/net21_12_ xsel_40_ XI11_4/XI0/XI0_40/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_2 XI11_4/net21_13_ xsel_40_ XI11_4/XI0/XI0_40/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_1 XI11_4/net21_14_ xsel_40_ XI11_4/XI0/XI0_40/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN0_0 XI11_4/net21_15_ xsel_40_ XI11_4/XI0/XI0_40/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_15 XI11_4/XI0/XI0_40/d__15_ xsel_40_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_14 XI11_4/XI0/XI0_40/d__14_ xsel_40_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_13 XI11_4/XI0/XI0_40/d__13_ xsel_40_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_12 XI11_4/XI0/XI0_40/d__12_ xsel_40_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_11 XI11_4/XI0/XI0_40/d__11_ xsel_40_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_10 XI11_4/XI0/XI0_40/d__10_ xsel_40_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_9 XI11_4/XI0/XI0_40/d__9_ xsel_40_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_8 XI11_4/XI0/XI0_40/d__8_ xsel_40_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_7 XI11_4/XI0/XI0_40/d__7_ xsel_40_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_6 XI11_4/XI0/XI0_40/d__6_ xsel_40_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_5 XI11_4/XI0/XI0_40/d__5_ xsel_40_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_4 XI11_4/XI0/XI0_40/d__4_ xsel_40_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_3 XI11_4/XI0/XI0_40/d__3_ xsel_40_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_2 XI11_4/XI0/XI0_40/d__2_ xsel_40_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_1 XI11_4/XI0/XI0_40/d__1_ xsel_40_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_40/MN1_0 XI11_4/XI0/XI0_40/d__0_ xsel_40_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_15 XI11_4/net21_0_ xsel_39_ XI11_4/XI0/XI0_39/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_14 XI11_4/net21_1_ xsel_39_ XI11_4/XI0/XI0_39/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_13 XI11_4/net21_2_ xsel_39_ XI11_4/XI0/XI0_39/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_12 XI11_4/net21_3_ xsel_39_ XI11_4/XI0/XI0_39/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_11 XI11_4/net21_4_ xsel_39_ XI11_4/XI0/XI0_39/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_10 XI11_4/net21_5_ xsel_39_ XI11_4/XI0/XI0_39/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_9 XI11_4/net21_6_ xsel_39_ XI11_4/XI0/XI0_39/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_8 XI11_4/net21_7_ xsel_39_ XI11_4/XI0/XI0_39/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_7 XI11_4/net21_8_ xsel_39_ XI11_4/XI0/XI0_39/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_6 XI11_4/net21_9_ xsel_39_ XI11_4/XI0/XI0_39/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_5 XI11_4/net21_10_ xsel_39_ XI11_4/XI0/XI0_39/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_4 XI11_4/net21_11_ xsel_39_ XI11_4/XI0/XI0_39/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_3 XI11_4/net21_12_ xsel_39_ XI11_4/XI0/XI0_39/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_2 XI11_4/net21_13_ xsel_39_ XI11_4/XI0/XI0_39/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_1 XI11_4/net21_14_ xsel_39_ XI11_4/XI0/XI0_39/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN0_0 XI11_4/net21_15_ xsel_39_ XI11_4/XI0/XI0_39/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_15 XI11_4/XI0/XI0_39/d__15_ xsel_39_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_14 XI11_4/XI0/XI0_39/d__14_ xsel_39_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_13 XI11_4/XI0/XI0_39/d__13_ xsel_39_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_12 XI11_4/XI0/XI0_39/d__12_ xsel_39_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_11 XI11_4/XI0/XI0_39/d__11_ xsel_39_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_10 XI11_4/XI0/XI0_39/d__10_ xsel_39_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_9 XI11_4/XI0/XI0_39/d__9_ xsel_39_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_8 XI11_4/XI0/XI0_39/d__8_ xsel_39_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_7 XI11_4/XI0/XI0_39/d__7_ xsel_39_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_6 XI11_4/XI0/XI0_39/d__6_ xsel_39_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_5 XI11_4/XI0/XI0_39/d__5_ xsel_39_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_4 XI11_4/XI0/XI0_39/d__4_ xsel_39_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_3 XI11_4/XI0/XI0_39/d__3_ xsel_39_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_2 XI11_4/XI0/XI0_39/d__2_ xsel_39_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_1 XI11_4/XI0/XI0_39/d__1_ xsel_39_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_39/MN1_0 XI11_4/XI0/XI0_39/d__0_ xsel_39_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_15 XI11_4/net21_0_ xsel_38_ XI11_4/XI0/XI0_38/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_14 XI11_4/net21_1_ xsel_38_ XI11_4/XI0/XI0_38/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_13 XI11_4/net21_2_ xsel_38_ XI11_4/XI0/XI0_38/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_12 XI11_4/net21_3_ xsel_38_ XI11_4/XI0/XI0_38/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_11 XI11_4/net21_4_ xsel_38_ XI11_4/XI0/XI0_38/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_10 XI11_4/net21_5_ xsel_38_ XI11_4/XI0/XI0_38/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_9 XI11_4/net21_6_ xsel_38_ XI11_4/XI0/XI0_38/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_8 XI11_4/net21_7_ xsel_38_ XI11_4/XI0/XI0_38/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_7 XI11_4/net21_8_ xsel_38_ XI11_4/XI0/XI0_38/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_6 XI11_4/net21_9_ xsel_38_ XI11_4/XI0/XI0_38/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_5 XI11_4/net21_10_ xsel_38_ XI11_4/XI0/XI0_38/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_4 XI11_4/net21_11_ xsel_38_ XI11_4/XI0/XI0_38/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_3 XI11_4/net21_12_ xsel_38_ XI11_4/XI0/XI0_38/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_2 XI11_4/net21_13_ xsel_38_ XI11_4/XI0/XI0_38/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_1 XI11_4/net21_14_ xsel_38_ XI11_4/XI0/XI0_38/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN0_0 XI11_4/net21_15_ xsel_38_ XI11_4/XI0/XI0_38/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_15 XI11_4/XI0/XI0_38/d__15_ xsel_38_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_14 XI11_4/XI0/XI0_38/d__14_ xsel_38_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_13 XI11_4/XI0/XI0_38/d__13_ xsel_38_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_12 XI11_4/XI0/XI0_38/d__12_ xsel_38_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_11 XI11_4/XI0/XI0_38/d__11_ xsel_38_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_10 XI11_4/XI0/XI0_38/d__10_ xsel_38_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_9 XI11_4/XI0/XI0_38/d__9_ xsel_38_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_8 XI11_4/XI0/XI0_38/d__8_ xsel_38_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_7 XI11_4/XI0/XI0_38/d__7_ xsel_38_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_6 XI11_4/XI0/XI0_38/d__6_ xsel_38_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_5 XI11_4/XI0/XI0_38/d__5_ xsel_38_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_4 XI11_4/XI0/XI0_38/d__4_ xsel_38_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_3 XI11_4/XI0/XI0_38/d__3_ xsel_38_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_2 XI11_4/XI0/XI0_38/d__2_ xsel_38_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_1 XI11_4/XI0/XI0_38/d__1_ xsel_38_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_38/MN1_0 XI11_4/XI0/XI0_38/d__0_ xsel_38_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_15 XI11_4/net21_0_ xsel_37_ XI11_4/XI0/XI0_37/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_14 XI11_4/net21_1_ xsel_37_ XI11_4/XI0/XI0_37/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_13 XI11_4/net21_2_ xsel_37_ XI11_4/XI0/XI0_37/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_12 XI11_4/net21_3_ xsel_37_ XI11_4/XI0/XI0_37/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_11 XI11_4/net21_4_ xsel_37_ XI11_4/XI0/XI0_37/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_10 XI11_4/net21_5_ xsel_37_ XI11_4/XI0/XI0_37/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_9 XI11_4/net21_6_ xsel_37_ XI11_4/XI0/XI0_37/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_8 XI11_4/net21_7_ xsel_37_ XI11_4/XI0/XI0_37/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_7 XI11_4/net21_8_ xsel_37_ XI11_4/XI0/XI0_37/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_6 XI11_4/net21_9_ xsel_37_ XI11_4/XI0/XI0_37/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_5 XI11_4/net21_10_ xsel_37_ XI11_4/XI0/XI0_37/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_4 XI11_4/net21_11_ xsel_37_ XI11_4/XI0/XI0_37/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_3 XI11_4/net21_12_ xsel_37_ XI11_4/XI0/XI0_37/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_2 XI11_4/net21_13_ xsel_37_ XI11_4/XI0/XI0_37/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_1 XI11_4/net21_14_ xsel_37_ XI11_4/XI0/XI0_37/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN0_0 XI11_4/net21_15_ xsel_37_ XI11_4/XI0/XI0_37/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_15 XI11_4/XI0/XI0_37/d__15_ xsel_37_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_14 XI11_4/XI0/XI0_37/d__14_ xsel_37_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_13 XI11_4/XI0/XI0_37/d__13_ xsel_37_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_12 XI11_4/XI0/XI0_37/d__12_ xsel_37_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_11 XI11_4/XI0/XI0_37/d__11_ xsel_37_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_10 XI11_4/XI0/XI0_37/d__10_ xsel_37_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_9 XI11_4/XI0/XI0_37/d__9_ xsel_37_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_8 XI11_4/XI0/XI0_37/d__8_ xsel_37_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_7 XI11_4/XI0/XI0_37/d__7_ xsel_37_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_6 XI11_4/XI0/XI0_37/d__6_ xsel_37_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_5 XI11_4/XI0/XI0_37/d__5_ xsel_37_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_4 XI11_4/XI0/XI0_37/d__4_ xsel_37_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_3 XI11_4/XI0/XI0_37/d__3_ xsel_37_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_2 XI11_4/XI0/XI0_37/d__2_ xsel_37_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_1 XI11_4/XI0/XI0_37/d__1_ xsel_37_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_37/MN1_0 XI11_4/XI0/XI0_37/d__0_ xsel_37_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_15 XI11_4/net21_0_ xsel_36_ XI11_4/XI0/XI0_36/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_14 XI11_4/net21_1_ xsel_36_ XI11_4/XI0/XI0_36/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_13 XI11_4/net21_2_ xsel_36_ XI11_4/XI0/XI0_36/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_12 XI11_4/net21_3_ xsel_36_ XI11_4/XI0/XI0_36/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_11 XI11_4/net21_4_ xsel_36_ XI11_4/XI0/XI0_36/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_10 XI11_4/net21_5_ xsel_36_ XI11_4/XI0/XI0_36/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_9 XI11_4/net21_6_ xsel_36_ XI11_4/XI0/XI0_36/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_8 XI11_4/net21_7_ xsel_36_ XI11_4/XI0/XI0_36/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_7 XI11_4/net21_8_ xsel_36_ XI11_4/XI0/XI0_36/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_6 XI11_4/net21_9_ xsel_36_ XI11_4/XI0/XI0_36/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_5 XI11_4/net21_10_ xsel_36_ XI11_4/XI0/XI0_36/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_4 XI11_4/net21_11_ xsel_36_ XI11_4/XI0/XI0_36/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_3 XI11_4/net21_12_ xsel_36_ XI11_4/XI0/XI0_36/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_2 XI11_4/net21_13_ xsel_36_ XI11_4/XI0/XI0_36/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_1 XI11_4/net21_14_ xsel_36_ XI11_4/XI0/XI0_36/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN0_0 XI11_4/net21_15_ xsel_36_ XI11_4/XI0/XI0_36/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_15 XI11_4/XI0/XI0_36/d__15_ xsel_36_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_14 XI11_4/XI0/XI0_36/d__14_ xsel_36_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_13 XI11_4/XI0/XI0_36/d__13_ xsel_36_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_12 XI11_4/XI0/XI0_36/d__12_ xsel_36_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_11 XI11_4/XI0/XI0_36/d__11_ xsel_36_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_10 XI11_4/XI0/XI0_36/d__10_ xsel_36_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_9 XI11_4/XI0/XI0_36/d__9_ xsel_36_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_8 XI11_4/XI0/XI0_36/d__8_ xsel_36_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_7 XI11_4/XI0/XI0_36/d__7_ xsel_36_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_6 XI11_4/XI0/XI0_36/d__6_ xsel_36_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_5 XI11_4/XI0/XI0_36/d__5_ xsel_36_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_4 XI11_4/XI0/XI0_36/d__4_ xsel_36_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_3 XI11_4/XI0/XI0_36/d__3_ xsel_36_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_2 XI11_4/XI0/XI0_36/d__2_ xsel_36_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_1 XI11_4/XI0/XI0_36/d__1_ xsel_36_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_36/MN1_0 XI11_4/XI0/XI0_36/d__0_ xsel_36_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_15 XI11_4/net21_0_ xsel_35_ XI11_4/XI0/XI0_35/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_14 XI11_4/net21_1_ xsel_35_ XI11_4/XI0/XI0_35/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_13 XI11_4/net21_2_ xsel_35_ XI11_4/XI0/XI0_35/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_12 XI11_4/net21_3_ xsel_35_ XI11_4/XI0/XI0_35/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_11 XI11_4/net21_4_ xsel_35_ XI11_4/XI0/XI0_35/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_10 XI11_4/net21_5_ xsel_35_ XI11_4/XI0/XI0_35/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_9 XI11_4/net21_6_ xsel_35_ XI11_4/XI0/XI0_35/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_8 XI11_4/net21_7_ xsel_35_ XI11_4/XI0/XI0_35/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_7 XI11_4/net21_8_ xsel_35_ XI11_4/XI0/XI0_35/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_6 XI11_4/net21_9_ xsel_35_ XI11_4/XI0/XI0_35/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_5 XI11_4/net21_10_ xsel_35_ XI11_4/XI0/XI0_35/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_4 XI11_4/net21_11_ xsel_35_ XI11_4/XI0/XI0_35/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_3 XI11_4/net21_12_ xsel_35_ XI11_4/XI0/XI0_35/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_2 XI11_4/net21_13_ xsel_35_ XI11_4/XI0/XI0_35/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_1 XI11_4/net21_14_ xsel_35_ XI11_4/XI0/XI0_35/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN0_0 XI11_4/net21_15_ xsel_35_ XI11_4/XI0/XI0_35/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_15 XI11_4/XI0/XI0_35/d__15_ xsel_35_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_14 XI11_4/XI0/XI0_35/d__14_ xsel_35_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_13 XI11_4/XI0/XI0_35/d__13_ xsel_35_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_12 XI11_4/XI0/XI0_35/d__12_ xsel_35_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_11 XI11_4/XI0/XI0_35/d__11_ xsel_35_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_10 XI11_4/XI0/XI0_35/d__10_ xsel_35_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_9 XI11_4/XI0/XI0_35/d__9_ xsel_35_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_8 XI11_4/XI0/XI0_35/d__8_ xsel_35_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_7 XI11_4/XI0/XI0_35/d__7_ xsel_35_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_6 XI11_4/XI0/XI0_35/d__6_ xsel_35_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_5 XI11_4/XI0/XI0_35/d__5_ xsel_35_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_4 XI11_4/XI0/XI0_35/d__4_ xsel_35_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_3 XI11_4/XI0/XI0_35/d__3_ xsel_35_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_2 XI11_4/XI0/XI0_35/d__2_ xsel_35_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_1 XI11_4/XI0/XI0_35/d__1_ xsel_35_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_35/MN1_0 XI11_4/XI0/XI0_35/d__0_ xsel_35_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_15 XI11_4/net21_0_ xsel_34_ XI11_4/XI0/XI0_34/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_14 XI11_4/net21_1_ xsel_34_ XI11_4/XI0/XI0_34/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_13 XI11_4/net21_2_ xsel_34_ XI11_4/XI0/XI0_34/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_12 XI11_4/net21_3_ xsel_34_ XI11_4/XI0/XI0_34/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_11 XI11_4/net21_4_ xsel_34_ XI11_4/XI0/XI0_34/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_10 XI11_4/net21_5_ xsel_34_ XI11_4/XI0/XI0_34/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_9 XI11_4/net21_6_ xsel_34_ XI11_4/XI0/XI0_34/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_8 XI11_4/net21_7_ xsel_34_ XI11_4/XI0/XI0_34/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_7 XI11_4/net21_8_ xsel_34_ XI11_4/XI0/XI0_34/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_6 XI11_4/net21_9_ xsel_34_ XI11_4/XI0/XI0_34/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_5 XI11_4/net21_10_ xsel_34_ XI11_4/XI0/XI0_34/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_4 XI11_4/net21_11_ xsel_34_ XI11_4/XI0/XI0_34/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_3 XI11_4/net21_12_ xsel_34_ XI11_4/XI0/XI0_34/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_2 XI11_4/net21_13_ xsel_34_ XI11_4/XI0/XI0_34/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_1 XI11_4/net21_14_ xsel_34_ XI11_4/XI0/XI0_34/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN0_0 XI11_4/net21_15_ xsel_34_ XI11_4/XI0/XI0_34/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_15 XI11_4/XI0/XI0_34/d__15_ xsel_34_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_14 XI11_4/XI0/XI0_34/d__14_ xsel_34_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_13 XI11_4/XI0/XI0_34/d__13_ xsel_34_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_12 XI11_4/XI0/XI0_34/d__12_ xsel_34_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_11 XI11_4/XI0/XI0_34/d__11_ xsel_34_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_10 XI11_4/XI0/XI0_34/d__10_ xsel_34_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_9 XI11_4/XI0/XI0_34/d__9_ xsel_34_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_8 XI11_4/XI0/XI0_34/d__8_ xsel_34_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_7 XI11_4/XI0/XI0_34/d__7_ xsel_34_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_6 XI11_4/XI0/XI0_34/d__6_ xsel_34_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_5 XI11_4/XI0/XI0_34/d__5_ xsel_34_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_4 XI11_4/XI0/XI0_34/d__4_ xsel_34_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_3 XI11_4/XI0/XI0_34/d__3_ xsel_34_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_2 XI11_4/XI0/XI0_34/d__2_ xsel_34_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_1 XI11_4/XI0/XI0_34/d__1_ xsel_34_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_34/MN1_0 XI11_4/XI0/XI0_34/d__0_ xsel_34_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_15 XI11_4/net21_0_ xsel_33_ XI11_4/XI0/XI0_33/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_14 XI11_4/net21_1_ xsel_33_ XI11_4/XI0/XI0_33/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_13 XI11_4/net21_2_ xsel_33_ XI11_4/XI0/XI0_33/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_12 XI11_4/net21_3_ xsel_33_ XI11_4/XI0/XI0_33/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_11 XI11_4/net21_4_ xsel_33_ XI11_4/XI0/XI0_33/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_10 XI11_4/net21_5_ xsel_33_ XI11_4/XI0/XI0_33/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_9 XI11_4/net21_6_ xsel_33_ XI11_4/XI0/XI0_33/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_8 XI11_4/net21_7_ xsel_33_ XI11_4/XI0/XI0_33/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_7 XI11_4/net21_8_ xsel_33_ XI11_4/XI0/XI0_33/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_6 XI11_4/net21_9_ xsel_33_ XI11_4/XI0/XI0_33/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_5 XI11_4/net21_10_ xsel_33_ XI11_4/XI0/XI0_33/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_4 XI11_4/net21_11_ xsel_33_ XI11_4/XI0/XI0_33/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_3 XI11_4/net21_12_ xsel_33_ XI11_4/XI0/XI0_33/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_2 XI11_4/net21_13_ xsel_33_ XI11_4/XI0/XI0_33/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_1 XI11_4/net21_14_ xsel_33_ XI11_4/XI0/XI0_33/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN0_0 XI11_4/net21_15_ xsel_33_ XI11_4/XI0/XI0_33/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_15 XI11_4/XI0/XI0_33/d__15_ xsel_33_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_14 XI11_4/XI0/XI0_33/d__14_ xsel_33_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_13 XI11_4/XI0/XI0_33/d__13_ xsel_33_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_12 XI11_4/XI0/XI0_33/d__12_ xsel_33_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_11 XI11_4/XI0/XI0_33/d__11_ xsel_33_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_10 XI11_4/XI0/XI0_33/d__10_ xsel_33_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_9 XI11_4/XI0/XI0_33/d__9_ xsel_33_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_8 XI11_4/XI0/XI0_33/d__8_ xsel_33_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_7 XI11_4/XI0/XI0_33/d__7_ xsel_33_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_6 XI11_4/XI0/XI0_33/d__6_ xsel_33_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_5 XI11_4/XI0/XI0_33/d__5_ xsel_33_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_4 XI11_4/XI0/XI0_33/d__4_ xsel_33_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_3 XI11_4/XI0/XI0_33/d__3_ xsel_33_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_2 XI11_4/XI0/XI0_33/d__2_ xsel_33_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_1 XI11_4/XI0/XI0_33/d__1_ xsel_33_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_33/MN1_0 XI11_4/XI0/XI0_33/d__0_ xsel_33_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_15 XI11_4/net21_0_ xsel_32_ XI11_4/XI0/XI0_32/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_14 XI11_4/net21_1_ xsel_32_ XI11_4/XI0/XI0_32/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_13 XI11_4/net21_2_ xsel_32_ XI11_4/XI0/XI0_32/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_12 XI11_4/net21_3_ xsel_32_ XI11_4/XI0/XI0_32/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_11 XI11_4/net21_4_ xsel_32_ XI11_4/XI0/XI0_32/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_10 XI11_4/net21_5_ xsel_32_ XI11_4/XI0/XI0_32/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_9 XI11_4/net21_6_ xsel_32_ XI11_4/XI0/XI0_32/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_8 XI11_4/net21_7_ xsel_32_ XI11_4/XI0/XI0_32/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_7 XI11_4/net21_8_ xsel_32_ XI11_4/XI0/XI0_32/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_6 XI11_4/net21_9_ xsel_32_ XI11_4/XI0/XI0_32/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_5 XI11_4/net21_10_ xsel_32_ XI11_4/XI0/XI0_32/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_4 XI11_4/net21_11_ xsel_32_ XI11_4/XI0/XI0_32/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_3 XI11_4/net21_12_ xsel_32_ XI11_4/XI0/XI0_32/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_2 XI11_4/net21_13_ xsel_32_ XI11_4/XI0/XI0_32/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_1 XI11_4/net21_14_ xsel_32_ XI11_4/XI0/XI0_32/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN0_0 XI11_4/net21_15_ xsel_32_ XI11_4/XI0/XI0_32/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_15 XI11_4/XI0/XI0_32/d__15_ xsel_32_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_14 XI11_4/XI0/XI0_32/d__14_ xsel_32_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_13 XI11_4/XI0/XI0_32/d__13_ xsel_32_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_12 XI11_4/XI0/XI0_32/d__12_ xsel_32_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_11 XI11_4/XI0/XI0_32/d__11_ xsel_32_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_10 XI11_4/XI0/XI0_32/d__10_ xsel_32_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_9 XI11_4/XI0/XI0_32/d__9_ xsel_32_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_8 XI11_4/XI0/XI0_32/d__8_ xsel_32_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_7 XI11_4/XI0/XI0_32/d__7_ xsel_32_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_6 XI11_4/XI0/XI0_32/d__6_ xsel_32_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_5 XI11_4/XI0/XI0_32/d__5_ xsel_32_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_4 XI11_4/XI0/XI0_32/d__4_ xsel_32_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_3 XI11_4/XI0/XI0_32/d__3_ xsel_32_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_2 XI11_4/XI0/XI0_32/d__2_ xsel_32_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_1 XI11_4/XI0/XI0_32/d__1_ xsel_32_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_32/MN1_0 XI11_4/XI0/XI0_32/d__0_ xsel_32_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_15 XI11_4/net21_0_ xsel_31_ XI11_4/XI0/XI0_31/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_14 XI11_4/net21_1_ xsel_31_ XI11_4/XI0/XI0_31/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_13 XI11_4/net21_2_ xsel_31_ XI11_4/XI0/XI0_31/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_12 XI11_4/net21_3_ xsel_31_ XI11_4/XI0/XI0_31/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_11 XI11_4/net21_4_ xsel_31_ XI11_4/XI0/XI0_31/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_10 XI11_4/net21_5_ xsel_31_ XI11_4/XI0/XI0_31/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_9 XI11_4/net21_6_ xsel_31_ XI11_4/XI0/XI0_31/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_8 XI11_4/net21_7_ xsel_31_ XI11_4/XI0/XI0_31/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_7 XI11_4/net21_8_ xsel_31_ XI11_4/XI0/XI0_31/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_6 XI11_4/net21_9_ xsel_31_ XI11_4/XI0/XI0_31/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_5 XI11_4/net21_10_ xsel_31_ XI11_4/XI0/XI0_31/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_4 XI11_4/net21_11_ xsel_31_ XI11_4/XI0/XI0_31/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_3 XI11_4/net21_12_ xsel_31_ XI11_4/XI0/XI0_31/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_2 XI11_4/net21_13_ xsel_31_ XI11_4/XI0/XI0_31/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_1 XI11_4/net21_14_ xsel_31_ XI11_4/XI0/XI0_31/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN0_0 XI11_4/net21_15_ xsel_31_ XI11_4/XI0/XI0_31/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_15 XI11_4/XI0/XI0_31/d__15_ xsel_31_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_14 XI11_4/XI0/XI0_31/d__14_ xsel_31_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_13 XI11_4/XI0/XI0_31/d__13_ xsel_31_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_12 XI11_4/XI0/XI0_31/d__12_ xsel_31_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_11 XI11_4/XI0/XI0_31/d__11_ xsel_31_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_10 XI11_4/XI0/XI0_31/d__10_ xsel_31_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_9 XI11_4/XI0/XI0_31/d__9_ xsel_31_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_8 XI11_4/XI0/XI0_31/d__8_ xsel_31_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_7 XI11_4/XI0/XI0_31/d__7_ xsel_31_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_6 XI11_4/XI0/XI0_31/d__6_ xsel_31_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_5 XI11_4/XI0/XI0_31/d__5_ xsel_31_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_4 XI11_4/XI0/XI0_31/d__4_ xsel_31_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_3 XI11_4/XI0/XI0_31/d__3_ xsel_31_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_2 XI11_4/XI0/XI0_31/d__2_ xsel_31_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_1 XI11_4/XI0/XI0_31/d__1_ xsel_31_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_31/MN1_0 XI11_4/XI0/XI0_31/d__0_ xsel_31_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_15 XI11_4/net21_0_ xsel_30_ XI11_4/XI0/XI0_30/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_14 XI11_4/net21_1_ xsel_30_ XI11_4/XI0/XI0_30/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_13 XI11_4/net21_2_ xsel_30_ XI11_4/XI0/XI0_30/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_12 XI11_4/net21_3_ xsel_30_ XI11_4/XI0/XI0_30/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_11 XI11_4/net21_4_ xsel_30_ XI11_4/XI0/XI0_30/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_10 XI11_4/net21_5_ xsel_30_ XI11_4/XI0/XI0_30/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_9 XI11_4/net21_6_ xsel_30_ XI11_4/XI0/XI0_30/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_8 XI11_4/net21_7_ xsel_30_ XI11_4/XI0/XI0_30/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_7 XI11_4/net21_8_ xsel_30_ XI11_4/XI0/XI0_30/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_6 XI11_4/net21_9_ xsel_30_ XI11_4/XI0/XI0_30/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_5 XI11_4/net21_10_ xsel_30_ XI11_4/XI0/XI0_30/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_4 XI11_4/net21_11_ xsel_30_ XI11_4/XI0/XI0_30/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_3 XI11_4/net21_12_ xsel_30_ XI11_4/XI0/XI0_30/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_2 XI11_4/net21_13_ xsel_30_ XI11_4/XI0/XI0_30/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_1 XI11_4/net21_14_ xsel_30_ XI11_4/XI0/XI0_30/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN0_0 XI11_4/net21_15_ xsel_30_ XI11_4/XI0/XI0_30/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_15 XI11_4/XI0/XI0_30/d__15_ xsel_30_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_14 XI11_4/XI0/XI0_30/d__14_ xsel_30_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_13 XI11_4/XI0/XI0_30/d__13_ xsel_30_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_12 XI11_4/XI0/XI0_30/d__12_ xsel_30_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_11 XI11_4/XI0/XI0_30/d__11_ xsel_30_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_10 XI11_4/XI0/XI0_30/d__10_ xsel_30_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_9 XI11_4/XI0/XI0_30/d__9_ xsel_30_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_8 XI11_4/XI0/XI0_30/d__8_ xsel_30_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_7 XI11_4/XI0/XI0_30/d__7_ xsel_30_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_6 XI11_4/XI0/XI0_30/d__6_ xsel_30_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_5 XI11_4/XI0/XI0_30/d__5_ xsel_30_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_4 XI11_4/XI0/XI0_30/d__4_ xsel_30_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_3 XI11_4/XI0/XI0_30/d__3_ xsel_30_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_2 XI11_4/XI0/XI0_30/d__2_ xsel_30_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_1 XI11_4/XI0/XI0_30/d__1_ xsel_30_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_30/MN1_0 XI11_4/XI0/XI0_30/d__0_ xsel_30_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_15 XI11_4/net21_0_ xsel_29_ XI11_4/XI0/XI0_29/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_14 XI11_4/net21_1_ xsel_29_ XI11_4/XI0/XI0_29/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_13 XI11_4/net21_2_ xsel_29_ XI11_4/XI0/XI0_29/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_12 XI11_4/net21_3_ xsel_29_ XI11_4/XI0/XI0_29/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_11 XI11_4/net21_4_ xsel_29_ XI11_4/XI0/XI0_29/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_10 XI11_4/net21_5_ xsel_29_ XI11_4/XI0/XI0_29/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_9 XI11_4/net21_6_ xsel_29_ XI11_4/XI0/XI0_29/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_8 XI11_4/net21_7_ xsel_29_ XI11_4/XI0/XI0_29/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_7 XI11_4/net21_8_ xsel_29_ XI11_4/XI0/XI0_29/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_6 XI11_4/net21_9_ xsel_29_ XI11_4/XI0/XI0_29/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_5 XI11_4/net21_10_ xsel_29_ XI11_4/XI0/XI0_29/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_4 XI11_4/net21_11_ xsel_29_ XI11_4/XI0/XI0_29/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_3 XI11_4/net21_12_ xsel_29_ XI11_4/XI0/XI0_29/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_2 XI11_4/net21_13_ xsel_29_ XI11_4/XI0/XI0_29/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_1 XI11_4/net21_14_ xsel_29_ XI11_4/XI0/XI0_29/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN0_0 XI11_4/net21_15_ xsel_29_ XI11_4/XI0/XI0_29/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_15 XI11_4/XI0/XI0_29/d__15_ xsel_29_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_14 XI11_4/XI0/XI0_29/d__14_ xsel_29_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_13 XI11_4/XI0/XI0_29/d__13_ xsel_29_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_12 XI11_4/XI0/XI0_29/d__12_ xsel_29_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_11 XI11_4/XI0/XI0_29/d__11_ xsel_29_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_10 XI11_4/XI0/XI0_29/d__10_ xsel_29_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_9 XI11_4/XI0/XI0_29/d__9_ xsel_29_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_8 XI11_4/XI0/XI0_29/d__8_ xsel_29_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_7 XI11_4/XI0/XI0_29/d__7_ xsel_29_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_6 XI11_4/XI0/XI0_29/d__6_ xsel_29_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_5 XI11_4/XI0/XI0_29/d__5_ xsel_29_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_4 XI11_4/XI0/XI0_29/d__4_ xsel_29_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_3 XI11_4/XI0/XI0_29/d__3_ xsel_29_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_2 XI11_4/XI0/XI0_29/d__2_ xsel_29_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_1 XI11_4/XI0/XI0_29/d__1_ xsel_29_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_29/MN1_0 XI11_4/XI0/XI0_29/d__0_ xsel_29_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_15 XI11_4/net21_0_ xsel_28_ XI11_4/XI0/XI0_28/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_14 XI11_4/net21_1_ xsel_28_ XI11_4/XI0/XI0_28/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_13 XI11_4/net21_2_ xsel_28_ XI11_4/XI0/XI0_28/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_12 XI11_4/net21_3_ xsel_28_ XI11_4/XI0/XI0_28/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_11 XI11_4/net21_4_ xsel_28_ XI11_4/XI0/XI0_28/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_10 XI11_4/net21_5_ xsel_28_ XI11_4/XI0/XI0_28/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_9 XI11_4/net21_6_ xsel_28_ XI11_4/XI0/XI0_28/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_8 XI11_4/net21_7_ xsel_28_ XI11_4/XI0/XI0_28/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_7 XI11_4/net21_8_ xsel_28_ XI11_4/XI0/XI0_28/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_6 XI11_4/net21_9_ xsel_28_ XI11_4/XI0/XI0_28/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_5 XI11_4/net21_10_ xsel_28_ XI11_4/XI0/XI0_28/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_4 XI11_4/net21_11_ xsel_28_ XI11_4/XI0/XI0_28/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_3 XI11_4/net21_12_ xsel_28_ XI11_4/XI0/XI0_28/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_2 XI11_4/net21_13_ xsel_28_ XI11_4/XI0/XI0_28/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_1 XI11_4/net21_14_ xsel_28_ XI11_4/XI0/XI0_28/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN0_0 XI11_4/net21_15_ xsel_28_ XI11_4/XI0/XI0_28/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_15 XI11_4/XI0/XI0_28/d__15_ xsel_28_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_14 XI11_4/XI0/XI0_28/d__14_ xsel_28_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_13 XI11_4/XI0/XI0_28/d__13_ xsel_28_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_12 XI11_4/XI0/XI0_28/d__12_ xsel_28_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_11 XI11_4/XI0/XI0_28/d__11_ xsel_28_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_10 XI11_4/XI0/XI0_28/d__10_ xsel_28_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_9 XI11_4/XI0/XI0_28/d__9_ xsel_28_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_8 XI11_4/XI0/XI0_28/d__8_ xsel_28_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_7 XI11_4/XI0/XI0_28/d__7_ xsel_28_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_6 XI11_4/XI0/XI0_28/d__6_ xsel_28_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_5 XI11_4/XI0/XI0_28/d__5_ xsel_28_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_4 XI11_4/XI0/XI0_28/d__4_ xsel_28_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_3 XI11_4/XI0/XI0_28/d__3_ xsel_28_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_2 XI11_4/XI0/XI0_28/d__2_ xsel_28_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_1 XI11_4/XI0/XI0_28/d__1_ xsel_28_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_28/MN1_0 XI11_4/XI0/XI0_28/d__0_ xsel_28_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_15 XI11_4/net21_0_ xsel_27_ XI11_4/XI0/XI0_27/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_14 XI11_4/net21_1_ xsel_27_ XI11_4/XI0/XI0_27/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_13 XI11_4/net21_2_ xsel_27_ XI11_4/XI0/XI0_27/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_12 XI11_4/net21_3_ xsel_27_ XI11_4/XI0/XI0_27/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_11 XI11_4/net21_4_ xsel_27_ XI11_4/XI0/XI0_27/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_10 XI11_4/net21_5_ xsel_27_ XI11_4/XI0/XI0_27/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_9 XI11_4/net21_6_ xsel_27_ XI11_4/XI0/XI0_27/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_8 XI11_4/net21_7_ xsel_27_ XI11_4/XI0/XI0_27/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_7 XI11_4/net21_8_ xsel_27_ XI11_4/XI0/XI0_27/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_6 XI11_4/net21_9_ xsel_27_ XI11_4/XI0/XI0_27/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_5 XI11_4/net21_10_ xsel_27_ XI11_4/XI0/XI0_27/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_4 XI11_4/net21_11_ xsel_27_ XI11_4/XI0/XI0_27/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_3 XI11_4/net21_12_ xsel_27_ XI11_4/XI0/XI0_27/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_2 XI11_4/net21_13_ xsel_27_ XI11_4/XI0/XI0_27/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_1 XI11_4/net21_14_ xsel_27_ XI11_4/XI0/XI0_27/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN0_0 XI11_4/net21_15_ xsel_27_ XI11_4/XI0/XI0_27/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_15 XI11_4/XI0/XI0_27/d__15_ xsel_27_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_14 XI11_4/XI0/XI0_27/d__14_ xsel_27_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_13 XI11_4/XI0/XI0_27/d__13_ xsel_27_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_12 XI11_4/XI0/XI0_27/d__12_ xsel_27_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_11 XI11_4/XI0/XI0_27/d__11_ xsel_27_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_10 XI11_4/XI0/XI0_27/d__10_ xsel_27_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_9 XI11_4/XI0/XI0_27/d__9_ xsel_27_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_8 XI11_4/XI0/XI0_27/d__8_ xsel_27_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_7 XI11_4/XI0/XI0_27/d__7_ xsel_27_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_6 XI11_4/XI0/XI0_27/d__6_ xsel_27_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_5 XI11_4/XI0/XI0_27/d__5_ xsel_27_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_4 XI11_4/XI0/XI0_27/d__4_ xsel_27_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_3 XI11_4/XI0/XI0_27/d__3_ xsel_27_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_2 XI11_4/XI0/XI0_27/d__2_ xsel_27_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_1 XI11_4/XI0/XI0_27/d__1_ xsel_27_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_27/MN1_0 XI11_4/XI0/XI0_27/d__0_ xsel_27_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_15 XI11_4/net21_0_ xsel_26_ XI11_4/XI0/XI0_26/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_14 XI11_4/net21_1_ xsel_26_ XI11_4/XI0/XI0_26/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_13 XI11_4/net21_2_ xsel_26_ XI11_4/XI0/XI0_26/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_12 XI11_4/net21_3_ xsel_26_ XI11_4/XI0/XI0_26/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_11 XI11_4/net21_4_ xsel_26_ XI11_4/XI0/XI0_26/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_10 XI11_4/net21_5_ xsel_26_ XI11_4/XI0/XI0_26/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_9 XI11_4/net21_6_ xsel_26_ XI11_4/XI0/XI0_26/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_8 XI11_4/net21_7_ xsel_26_ XI11_4/XI0/XI0_26/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_7 XI11_4/net21_8_ xsel_26_ XI11_4/XI0/XI0_26/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_6 XI11_4/net21_9_ xsel_26_ XI11_4/XI0/XI0_26/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_5 XI11_4/net21_10_ xsel_26_ XI11_4/XI0/XI0_26/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_4 XI11_4/net21_11_ xsel_26_ XI11_4/XI0/XI0_26/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_3 XI11_4/net21_12_ xsel_26_ XI11_4/XI0/XI0_26/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_2 XI11_4/net21_13_ xsel_26_ XI11_4/XI0/XI0_26/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_1 XI11_4/net21_14_ xsel_26_ XI11_4/XI0/XI0_26/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN0_0 XI11_4/net21_15_ xsel_26_ XI11_4/XI0/XI0_26/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_15 XI11_4/XI0/XI0_26/d__15_ xsel_26_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_14 XI11_4/XI0/XI0_26/d__14_ xsel_26_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_13 XI11_4/XI0/XI0_26/d__13_ xsel_26_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_12 XI11_4/XI0/XI0_26/d__12_ xsel_26_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_11 XI11_4/XI0/XI0_26/d__11_ xsel_26_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_10 XI11_4/XI0/XI0_26/d__10_ xsel_26_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_9 XI11_4/XI0/XI0_26/d__9_ xsel_26_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_8 XI11_4/XI0/XI0_26/d__8_ xsel_26_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_7 XI11_4/XI0/XI0_26/d__7_ xsel_26_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_6 XI11_4/XI0/XI0_26/d__6_ xsel_26_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_5 XI11_4/XI0/XI0_26/d__5_ xsel_26_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_4 XI11_4/XI0/XI0_26/d__4_ xsel_26_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_3 XI11_4/XI0/XI0_26/d__3_ xsel_26_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_2 XI11_4/XI0/XI0_26/d__2_ xsel_26_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_1 XI11_4/XI0/XI0_26/d__1_ xsel_26_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_26/MN1_0 XI11_4/XI0/XI0_26/d__0_ xsel_26_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_15 XI11_4/net21_0_ xsel_25_ XI11_4/XI0/XI0_25/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_14 XI11_4/net21_1_ xsel_25_ XI11_4/XI0/XI0_25/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_13 XI11_4/net21_2_ xsel_25_ XI11_4/XI0/XI0_25/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_12 XI11_4/net21_3_ xsel_25_ XI11_4/XI0/XI0_25/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_11 XI11_4/net21_4_ xsel_25_ XI11_4/XI0/XI0_25/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_10 XI11_4/net21_5_ xsel_25_ XI11_4/XI0/XI0_25/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_9 XI11_4/net21_6_ xsel_25_ XI11_4/XI0/XI0_25/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_8 XI11_4/net21_7_ xsel_25_ XI11_4/XI0/XI0_25/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_7 XI11_4/net21_8_ xsel_25_ XI11_4/XI0/XI0_25/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_6 XI11_4/net21_9_ xsel_25_ XI11_4/XI0/XI0_25/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_5 XI11_4/net21_10_ xsel_25_ XI11_4/XI0/XI0_25/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_4 XI11_4/net21_11_ xsel_25_ XI11_4/XI0/XI0_25/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_3 XI11_4/net21_12_ xsel_25_ XI11_4/XI0/XI0_25/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_2 XI11_4/net21_13_ xsel_25_ XI11_4/XI0/XI0_25/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_1 XI11_4/net21_14_ xsel_25_ XI11_4/XI0/XI0_25/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN0_0 XI11_4/net21_15_ xsel_25_ XI11_4/XI0/XI0_25/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_15 XI11_4/XI0/XI0_25/d__15_ xsel_25_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_14 XI11_4/XI0/XI0_25/d__14_ xsel_25_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_13 XI11_4/XI0/XI0_25/d__13_ xsel_25_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_12 XI11_4/XI0/XI0_25/d__12_ xsel_25_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_11 XI11_4/XI0/XI0_25/d__11_ xsel_25_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_10 XI11_4/XI0/XI0_25/d__10_ xsel_25_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_9 XI11_4/XI0/XI0_25/d__9_ xsel_25_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_8 XI11_4/XI0/XI0_25/d__8_ xsel_25_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_7 XI11_4/XI0/XI0_25/d__7_ xsel_25_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_6 XI11_4/XI0/XI0_25/d__6_ xsel_25_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_5 XI11_4/XI0/XI0_25/d__5_ xsel_25_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_4 XI11_4/XI0/XI0_25/d__4_ xsel_25_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_3 XI11_4/XI0/XI0_25/d__3_ xsel_25_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_2 XI11_4/XI0/XI0_25/d__2_ xsel_25_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_1 XI11_4/XI0/XI0_25/d__1_ xsel_25_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_25/MN1_0 XI11_4/XI0/XI0_25/d__0_ xsel_25_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_15 XI11_4/net21_0_ xsel_24_ XI11_4/XI0/XI0_24/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_14 XI11_4/net21_1_ xsel_24_ XI11_4/XI0/XI0_24/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_13 XI11_4/net21_2_ xsel_24_ XI11_4/XI0/XI0_24/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_12 XI11_4/net21_3_ xsel_24_ XI11_4/XI0/XI0_24/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_11 XI11_4/net21_4_ xsel_24_ XI11_4/XI0/XI0_24/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_10 XI11_4/net21_5_ xsel_24_ XI11_4/XI0/XI0_24/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_9 XI11_4/net21_6_ xsel_24_ XI11_4/XI0/XI0_24/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_8 XI11_4/net21_7_ xsel_24_ XI11_4/XI0/XI0_24/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_7 XI11_4/net21_8_ xsel_24_ XI11_4/XI0/XI0_24/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_6 XI11_4/net21_9_ xsel_24_ XI11_4/XI0/XI0_24/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_5 XI11_4/net21_10_ xsel_24_ XI11_4/XI0/XI0_24/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_4 XI11_4/net21_11_ xsel_24_ XI11_4/XI0/XI0_24/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_3 XI11_4/net21_12_ xsel_24_ XI11_4/XI0/XI0_24/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_2 XI11_4/net21_13_ xsel_24_ XI11_4/XI0/XI0_24/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_1 XI11_4/net21_14_ xsel_24_ XI11_4/XI0/XI0_24/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN0_0 XI11_4/net21_15_ xsel_24_ XI11_4/XI0/XI0_24/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_15 XI11_4/XI0/XI0_24/d__15_ xsel_24_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_14 XI11_4/XI0/XI0_24/d__14_ xsel_24_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_13 XI11_4/XI0/XI0_24/d__13_ xsel_24_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_12 XI11_4/XI0/XI0_24/d__12_ xsel_24_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_11 XI11_4/XI0/XI0_24/d__11_ xsel_24_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_10 XI11_4/XI0/XI0_24/d__10_ xsel_24_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_9 XI11_4/XI0/XI0_24/d__9_ xsel_24_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_8 XI11_4/XI0/XI0_24/d__8_ xsel_24_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_7 XI11_4/XI0/XI0_24/d__7_ xsel_24_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_6 XI11_4/XI0/XI0_24/d__6_ xsel_24_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_5 XI11_4/XI0/XI0_24/d__5_ xsel_24_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_4 XI11_4/XI0/XI0_24/d__4_ xsel_24_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_3 XI11_4/XI0/XI0_24/d__3_ xsel_24_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_2 XI11_4/XI0/XI0_24/d__2_ xsel_24_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_1 XI11_4/XI0/XI0_24/d__1_ xsel_24_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_24/MN1_0 XI11_4/XI0/XI0_24/d__0_ xsel_24_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_15 XI11_4/net21_0_ xsel_23_ XI11_4/XI0/XI0_23/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_14 XI11_4/net21_1_ xsel_23_ XI11_4/XI0/XI0_23/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_13 XI11_4/net21_2_ xsel_23_ XI11_4/XI0/XI0_23/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_12 XI11_4/net21_3_ xsel_23_ XI11_4/XI0/XI0_23/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_11 XI11_4/net21_4_ xsel_23_ XI11_4/XI0/XI0_23/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_10 XI11_4/net21_5_ xsel_23_ XI11_4/XI0/XI0_23/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_9 XI11_4/net21_6_ xsel_23_ XI11_4/XI0/XI0_23/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_8 XI11_4/net21_7_ xsel_23_ XI11_4/XI0/XI0_23/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_7 XI11_4/net21_8_ xsel_23_ XI11_4/XI0/XI0_23/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_6 XI11_4/net21_9_ xsel_23_ XI11_4/XI0/XI0_23/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_5 XI11_4/net21_10_ xsel_23_ XI11_4/XI0/XI0_23/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_4 XI11_4/net21_11_ xsel_23_ XI11_4/XI0/XI0_23/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_3 XI11_4/net21_12_ xsel_23_ XI11_4/XI0/XI0_23/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_2 XI11_4/net21_13_ xsel_23_ XI11_4/XI0/XI0_23/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_1 XI11_4/net21_14_ xsel_23_ XI11_4/XI0/XI0_23/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN0_0 XI11_4/net21_15_ xsel_23_ XI11_4/XI0/XI0_23/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_15 XI11_4/XI0/XI0_23/d__15_ xsel_23_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_14 XI11_4/XI0/XI0_23/d__14_ xsel_23_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_13 XI11_4/XI0/XI0_23/d__13_ xsel_23_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_12 XI11_4/XI0/XI0_23/d__12_ xsel_23_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_11 XI11_4/XI0/XI0_23/d__11_ xsel_23_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_10 XI11_4/XI0/XI0_23/d__10_ xsel_23_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_9 XI11_4/XI0/XI0_23/d__9_ xsel_23_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_8 XI11_4/XI0/XI0_23/d__8_ xsel_23_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_7 XI11_4/XI0/XI0_23/d__7_ xsel_23_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_6 XI11_4/XI0/XI0_23/d__6_ xsel_23_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_5 XI11_4/XI0/XI0_23/d__5_ xsel_23_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_4 XI11_4/XI0/XI0_23/d__4_ xsel_23_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_3 XI11_4/XI0/XI0_23/d__3_ xsel_23_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_2 XI11_4/XI0/XI0_23/d__2_ xsel_23_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_1 XI11_4/XI0/XI0_23/d__1_ xsel_23_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_23/MN1_0 XI11_4/XI0/XI0_23/d__0_ xsel_23_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_15 XI11_4/net21_0_ xsel_22_ XI11_4/XI0/XI0_22/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_14 XI11_4/net21_1_ xsel_22_ XI11_4/XI0/XI0_22/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_13 XI11_4/net21_2_ xsel_22_ XI11_4/XI0/XI0_22/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_12 XI11_4/net21_3_ xsel_22_ XI11_4/XI0/XI0_22/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_11 XI11_4/net21_4_ xsel_22_ XI11_4/XI0/XI0_22/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_10 XI11_4/net21_5_ xsel_22_ XI11_4/XI0/XI0_22/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_9 XI11_4/net21_6_ xsel_22_ XI11_4/XI0/XI0_22/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_8 XI11_4/net21_7_ xsel_22_ XI11_4/XI0/XI0_22/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_7 XI11_4/net21_8_ xsel_22_ XI11_4/XI0/XI0_22/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_6 XI11_4/net21_9_ xsel_22_ XI11_4/XI0/XI0_22/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_5 XI11_4/net21_10_ xsel_22_ XI11_4/XI0/XI0_22/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_4 XI11_4/net21_11_ xsel_22_ XI11_4/XI0/XI0_22/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_3 XI11_4/net21_12_ xsel_22_ XI11_4/XI0/XI0_22/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_2 XI11_4/net21_13_ xsel_22_ XI11_4/XI0/XI0_22/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_1 XI11_4/net21_14_ xsel_22_ XI11_4/XI0/XI0_22/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN0_0 XI11_4/net21_15_ xsel_22_ XI11_4/XI0/XI0_22/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_15 XI11_4/XI0/XI0_22/d__15_ xsel_22_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_14 XI11_4/XI0/XI0_22/d__14_ xsel_22_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_13 XI11_4/XI0/XI0_22/d__13_ xsel_22_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_12 XI11_4/XI0/XI0_22/d__12_ xsel_22_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_11 XI11_4/XI0/XI0_22/d__11_ xsel_22_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_10 XI11_4/XI0/XI0_22/d__10_ xsel_22_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_9 XI11_4/XI0/XI0_22/d__9_ xsel_22_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_8 XI11_4/XI0/XI0_22/d__8_ xsel_22_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_7 XI11_4/XI0/XI0_22/d__7_ xsel_22_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_6 XI11_4/XI0/XI0_22/d__6_ xsel_22_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_5 XI11_4/XI0/XI0_22/d__5_ xsel_22_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_4 XI11_4/XI0/XI0_22/d__4_ xsel_22_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_3 XI11_4/XI0/XI0_22/d__3_ xsel_22_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_2 XI11_4/XI0/XI0_22/d__2_ xsel_22_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_1 XI11_4/XI0/XI0_22/d__1_ xsel_22_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_22/MN1_0 XI11_4/XI0/XI0_22/d__0_ xsel_22_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_15 XI11_4/net21_0_ xsel_21_ XI11_4/XI0/XI0_21/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_14 XI11_4/net21_1_ xsel_21_ XI11_4/XI0/XI0_21/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_13 XI11_4/net21_2_ xsel_21_ XI11_4/XI0/XI0_21/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_12 XI11_4/net21_3_ xsel_21_ XI11_4/XI0/XI0_21/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_11 XI11_4/net21_4_ xsel_21_ XI11_4/XI0/XI0_21/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_10 XI11_4/net21_5_ xsel_21_ XI11_4/XI0/XI0_21/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_9 XI11_4/net21_6_ xsel_21_ XI11_4/XI0/XI0_21/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_8 XI11_4/net21_7_ xsel_21_ XI11_4/XI0/XI0_21/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_7 XI11_4/net21_8_ xsel_21_ XI11_4/XI0/XI0_21/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_6 XI11_4/net21_9_ xsel_21_ XI11_4/XI0/XI0_21/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_5 XI11_4/net21_10_ xsel_21_ XI11_4/XI0/XI0_21/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_4 XI11_4/net21_11_ xsel_21_ XI11_4/XI0/XI0_21/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_3 XI11_4/net21_12_ xsel_21_ XI11_4/XI0/XI0_21/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_2 XI11_4/net21_13_ xsel_21_ XI11_4/XI0/XI0_21/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_1 XI11_4/net21_14_ xsel_21_ XI11_4/XI0/XI0_21/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN0_0 XI11_4/net21_15_ xsel_21_ XI11_4/XI0/XI0_21/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_15 XI11_4/XI0/XI0_21/d__15_ xsel_21_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_14 XI11_4/XI0/XI0_21/d__14_ xsel_21_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_13 XI11_4/XI0/XI0_21/d__13_ xsel_21_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_12 XI11_4/XI0/XI0_21/d__12_ xsel_21_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_11 XI11_4/XI0/XI0_21/d__11_ xsel_21_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_10 XI11_4/XI0/XI0_21/d__10_ xsel_21_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_9 XI11_4/XI0/XI0_21/d__9_ xsel_21_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_8 XI11_4/XI0/XI0_21/d__8_ xsel_21_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_7 XI11_4/XI0/XI0_21/d__7_ xsel_21_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_6 XI11_4/XI0/XI0_21/d__6_ xsel_21_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_5 XI11_4/XI0/XI0_21/d__5_ xsel_21_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_4 XI11_4/XI0/XI0_21/d__4_ xsel_21_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_3 XI11_4/XI0/XI0_21/d__3_ xsel_21_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_2 XI11_4/XI0/XI0_21/d__2_ xsel_21_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_1 XI11_4/XI0/XI0_21/d__1_ xsel_21_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_21/MN1_0 XI11_4/XI0/XI0_21/d__0_ xsel_21_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_15 XI11_4/net21_0_ xsel_20_ XI11_4/XI0/XI0_20/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_14 XI11_4/net21_1_ xsel_20_ XI11_4/XI0/XI0_20/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_13 XI11_4/net21_2_ xsel_20_ XI11_4/XI0/XI0_20/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_12 XI11_4/net21_3_ xsel_20_ XI11_4/XI0/XI0_20/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_11 XI11_4/net21_4_ xsel_20_ XI11_4/XI0/XI0_20/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_10 XI11_4/net21_5_ xsel_20_ XI11_4/XI0/XI0_20/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_9 XI11_4/net21_6_ xsel_20_ XI11_4/XI0/XI0_20/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_8 XI11_4/net21_7_ xsel_20_ XI11_4/XI0/XI0_20/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_7 XI11_4/net21_8_ xsel_20_ XI11_4/XI0/XI0_20/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_6 XI11_4/net21_9_ xsel_20_ XI11_4/XI0/XI0_20/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_5 XI11_4/net21_10_ xsel_20_ XI11_4/XI0/XI0_20/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_4 XI11_4/net21_11_ xsel_20_ XI11_4/XI0/XI0_20/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_3 XI11_4/net21_12_ xsel_20_ XI11_4/XI0/XI0_20/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_2 XI11_4/net21_13_ xsel_20_ XI11_4/XI0/XI0_20/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_1 XI11_4/net21_14_ xsel_20_ XI11_4/XI0/XI0_20/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN0_0 XI11_4/net21_15_ xsel_20_ XI11_4/XI0/XI0_20/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_15 XI11_4/XI0/XI0_20/d__15_ xsel_20_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_14 XI11_4/XI0/XI0_20/d__14_ xsel_20_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_13 XI11_4/XI0/XI0_20/d__13_ xsel_20_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_12 XI11_4/XI0/XI0_20/d__12_ xsel_20_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_11 XI11_4/XI0/XI0_20/d__11_ xsel_20_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_10 XI11_4/XI0/XI0_20/d__10_ xsel_20_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_9 XI11_4/XI0/XI0_20/d__9_ xsel_20_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_8 XI11_4/XI0/XI0_20/d__8_ xsel_20_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_7 XI11_4/XI0/XI0_20/d__7_ xsel_20_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_6 XI11_4/XI0/XI0_20/d__6_ xsel_20_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_5 XI11_4/XI0/XI0_20/d__5_ xsel_20_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_4 XI11_4/XI0/XI0_20/d__4_ xsel_20_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_3 XI11_4/XI0/XI0_20/d__3_ xsel_20_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_2 XI11_4/XI0/XI0_20/d__2_ xsel_20_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_1 XI11_4/XI0/XI0_20/d__1_ xsel_20_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_20/MN1_0 XI11_4/XI0/XI0_20/d__0_ xsel_20_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_15 XI11_4/net21_0_ xsel_19_ XI11_4/XI0/XI0_19/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_14 XI11_4/net21_1_ xsel_19_ XI11_4/XI0/XI0_19/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_13 XI11_4/net21_2_ xsel_19_ XI11_4/XI0/XI0_19/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_12 XI11_4/net21_3_ xsel_19_ XI11_4/XI0/XI0_19/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_11 XI11_4/net21_4_ xsel_19_ XI11_4/XI0/XI0_19/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_10 XI11_4/net21_5_ xsel_19_ XI11_4/XI0/XI0_19/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_9 XI11_4/net21_6_ xsel_19_ XI11_4/XI0/XI0_19/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_8 XI11_4/net21_7_ xsel_19_ XI11_4/XI0/XI0_19/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_7 XI11_4/net21_8_ xsel_19_ XI11_4/XI0/XI0_19/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_6 XI11_4/net21_9_ xsel_19_ XI11_4/XI0/XI0_19/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_5 XI11_4/net21_10_ xsel_19_ XI11_4/XI0/XI0_19/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_4 XI11_4/net21_11_ xsel_19_ XI11_4/XI0/XI0_19/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_3 XI11_4/net21_12_ xsel_19_ XI11_4/XI0/XI0_19/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_2 XI11_4/net21_13_ xsel_19_ XI11_4/XI0/XI0_19/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_1 XI11_4/net21_14_ xsel_19_ XI11_4/XI0/XI0_19/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN0_0 XI11_4/net21_15_ xsel_19_ XI11_4/XI0/XI0_19/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_15 XI11_4/XI0/XI0_19/d__15_ xsel_19_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_14 XI11_4/XI0/XI0_19/d__14_ xsel_19_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_13 XI11_4/XI0/XI0_19/d__13_ xsel_19_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_12 XI11_4/XI0/XI0_19/d__12_ xsel_19_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_11 XI11_4/XI0/XI0_19/d__11_ xsel_19_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_10 XI11_4/XI0/XI0_19/d__10_ xsel_19_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_9 XI11_4/XI0/XI0_19/d__9_ xsel_19_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_8 XI11_4/XI0/XI0_19/d__8_ xsel_19_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_7 XI11_4/XI0/XI0_19/d__7_ xsel_19_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_6 XI11_4/XI0/XI0_19/d__6_ xsel_19_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_5 XI11_4/XI0/XI0_19/d__5_ xsel_19_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_4 XI11_4/XI0/XI0_19/d__4_ xsel_19_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_3 XI11_4/XI0/XI0_19/d__3_ xsel_19_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_2 XI11_4/XI0/XI0_19/d__2_ xsel_19_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_1 XI11_4/XI0/XI0_19/d__1_ xsel_19_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_19/MN1_0 XI11_4/XI0/XI0_19/d__0_ xsel_19_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_15 XI11_4/net21_0_ xsel_18_ XI11_4/XI0/XI0_18/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_14 XI11_4/net21_1_ xsel_18_ XI11_4/XI0/XI0_18/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_13 XI11_4/net21_2_ xsel_18_ XI11_4/XI0/XI0_18/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_12 XI11_4/net21_3_ xsel_18_ XI11_4/XI0/XI0_18/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_11 XI11_4/net21_4_ xsel_18_ XI11_4/XI0/XI0_18/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_10 XI11_4/net21_5_ xsel_18_ XI11_4/XI0/XI0_18/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_9 XI11_4/net21_6_ xsel_18_ XI11_4/XI0/XI0_18/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_8 XI11_4/net21_7_ xsel_18_ XI11_4/XI0/XI0_18/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_7 XI11_4/net21_8_ xsel_18_ XI11_4/XI0/XI0_18/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_6 XI11_4/net21_9_ xsel_18_ XI11_4/XI0/XI0_18/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_5 XI11_4/net21_10_ xsel_18_ XI11_4/XI0/XI0_18/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_4 XI11_4/net21_11_ xsel_18_ XI11_4/XI0/XI0_18/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_3 XI11_4/net21_12_ xsel_18_ XI11_4/XI0/XI0_18/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_2 XI11_4/net21_13_ xsel_18_ XI11_4/XI0/XI0_18/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_1 XI11_4/net21_14_ xsel_18_ XI11_4/XI0/XI0_18/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN0_0 XI11_4/net21_15_ xsel_18_ XI11_4/XI0/XI0_18/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_15 XI11_4/XI0/XI0_18/d__15_ xsel_18_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_14 XI11_4/XI0/XI0_18/d__14_ xsel_18_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_13 XI11_4/XI0/XI0_18/d__13_ xsel_18_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_12 XI11_4/XI0/XI0_18/d__12_ xsel_18_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_11 XI11_4/XI0/XI0_18/d__11_ xsel_18_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_10 XI11_4/XI0/XI0_18/d__10_ xsel_18_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_9 XI11_4/XI0/XI0_18/d__9_ xsel_18_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_8 XI11_4/XI0/XI0_18/d__8_ xsel_18_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_7 XI11_4/XI0/XI0_18/d__7_ xsel_18_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_6 XI11_4/XI0/XI0_18/d__6_ xsel_18_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_5 XI11_4/XI0/XI0_18/d__5_ xsel_18_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_4 XI11_4/XI0/XI0_18/d__4_ xsel_18_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_3 XI11_4/XI0/XI0_18/d__3_ xsel_18_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_2 XI11_4/XI0/XI0_18/d__2_ xsel_18_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_1 XI11_4/XI0/XI0_18/d__1_ xsel_18_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_18/MN1_0 XI11_4/XI0/XI0_18/d__0_ xsel_18_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_15 XI11_4/net21_0_ xsel_17_ XI11_4/XI0/XI0_17/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_14 XI11_4/net21_1_ xsel_17_ XI11_4/XI0/XI0_17/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_13 XI11_4/net21_2_ xsel_17_ XI11_4/XI0/XI0_17/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_12 XI11_4/net21_3_ xsel_17_ XI11_4/XI0/XI0_17/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_11 XI11_4/net21_4_ xsel_17_ XI11_4/XI0/XI0_17/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_10 XI11_4/net21_5_ xsel_17_ XI11_4/XI0/XI0_17/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_9 XI11_4/net21_6_ xsel_17_ XI11_4/XI0/XI0_17/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_8 XI11_4/net21_7_ xsel_17_ XI11_4/XI0/XI0_17/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_7 XI11_4/net21_8_ xsel_17_ XI11_4/XI0/XI0_17/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_6 XI11_4/net21_9_ xsel_17_ XI11_4/XI0/XI0_17/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_5 XI11_4/net21_10_ xsel_17_ XI11_4/XI0/XI0_17/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_4 XI11_4/net21_11_ xsel_17_ XI11_4/XI0/XI0_17/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_3 XI11_4/net21_12_ xsel_17_ XI11_4/XI0/XI0_17/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_2 XI11_4/net21_13_ xsel_17_ XI11_4/XI0/XI0_17/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_1 XI11_4/net21_14_ xsel_17_ XI11_4/XI0/XI0_17/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN0_0 XI11_4/net21_15_ xsel_17_ XI11_4/XI0/XI0_17/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_15 XI11_4/XI0/XI0_17/d__15_ xsel_17_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_14 XI11_4/XI0/XI0_17/d__14_ xsel_17_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_13 XI11_4/XI0/XI0_17/d__13_ xsel_17_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_12 XI11_4/XI0/XI0_17/d__12_ xsel_17_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_11 XI11_4/XI0/XI0_17/d__11_ xsel_17_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_10 XI11_4/XI0/XI0_17/d__10_ xsel_17_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_9 XI11_4/XI0/XI0_17/d__9_ xsel_17_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_8 XI11_4/XI0/XI0_17/d__8_ xsel_17_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_7 XI11_4/XI0/XI0_17/d__7_ xsel_17_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_6 XI11_4/XI0/XI0_17/d__6_ xsel_17_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_5 XI11_4/XI0/XI0_17/d__5_ xsel_17_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_4 XI11_4/XI0/XI0_17/d__4_ xsel_17_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_3 XI11_4/XI0/XI0_17/d__3_ xsel_17_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_2 XI11_4/XI0/XI0_17/d__2_ xsel_17_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_1 XI11_4/XI0/XI0_17/d__1_ xsel_17_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_17/MN1_0 XI11_4/XI0/XI0_17/d__0_ xsel_17_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_15 XI11_4/net21_0_ xsel_16_ XI11_4/XI0/XI0_16/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_14 XI11_4/net21_1_ xsel_16_ XI11_4/XI0/XI0_16/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_13 XI11_4/net21_2_ xsel_16_ XI11_4/XI0/XI0_16/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_12 XI11_4/net21_3_ xsel_16_ XI11_4/XI0/XI0_16/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_11 XI11_4/net21_4_ xsel_16_ XI11_4/XI0/XI0_16/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_10 XI11_4/net21_5_ xsel_16_ XI11_4/XI0/XI0_16/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_9 XI11_4/net21_6_ xsel_16_ XI11_4/XI0/XI0_16/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_8 XI11_4/net21_7_ xsel_16_ XI11_4/XI0/XI0_16/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_7 XI11_4/net21_8_ xsel_16_ XI11_4/XI0/XI0_16/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_6 XI11_4/net21_9_ xsel_16_ XI11_4/XI0/XI0_16/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_5 XI11_4/net21_10_ xsel_16_ XI11_4/XI0/XI0_16/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_4 XI11_4/net21_11_ xsel_16_ XI11_4/XI0/XI0_16/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_3 XI11_4/net21_12_ xsel_16_ XI11_4/XI0/XI0_16/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_2 XI11_4/net21_13_ xsel_16_ XI11_4/XI0/XI0_16/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_1 XI11_4/net21_14_ xsel_16_ XI11_4/XI0/XI0_16/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN0_0 XI11_4/net21_15_ xsel_16_ XI11_4/XI0/XI0_16/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_15 XI11_4/XI0/XI0_16/d__15_ xsel_16_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_14 XI11_4/XI0/XI0_16/d__14_ xsel_16_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_13 XI11_4/XI0/XI0_16/d__13_ xsel_16_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_12 XI11_4/XI0/XI0_16/d__12_ xsel_16_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_11 XI11_4/XI0/XI0_16/d__11_ xsel_16_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_10 XI11_4/XI0/XI0_16/d__10_ xsel_16_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_9 XI11_4/XI0/XI0_16/d__9_ xsel_16_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_8 XI11_4/XI0/XI0_16/d__8_ xsel_16_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_7 XI11_4/XI0/XI0_16/d__7_ xsel_16_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_6 XI11_4/XI0/XI0_16/d__6_ xsel_16_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_5 XI11_4/XI0/XI0_16/d__5_ xsel_16_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_4 XI11_4/XI0/XI0_16/d__4_ xsel_16_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_3 XI11_4/XI0/XI0_16/d__3_ xsel_16_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_2 XI11_4/XI0/XI0_16/d__2_ xsel_16_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_1 XI11_4/XI0/XI0_16/d__1_ xsel_16_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_16/MN1_0 XI11_4/XI0/XI0_16/d__0_ xsel_16_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_15 XI11_4/net21_0_ xsel_15_ XI11_4/XI0/XI0_15/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_14 XI11_4/net21_1_ xsel_15_ XI11_4/XI0/XI0_15/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_13 XI11_4/net21_2_ xsel_15_ XI11_4/XI0/XI0_15/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_12 XI11_4/net21_3_ xsel_15_ XI11_4/XI0/XI0_15/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_11 XI11_4/net21_4_ xsel_15_ XI11_4/XI0/XI0_15/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_10 XI11_4/net21_5_ xsel_15_ XI11_4/XI0/XI0_15/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_9 XI11_4/net21_6_ xsel_15_ XI11_4/XI0/XI0_15/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_8 XI11_4/net21_7_ xsel_15_ XI11_4/XI0/XI0_15/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_7 XI11_4/net21_8_ xsel_15_ XI11_4/XI0/XI0_15/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_6 XI11_4/net21_9_ xsel_15_ XI11_4/XI0/XI0_15/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_5 XI11_4/net21_10_ xsel_15_ XI11_4/XI0/XI0_15/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_4 XI11_4/net21_11_ xsel_15_ XI11_4/XI0/XI0_15/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_3 XI11_4/net21_12_ xsel_15_ XI11_4/XI0/XI0_15/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_2 XI11_4/net21_13_ xsel_15_ XI11_4/XI0/XI0_15/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_1 XI11_4/net21_14_ xsel_15_ XI11_4/XI0/XI0_15/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN0_0 XI11_4/net21_15_ xsel_15_ XI11_4/XI0/XI0_15/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_15 XI11_4/XI0/XI0_15/d__15_ xsel_15_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_14 XI11_4/XI0/XI0_15/d__14_ xsel_15_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_13 XI11_4/XI0/XI0_15/d__13_ xsel_15_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_12 XI11_4/XI0/XI0_15/d__12_ xsel_15_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_11 XI11_4/XI0/XI0_15/d__11_ xsel_15_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_10 XI11_4/XI0/XI0_15/d__10_ xsel_15_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_9 XI11_4/XI0/XI0_15/d__9_ xsel_15_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_8 XI11_4/XI0/XI0_15/d__8_ xsel_15_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_7 XI11_4/XI0/XI0_15/d__7_ xsel_15_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_6 XI11_4/XI0/XI0_15/d__6_ xsel_15_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_5 XI11_4/XI0/XI0_15/d__5_ xsel_15_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_4 XI11_4/XI0/XI0_15/d__4_ xsel_15_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_3 XI11_4/XI0/XI0_15/d__3_ xsel_15_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_2 XI11_4/XI0/XI0_15/d__2_ xsel_15_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_1 XI11_4/XI0/XI0_15/d__1_ xsel_15_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_15/MN1_0 XI11_4/XI0/XI0_15/d__0_ xsel_15_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_15 XI11_4/net21_0_ xsel_14_ XI11_4/XI0/XI0_14/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_14 XI11_4/net21_1_ xsel_14_ XI11_4/XI0/XI0_14/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_13 XI11_4/net21_2_ xsel_14_ XI11_4/XI0/XI0_14/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_12 XI11_4/net21_3_ xsel_14_ XI11_4/XI0/XI0_14/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_11 XI11_4/net21_4_ xsel_14_ XI11_4/XI0/XI0_14/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_10 XI11_4/net21_5_ xsel_14_ XI11_4/XI0/XI0_14/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_9 XI11_4/net21_6_ xsel_14_ XI11_4/XI0/XI0_14/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_8 XI11_4/net21_7_ xsel_14_ XI11_4/XI0/XI0_14/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_7 XI11_4/net21_8_ xsel_14_ XI11_4/XI0/XI0_14/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_6 XI11_4/net21_9_ xsel_14_ XI11_4/XI0/XI0_14/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_5 XI11_4/net21_10_ xsel_14_ XI11_4/XI0/XI0_14/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_4 XI11_4/net21_11_ xsel_14_ XI11_4/XI0/XI0_14/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_3 XI11_4/net21_12_ xsel_14_ XI11_4/XI0/XI0_14/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_2 XI11_4/net21_13_ xsel_14_ XI11_4/XI0/XI0_14/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_1 XI11_4/net21_14_ xsel_14_ XI11_4/XI0/XI0_14/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN0_0 XI11_4/net21_15_ xsel_14_ XI11_4/XI0/XI0_14/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_15 XI11_4/XI0/XI0_14/d__15_ xsel_14_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_14 XI11_4/XI0/XI0_14/d__14_ xsel_14_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_13 XI11_4/XI0/XI0_14/d__13_ xsel_14_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_12 XI11_4/XI0/XI0_14/d__12_ xsel_14_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_11 XI11_4/XI0/XI0_14/d__11_ xsel_14_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_10 XI11_4/XI0/XI0_14/d__10_ xsel_14_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_9 XI11_4/XI0/XI0_14/d__9_ xsel_14_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_8 XI11_4/XI0/XI0_14/d__8_ xsel_14_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_7 XI11_4/XI0/XI0_14/d__7_ xsel_14_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_6 XI11_4/XI0/XI0_14/d__6_ xsel_14_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_5 XI11_4/XI0/XI0_14/d__5_ xsel_14_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_4 XI11_4/XI0/XI0_14/d__4_ xsel_14_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_3 XI11_4/XI0/XI0_14/d__3_ xsel_14_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_2 XI11_4/XI0/XI0_14/d__2_ xsel_14_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_1 XI11_4/XI0/XI0_14/d__1_ xsel_14_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_14/MN1_0 XI11_4/XI0/XI0_14/d__0_ xsel_14_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_15 XI11_4/net21_0_ xsel_13_ XI11_4/XI0/XI0_13/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_14 XI11_4/net21_1_ xsel_13_ XI11_4/XI0/XI0_13/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_13 XI11_4/net21_2_ xsel_13_ XI11_4/XI0/XI0_13/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_12 XI11_4/net21_3_ xsel_13_ XI11_4/XI0/XI0_13/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_11 XI11_4/net21_4_ xsel_13_ XI11_4/XI0/XI0_13/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_10 XI11_4/net21_5_ xsel_13_ XI11_4/XI0/XI0_13/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_9 XI11_4/net21_6_ xsel_13_ XI11_4/XI0/XI0_13/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_8 XI11_4/net21_7_ xsel_13_ XI11_4/XI0/XI0_13/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_7 XI11_4/net21_8_ xsel_13_ XI11_4/XI0/XI0_13/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_6 XI11_4/net21_9_ xsel_13_ XI11_4/XI0/XI0_13/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_5 XI11_4/net21_10_ xsel_13_ XI11_4/XI0/XI0_13/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_4 XI11_4/net21_11_ xsel_13_ XI11_4/XI0/XI0_13/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_3 XI11_4/net21_12_ xsel_13_ XI11_4/XI0/XI0_13/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_2 XI11_4/net21_13_ xsel_13_ XI11_4/XI0/XI0_13/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_1 XI11_4/net21_14_ xsel_13_ XI11_4/XI0/XI0_13/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN0_0 XI11_4/net21_15_ xsel_13_ XI11_4/XI0/XI0_13/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_15 XI11_4/XI0/XI0_13/d__15_ xsel_13_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_14 XI11_4/XI0/XI0_13/d__14_ xsel_13_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_13 XI11_4/XI0/XI0_13/d__13_ xsel_13_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_12 XI11_4/XI0/XI0_13/d__12_ xsel_13_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_11 XI11_4/XI0/XI0_13/d__11_ xsel_13_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_10 XI11_4/XI0/XI0_13/d__10_ xsel_13_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_9 XI11_4/XI0/XI0_13/d__9_ xsel_13_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_8 XI11_4/XI0/XI0_13/d__8_ xsel_13_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_7 XI11_4/XI0/XI0_13/d__7_ xsel_13_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_6 XI11_4/XI0/XI0_13/d__6_ xsel_13_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_5 XI11_4/XI0/XI0_13/d__5_ xsel_13_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_4 XI11_4/XI0/XI0_13/d__4_ xsel_13_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_3 XI11_4/XI0/XI0_13/d__3_ xsel_13_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_2 XI11_4/XI0/XI0_13/d__2_ xsel_13_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_1 XI11_4/XI0/XI0_13/d__1_ xsel_13_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_13/MN1_0 XI11_4/XI0/XI0_13/d__0_ xsel_13_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_15 XI11_4/net21_0_ xsel_12_ XI11_4/XI0/XI0_12/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_14 XI11_4/net21_1_ xsel_12_ XI11_4/XI0/XI0_12/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_13 XI11_4/net21_2_ xsel_12_ XI11_4/XI0/XI0_12/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_12 XI11_4/net21_3_ xsel_12_ XI11_4/XI0/XI0_12/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_11 XI11_4/net21_4_ xsel_12_ XI11_4/XI0/XI0_12/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_10 XI11_4/net21_5_ xsel_12_ XI11_4/XI0/XI0_12/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_9 XI11_4/net21_6_ xsel_12_ XI11_4/XI0/XI0_12/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_8 XI11_4/net21_7_ xsel_12_ XI11_4/XI0/XI0_12/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_7 XI11_4/net21_8_ xsel_12_ XI11_4/XI0/XI0_12/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_6 XI11_4/net21_9_ xsel_12_ XI11_4/XI0/XI0_12/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_5 XI11_4/net21_10_ xsel_12_ XI11_4/XI0/XI0_12/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_4 XI11_4/net21_11_ xsel_12_ XI11_4/XI0/XI0_12/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_3 XI11_4/net21_12_ xsel_12_ XI11_4/XI0/XI0_12/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_2 XI11_4/net21_13_ xsel_12_ XI11_4/XI0/XI0_12/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_1 XI11_4/net21_14_ xsel_12_ XI11_4/XI0/XI0_12/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN0_0 XI11_4/net21_15_ xsel_12_ XI11_4/XI0/XI0_12/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_15 XI11_4/XI0/XI0_12/d__15_ xsel_12_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_14 XI11_4/XI0/XI0_12/d__14_ xsel_12_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_13 XI11_4/XI0/XI0_12/d__13_ xsel_12_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_12 XI11_4/XI0/XI0_12/d__12_ xsel_12_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_11 XI11_4/XI0/XI0_12/d__11_ xsel_12_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_10 XI11_4/XI0/XI0_12/d__10_ xsel_12_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_9 XI11_4/XI0/XI0_12/d__9_ xsel_12_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_8 XI11_4/XI0/XI0_12/d__8_ xsel_12_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_7 XI11_4/XI0/XI0_12/d__7_ xsel_12_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_6 XI11_4/XI0/XI0_12/d__6_ xsel_12_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_5 XI11_4/XI0/XI0_12/d__5_ xsel_12_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_4 XI11_4/XI0/XI0_12/d__4_ xsel_12_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_3 XI11_4/XI0/XI0_12/d__3_ xsel_12_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_2 XI11_4/XI0/XI0_12/d__2_ xsel_12_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_1 XI11_4/XI0/XI0_12/d__1_ xsel_12_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_12/MN1_0 XI11_4/XI0/XI0_12/d__0_ xsel_12_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_15 XI11_4/net21_0_ xsel_11_ XI11_4/XI0/XI0_11/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_14 XI11_4/net21_1_ xsel_11_ XI11_4/XI0/XI0_11/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_13 XI11_4/net21_2_ xsel_11_ XI11_4/XI0/XI0_11/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_12 XI11_4/net21_3_ xsel_11_ XI11_4/XI0/XI0_11/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_11 XI11_4/net21_4_ xsel_11_ XI11_4/XI0/XI0_11/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_10 XI11_4/net21_5_ xsel_11_ XI11_4/XI0/XI0_11/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_9 XI11_4/net21_6_ xsel_11_ XI11_4/XI0/XI0_11/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_8 XI11_4/net21_7_ xsel_11_ XI11_4/XI0/XI0_11/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_7 XI11_4/net21_8_ xsel_11_ XI11_4/XI0/XI0_11/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_6 XI11_4/net21_9_ xsel_11_ XI11_4/XI0/XI0_11/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_5 XI11_4/net21_10_ xsel_11_ XI11_4/XI0/XI0_11/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_4 XI11_4/net21_11_ xsel_11_ XI11_4/XI0/XI0_11/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_3 XI11_4/net21_12_ xsel_11_ XI11_4/XI0/XI0_11/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_2 XI11_4/net21_13_ xsel_11_ XI11_4/XI0/XI0_11/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_1 XI11_4/net21_14_ xsel_11_ XI11_4/XI0/XI0_11/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN0_0 XI11_4/net21_15_ xsel_11_ XI11_4/XI0/XI0_11/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_15 XI11_4/XI0/XI0_11/d__15_ xsel_11_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_14 XI11_4/XI0/XI0_11/d__14_ xsel_11_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_13 XI11_4/XI0/XI0_11/d__13_ xsel_11_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_12 XI11_4/XI0/XI0_11/d__12_ xsel_11_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_11 XI11_4/XI0/XI0_11/d__11_ xsel_11_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_10 XI11_4/XI0/XI0_11/d__10_ xsel_11_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_9 XI11_4/XI0/XI0_11/d__9_ xsel_11_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_8 XI11_4/XI0/XI0_11/d__8_ xsel_11_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_7 XI11_4/XI0/XI0_11/d__7_ xsel_11_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_6 XI11_4/XI0/XI0_11/d__6_ xsel_11_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_5 XI11_4/XI0/XI0_11/d__5_ xsel_11_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_4 XI11_4/XI0/XI0_11/d__4_ xsel_11_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_3 XI11_4/XI0/XI0_11/d__3_ xsel_11_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_2 XI11_4/XI0/XI0_11/d__2_ xsel_11_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_1 XI11_4/XI0/XI0_11/d__1_ xsel_11_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_11/MN1_0 XI11_4/XI0/XI0_11/d__0_ xsel_11_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_15 XI11_4/net21_0_ xsel_10_ XI11_4/XI0/XI0_10/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_14 XI11_4/net21_1_ xsel_10_ XI11_4/XI0/XI0_10/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_13 XI11_4/net21_2_ xsel_10_ XI11_4/XI0/XI0_10/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_12 XI11_4/net21_3_ xsel_10_ XI11_4/XI0/XI0_10/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_11 XI11_4/net21_4_ xsel_10_ XI11_4/XI0/XI0_10/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_10 XI11_4/net21_5_ xsel_10_ XI11_4/XI0/XI0_10/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_9 XI11_4/net21_6_ xsel_10_ XI11_4/XI0/XI0_10/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_8 XI11_4/net21_7_ xsel_10_ XI11_4/XI0/XI0_10/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_7 XI11_4/net21_8_ xsel_10_ XI11_4/XI0/XI0_10/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_6 XI11_4/net21_9_ xsel_10_ XI11_4/XI0/XI0_10/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_5 XI11_4/net21_10_ xsel_10_ XI11_4/XI0/XI0_10/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_4 XI11_4/net21_11_ xsel_10_ XI11_4/XI0/XI0_10/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_3 XI11_4/net21_12_ xsel_10_ XI11_4/XI0/XI0_10/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_2 XI11_4/net21_13_ xsel_10_ XI11_4/XI0/XI0_10/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_1 XI11_4/net21_14_ xsel_10_ XI11_4/XI0/XI0_10/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN0_0 XI11_4/net21_15_ xsel_10_ XI11_4/XI0/XI0_10/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_15 XI11_4/XI0/XI0_10/d__15_ xsel_10_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_14 XI11_4/XI0/XI0_10/d__14_ xsel_10_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_13 XI11_4/XI0/XI0_10/d__13_ xsel_10_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_12 XI11_4/XI0/XI0_10/d__12_ xsel_10_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_11 XI11_4/XI0/XI0_10/d__11_ xsel_10_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_10 XI11_4/XI0/XI0_10/d__10_ xsel_10_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_9 XI11_4/XI0/XI0_10/d__9_ xsel_10_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_8 XI11_4/XI0/XI0_10/d__8_ xsel_10_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_7 XI11_4/XI0/XI0_10/d__7_ xsel_10_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_6 XI11_4/XI0/XI0_10/d__6_ xsel_10_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_5 XI11_4/XI0/XI0_10/d__5_ xsel_10_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_4 XI11_4/XI0/XI0_10/d__4_ xsel_10_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_3 XI11_4/XI0/XI0_10/d__3_ xsel_10_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_2 XI11_4/XI0/XI0_10/d__2_ xsel_10_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_1 XI11_4/XI0/XI0_10/d__1_ xsel_10_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_10/MN1_0 XI11_4/XI0/XI0_10/d__0_ xsel_10_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_15 XI11_4/net21_0_ xsel_9_ XI11_4/XI0/XI0_9/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_14 XI11_4/net21_1_ xsel_9_ XI11_4/XI0/XI0_9/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_13 XI11_4/net21_2_ xsel_9_ XI11_4/XI0/XI0_9/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_12 XI11_4/net21_3_ xsel_9_ XI11_4/XI0/XI0_9/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_11 XI11_4/net21_4_ xsel_9_ XI11_4/XI0/XI0_9/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_10 XI11_4/net21_5_ xsel_9_ XI11_4/XI0/XI0_9/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_9 XI11_4/net21_6_ xsel_9_ XI11_4/XI0/XI0_9/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_8 XI11_4/net21_7_ xsel_9_ XI11_4/XI0/XI0_9/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_7 XI11_4/net21_8_ xsel_9_ XI11_4/XI0/XI0_9/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_6 XI11_4/net21_9_ xsel_9_ XI11_4/XI0/XI0_9/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_5 XI11_4/net21_10_ xsel_9_ XI11_4/XI0/XI0_9/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_4 XI11_4/net21_11_ xsel_9_ XI11_4/XI0/XI0_9/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_3 XI11_4/net21_12_ xsel_9_ XI11_4/XI0/XI0_9/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_2 XI11_4/net21_13_ xsel_9_ XI11_4/XI0/XI0_9/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_1 XI11_4/net21_14_ xsel_9_ XI11_4/XI0/XI0_9/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN0_0 XI11_4/net21_15_ xsel_9_ XI11_4/XI0/XI0_9/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_15 XI11_4/XI0/XI0_9/d__15_ xsel_9_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_14 XI11_4/XI0/XI0_9/d__14_ xsel_9_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_13 XI11_4/XI0/XI0_9/d__13_ xsel_9_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_12 XI11_4/XI0/XI0_9/d__12_ xsel_9_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_11 XI11_4/XI0/XI0_9/d__11_ xsel_9_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_10 XI11_4/XI0/XI0_9/d__10_ xsel_9_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_9 XI11_4/XI0/XI0_9/d__9_ xsel_9_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_8 XI11_4/XI0/XI0_9/d__8_ xsel_9_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_7 XI11_4/XI0/XI0_9/d__7_ xsel_9_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_6 XI11_4/XI0/XI0_9/d__6_ xsel_9_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_5 XI11_4/XI0/XI0_9/d__5_ xsel_9_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_4 XI11_4/XI0/XI0_9/d__4_ xsel_9_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_3 XI11_4/XI0/XI0_9/d__3_ xsel_9_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_2 XI11_4/XI0/XI0_9/d__2_ xsel_9_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_1 XI11_4/XI0/XI0_9/d__1_ xsel_9_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_9/MN1_0 XI11_4/XI0/XI0_9/d__0_ xsel_9_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_15 XI11_4/net21_0_ xsel_8_ XI11_4/XI0/XI0_8/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_14 XI11_4/net21_1_ xsel_8_ XI11_4/XI0/XI0_8/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_13 XI11_4/net21_2_ xsel_8_ XI11_4/XI0/XI0_8/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_12 XI11_4/net21_3_ xsel_8_ XI11_4/XI0/XI0_8/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_11 XI11_4/net21_4_ xsel_8_ XI11_4/XI0/XI0_8/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_10 XI11_4/net21_5_ xsel_8_ XI11_4/XI0/XI0_8/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_9 XI11_4/net21_6_ xsel_8_ XI11_4/XI0/XI0_8/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_8 XI11_4/net21_7_ xsel_8_ XI11_4/XI0/XI0_8/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_7 XI11_4/net21_8_ xsel_8_ XI11_4/XI0/XI0_8/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_6 XI11_4/net21_9_ xsel_8_ XI11_4/XI0/XI0_8/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_5 XI11_4/net21_10_ xsel_8_ XI11_4/XI0/XI0_8/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_4 XI11_4/net21_11_ xsel_8_ XI11_4/XI0/XI0_8/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_3 XI11_4/net21_12_ xsel_8_ XI11_4/XI0/XI0_8/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_2 XI11_4/net21_13_ xsel_8_ XI11_4/XI0/XI0_8/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_1 XI11_4/net21_14_ xsel_8_ XI11_4/XI0/XI0_8/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN0_0 XI11_4/net21_15_ xsel_8_ XI11_4/XI0/XI0_8/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_15 XI11_4/XI0/XI0_8/d__15_ xsel_8_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_14 XI11_4/XI0/XI0_8/d__14_ xsel_8_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_13 XI11_4/XI0/XI0_8/d__13_ xsel_8_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_12 XI11_4/XI0/XI0_8/d__12_ xsel_8_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_11 XI11_4/XI0/XI0_8/d__11_ xsel_8_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_10 XI11_4/XI0/XI0_8/d__10_ xsel_8_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_9 XI11_4/XI0/XI0_8/d__9_ xsel_8_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_8 XI11_4/XI0/XI0_8/d__8_ xsel_8_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_7 XI11_4/XI0/XI0_8/d__7_ xsel_8_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_6 XI11_4/XI0/XI0_8/d__6_ xsel_8_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_5 XI11_4/XI0/XI0_8/d__5_ xsel_8_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_4 XI11_4/XI0/XI0_8/d__4_ xsel_8_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_3 XI11_4/XI0/XI0_8/d__3_ xsel_8_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_2 XI11_4/XI0/XI0_8/d__2_ xsel_8_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_1 XI11_4/XI0/XI0_8/d__1_ xsel_8_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_8/MN1_0 XI11_4/XI0/XI0_8/d__0_ xsel_8_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_15 XI11_4/net21_0_ xsel_7_ XI11_4/XI0/XI0_7/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_14 XI11_4/net21_1_ xsel_7_ XI11_4/XI0/XI0_7/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_13 XI11_4/net21_2_ xsel_7_ XI11_4/XI0/XI0_7/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_12 XI11_4/net21_3_ xsel_7_ XI11_4/XI0/XI0_7/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_11 XI11_4/net21_4_ xsel_7_ XI11_4/XI0/XI0_7/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_10 XI11_4/net21_5_ xsel_7_ XI11_4/XI0/XI0_7/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_9 XI11_4/net21_6_ xsel_7_ XI11_4/XI0/XI0_7/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_8 XI11_4/net21_7_ xsel_7_ XI11_4/XI0/XI0_7/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_7 XI11_4/net21_8_ xsel_7_ XI11_4/XI0/XI0_7/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_6 XI11_4/net21_9_ xsel_7_ XI11_4/XI0/XI0_7/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_5 XI11_4/net21_10_ xsel_7_ XI11_4/XI0/XI0_7/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_4 XI11_4/net21_11_ xsel_7_ XI11_4/XI0/XI0_7/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_3 XI11_4/net21_12_ xsel_7_ XI11_4/XI0/XI0_7/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_2 XI11_4/net21_13_ xsel_7_ XI11_4/XI0/XI0_7/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_1 XI11_4/net21_14_ xsel_7_ XI11_4/XI0/XI0_7/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN0_0 XI11_4/net21_15_ xsel_7_ XI11_4/XI0/XI0_7/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_15 XI11_4/XI0/XI0_7/d__15_ xsel_7_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_14 XI11_4/XI0/XI0_7/d__14_ xsel_7_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_13 XI11_4/XI0/XI0_7/d__13_ xsel_7_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_12 XI11_4/XI0/XI0_7/d__12_ xsel_7_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_11 XI11_4/XI0/XI0_7/d__11_ xsel_7_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_10 XI11_4/XI0/XI0_7/d__10_ xsel_7_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_9 XI11_4/XI0/XI0_7/d__9_ xsel_7_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_8 XI11_4/XI0/XI0_7/d__8_ xsel_7_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_7 XI11_4/XI0/XI0_7/d__7_ xsel_7_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_6 XI11_4/XI0/XI0_7/d__6_ xsel_7_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_5 XI11_4/XI0/XI0_7/d__5_ xsel_7_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_4 XI11_4/XI0/XI0_7/d__4_ xsel_7_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_3 XI11_4/XI0/XI0_7/d__3_ xsel_7_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_2 XI11_4/XI0/XI0_7/d__2_ xsel_7_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_1 XI11_4/XI0/XI0_7/d__1_ xsel_7_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_7/MN1_0 XI11_4/XI0/XI0_7/d__0_ xsel_7_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_15 XI11_4/net21_0_ xsel_6_ XI11_4/XI0/XI0_6/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_14 XI11_4/net21_1_ xsel_6_ XI11_4/XI0/XI0_6/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_13 XI11_4/net21_2_ xsel_6_ XI11_4/XI0/XI0_6/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_12 XI11_4/net21_3_ xsel_6_ XI11_4/XI0/XI0_6/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_11 XI11_4/net21_4_ xsel_6_ XI11_4/XI0/XI0_6/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_10 XI11_4/net21_5_ xsel_6_ XI11_4/XI0/XI0_6/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_9 XI11_4/net21_6_ xsel_6_ XI11_4/XI0/XI0_6/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_8 XI11_4/net21_7_ xsel_6_ XI11_4/XI0/XI0_6/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_7 XI11_4/net21_8_ xsel_6_ XI11_4/XI0/XI0_6/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_6 XI11_4/net21_9_ xsel_6_ XI11_4/XI0/XI0_6/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_5 XI11_4/net21_10_ xsel_6_ XI11_4/XI0/XI0_6/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_4 XI11_4/net21_11_ xsel_6_ XI11_4/XI0/XI0_6/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_3 XI11_4/net21_12_ xsel_6_ XI11_4/XI0/XI0_6/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_2 XI11_4/net21_13_ xsel_6_ XI11_4/XI0/XI0_6/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_1 XI11_4/net21_14_ xsel_6_ XI11_4/XI0/XI0_6/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN0_0 XI11_4/net21_15_ xsel_6_ XI11_4/XI0/XI0_6/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_15 XI11_4/XI0/XI0_6/d__15_ xsel_6_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_14 XI11_4/XI0/XI0_6/d__14_ xsel_6_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_13 XI11_4/XI0/XI0_6/d__13_ xsel_6_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_12 XI11_4/XI0/XI0_6/d__12_ xsel_6_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_11 XI11_4/XI0/XI0_6/d__11_ xsel_6_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_10 XI11_4/XI0/XI0_6/d__10_ xsel_6_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_9 XI11_4/XI0/XI0_6/d__9_ xsel_6_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_8 XI11_4/XI0/XI0_6/d__8_ xsel_6_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_7 XI11_4/XI0/XI0_6/d__7_ xsel_6_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_6 XI11_4/XI0/XI0_6/d__6_ xsel_6_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_5 XI11_4/XI0/XI0_6/d__5_ xsel_6_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_4 XI11_4/XI0/XI0_6/d__4_ xsel_6_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_3 XI11_4/XI0/XI0_6/d__3_ xsel_6_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_2 XI11_4/XI0/XI0_6/d__2_ xsel_6_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_1 XI11_4/XI0/XI0_6/d__1_ xsel_6_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_6/MN1_0 XI11_4/XI0/XI0_6/d__0_ xsel_6_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_15 XI11_4/net21_0_ xsel_5_ XI11_4/XI0/XI0_5/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_14 XI11_4/net21_1_ xsel_5_ XI11_4/XI0/XI0_5/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_13 XI11_4/net21_2_ xsel_5_ XI11_4/XI0/XI0_5/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_12 XI11_4/net21_3_ xsel_5_ XI11_4/XI0/XI0_5/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_11 XI11_4/net21_4_ xsel_5_ XI11_4/XI0/XI0_5/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_10 XI11_4/net21_5_ xsel_5_ XI11_4/XI0/XI0_5/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_9 XI11_4/net21_6_ xsel_5_ XI11_4/XI0/XI0_5/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_8 XI11_4/net21_7_ xsel_5_ XI11_4/XI0/XI0_5/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_7 XI11_4/net21_8_ xsel_5_ XI11_4/XI0/XI0_5/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_6 XI11_4/net21_9_ xsel_5_ XI11_4/XI0/XI0_5/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_5 XI11_4/net21_10_ xsel_5_ XI11_4/XI0/XI0_5/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_4 XI11_4/net21_11_ xsel_5_ XI11_4/XI0/XI0_5/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_3 XI11_4/net21_12_ xsel_5_ XI11_4/XI0/XI0_5/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_2 XI11_4/net21_13_ xsel_5_ XI11_4/XI0/XI0_5/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_1 XI11_4/net21_14_ xsel_5_ XI11_4/XI0/XI0_5/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN0_0 XI11_4/net21_15_ xsel_5_ XI11_4/XI0/XI0_5/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_15 XI11_4/XI0/XI0_5/d__15_ xsel_5_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_14 XI11_4/XI0/XI0_5/d__14_ xsel_5_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_13 XI11_4/XI0/XI0_5/d__13_ xsel_5_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_12 XI11_4/XI0/XI0_5/d__12_ xsel_5_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_11 XI11_4/XI0/XI0_5/d__11_ xsel_5_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_10 XI11_4/XI0/XI0_5/d__10_ xsel_5_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_9 XI11_4/XI0/XI0_5/d__9_ xsel_5_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_8 XI11_4/XI0/XI0_5/d__8_ xsel_5_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_7 XI11_4/XI0/XI0_5/d__7_ xsel_5_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_6 XI11_4/XI0/XI0_5/d__6_ xsel_5_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_5 XI11_4/XI0/XI0_5/d__5_ xsel_5_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_4 XI11_4/XI0/XI0_5/d__4_ xsel_5_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_3 XI11_4/XI0/XI0_5/d__3_ xsel_5_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_2 XI11_4/XI0/XI0_5/d__2_ xsel_5_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_1 XI11_4/XI0/XI0_5/d__1_ xsel_5_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_5/MN1_0 XI11_4/XI0/XI0_5/d__0_ xsel_5_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_15 XI11_4/net21_0_ xsel_4_ XI11_4/XI0/XI0_4/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_14 XI11_4/net21_1_ xsel_4_ XI11_4/XI0/XI0_4/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_13 XI11_4/net21_2_ xsel_4_ XI11_4/XI0/XI0_4/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_12 XI11_4/net21_3_ xsel_4_ XI11_4/XI0/XI0_4/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_11 XI11_4/net21_4_ xsel_4_ XI11_4/XI0/XI0_4/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_10 XI11_4/net21_5_ xsel_4_ XI11_4/XI0/XI0_4/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_9 XI11_4/net21_6_ xsel_4_ XI11_4/XI0/XI0_4/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_8 XI11_4/net21_7_ xsel_4_ XI11_4/XI0/XI0_4/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_7 XI11_4/net21_8_ xsel_4_ XI11_4/XI0/XI0_4/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_6 XI11_4/net21_9_ xsel_4_ XI11_4/XI0/XI0_4/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_5 XI11_4/net21_10_ xsel_4_ XI11_4/XI0/XI0_4/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_4 XI11_4/net21_11_ xsel_4_ XI11_4/XI0/XI0_4/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_3 XI11_4/net21_12_ xsel_4_ XI11_4/XI0/XI0_4/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_2 XI11_4/net21_13_ xsel_4_ XI11_4/XI0/XI0_4/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_1 XI11_4/net21_14_ xsel_4_ XI11_4/XI0/XI0_4/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN0_0 XI11_4/net21_15_ xsel_4_ XI11_4/XI0/XI0_4/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_15 XI11_4/XI0/XI0_4/d__15_ xsel_4_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_14 XI11_4/XI0/XI0_4/d__14_ xsel_4_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_13 XI11_4/XI0/XI0_4/d__13_ xsel_4_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_12 XI11_4/XI0/XI0_4/d__12_ xsel_4_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_11 XI11_4/XI0/XI0_4/d__11_ xsel_4_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_10 XI11_4/XI0/XI0_4/d__10_ xsel_4_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_9 XI11_4/XI0/XI0_4/d__9_ xsel_4_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_8 XI11_4/XI0/XI0_4/d__8_ xsel_4_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_7 XI11_4/XI0/XI0_4/d__7_ xsel_4_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_6 XI11_4/XI0/XI0_4/d__6_ xsel_4_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_5 XI11_4/XI0/XI0_4/d__5_ xsel_4_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_4 XI11_4/XI0/XI0_4/d__4_ xsel_4_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_3 XI11_4/XI0/XI0_4/d__3_ xsel_4_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_2 XI11_4/XI0/XI0_4/d__2_ xsel_4_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_1 XI11_4/XI0/XI0_4/d__1_ xsel_4_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_4/MN1_0 XI11_4/XI0/XI0_4/d__0_ xsel_4_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_15 XI11_4/net21_0_ xsel_3_ XI11_4/XI0/XI0_3/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_14 XI11_4/net21_1_ xsel_3_ XI11_4/XI0/XI0_3/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_13 XI11_4/net21_2_ xsel_3_ XI11_4/XI0/XI0_3/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_12 XI11_4/net21_3_ xsel_3_ XI11_4/XI0/XI0_3/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_11 XI11_4/net21_4_ xsel_3_ XI11_4/XI0/XI0_3/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_10 XI11_4/net21_5_ xsel_3_ XI11_4/XI0/XI0_3/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_9 XI11_4/net21_6_ xsel_3_ XI11_4/XI0/XI0_3/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_8 XI11_4/net21_7_ xsel_3_ XI11_4/XI0/XI0_3/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_7 XI11_4/net21_8_ xsel_3_ XI11_4/XI0/XI0_3/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_6 XI11_4/net21_9_ xsel_3_ XI11_4/XI0/XI0_3/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_5 XI11_4/net21_10_ xsel_3_ XI11_4/XI0/XI0_3/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_4 XI11_4/net21_11_ xsel_3_ XI11_4/XI0/XI0_3/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_3 XI11_4/net21_12_ xsel_3_ XI11_4/XI0/XI0_3/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_2 XI11_4/net21_13_ xsel_3_ XI11_4/XI0/XI0_3/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_1 XI11_4/net21_14_ xsel_3_ XI11_4/XI0/XI0_3/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN0_0 XI11_4/net21_15_ xsel_3_ XI11_4/XI0/XI0_3/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_15 XI11_4/XI0/XI0_3/d__15_ xsel_3_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_14 XI11_4/XI0/XI0_3/d__14_ xsel_3_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_13 XI11_4/XI0/XI0_3/d__13_ xsel_3_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_12 XI11_4/XI0/XI0_3/d__12_ xsel_3_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_11 XI11_4/XI0/XI0_3/d__11_ xsel_3_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_10 XI11_4/XI0/XI0_3/d__10_ xsel_3_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_9 XI11_4/XI0/XI0_3/d__9_ xsel_3_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_8 XI11_4/XI0/XI0_3/d__8_ xsel_3_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_7 XI11_4/XI0/XI0_3/d__7_ xsel_3_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_6 XI11_4/XI0/XI0_3/d__6_ xsel_3_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_5 XI11_4/XI0/XI0_3/d__5_ xsel_3_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_4 XI11_4/XI0/XI0_3/d__4_ xsel_3_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_3 XI11_4/XI0/XI0_3/d__3_ xsel_3_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_2 XI11_4/XI0/XI0_3/d__2_ xsel_3_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_1 XI11_4/XI0/XI0_3/d__1_ xsel_3_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_3/MN1_0 XI11_4/XI0/XI0_3/d__0_ xsel_3_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_15 XI11_4/net21_0_ xsel_2_ XI11_4/XI0/XI0_2/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_14 XI11_4/net21_1_ xsel_2_ XI11_4/XI0/XI0_2/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_13 XI11_4/net21_2_ xsel_2_ XI11_4/XI0/XI0_2/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_12 XI11_4/net21_3_ xsel_2_ XI11_4/XI0/XI0_2/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_11 XI11_4/net21_4_ xsel_2_ XI11_4/XI0/XI0_2/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_10 XI11_4/net21_5_ xsel_2_ XI11_4/XI0/XI0_2/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_9 XI11_4/net21_6_ xsel_2_ XI11_4/XI0/XI0_2/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_8 XI11_4/net21_7_ xsel_2_ XI11_4/XI0/XI0_2/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_7 XI11_4/net21_8_ xsel_2_ XI11_4/XI0/XI0_2/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_6 XI11_4/net21_9_ xsel_2_ XI11_4/XI0/XI0_2/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_5 XI11_4/net21_10_ xsel_2_ XI11_4/XI0/XI0_2/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_4 XI11_4/net21_11_ xsel_2_ XI11_4/XI0/XI0_2/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_3 XI11_4/net21_12_ xsel_2_ XI11_4/XI0/XI0_2/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_2 XI11_4/net21_13_ xsel_2_ XI11_4/XI0/XI0_2/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_1 XI11_4/net21_14_ xsel_2_ XI11_4/XI0/XI0_2/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN0_0 XI11_4/net21_15_ xsel_2_ XI11_4/XI0/XI0_2/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_15 XI11_4/XI0/XI0_2/d__15_ xsel_2_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_14 XI11_4/XI0/XI0_2/d__14_ xsel_2_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_13 XI11_4/XI0/XI0_2/d__13_ xsel_2_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_12 XI11_4/XI0/XI0_2/d__12_ xsel_2_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_11 XI11_4/XI0/XI0_2/d__11_ xsel_2_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_10 XI11_4/XI0/XI0_2/d__10_ xsel_2_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_9 XI11_4/XI0/XI0_2/d__9_ xsel_2_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_8 XI11_4/XI0/XI0_2/d__8_ xsel_2_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_7 XI11_4/XI0/XI0_2/d__7_ xsel_2_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_6 XI11_4/XI0/XI0_2/d__6_ xsel_2_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_5 XI11_4/XI0/XI0_2/d__5_ xsel_2_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_4 XI11_4/XI0/XI0_2/d__4_ xsel_2_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_3 XI11_4/XI0/XI0_2/d__3_ xsel_2_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_2 XI11_4/XI0/XI0_2/d__2_ xsel_2_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_1 XI11_4/XI0/XI0_2/d__1_ xsel_2_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_2/MN1_0 XI11_4/XI0/XI0_2/d__0_ xsel_2_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_15 XI11_4/net21_0_ xsel_1_ XI11_4/XI0/XI0_1/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_14 XI11_4/net21_1_ xsel_1_ XI11_4/XI0/XI0_1/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_13 XI11_4/net21_2_ xsel_1_ XI11_4/XI0/XI0_1/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_12 XI11_4/net21_3_ xsel_1_ XI11_4/XI0/XI0_1/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_11 XI11_4/net21_4_ xsel_1_ XI11_4/XI0/XI0_1/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_10 XI11_4/net21_5_ xsel_1_ XI11_4/XI0/XI0_1/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_9 XI11_4/net21_6_ xsel_1_ XI11_4/XI0/XI0_1/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_8 XI11_4/net21_7_ xsel_1_ XI11_4/XI0/XI0_1/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_7 XI11_4/net21_8_ xsel_1_ XI11_4/XI0/XI0_1/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_6 XI11_4/net21_9_ xsel_1_ XI11_4/XI0/XI0_1/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_5 XI11_4/net21_10_ xsel_1_ XI11_4/XI0/XI0_1/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_4 XI11_4/net21_11_ xsel_1_ XI11_4/XI0/XI0_1/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_3 XI11_4/net21_12_ xsel_1_ XI11_4/XI0/XI0_1/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_2 XI11_4/net21_13_ xsel_1_ XI11_4/XI0/XI0_1/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_1 XI11_4/net21_14_ xsel_1_ XI11_4/XI0/XI0_1/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN0_0 XI11_4/net21_15_ xsel_1_ XI11_4/XI0/XI0_1/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_15 XI11_4/XI0/XI0_1/d__15_ xsel_1_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_14 XI11_4/XI0/XI0_1/d__14_ xsel_1_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_13 XI11_4/XI0/XI0_1/d__13_ xsel_1_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_12 XI11_4/XI0/XI0_1/d__12_ xsel_1_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_11 XI11_4/XI0/XI0_1/d__11_ xsel_1_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_10 XI11_4/XI0/XI0_1/d__10_ xsel_1_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_9 XI11_4/XI0/XI0_1/d__9_ xsel_1_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_8 XI11_4/XI0/XI0_1/d__8_ xsel_1_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_7 XI11_4/XI0/XI0_1/d__7_ xsel_1_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_6 XI11_4/XI0/XI0_1/d__6_ xsel_1_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_5 XI11_4/XI0/XI0_1/d__5_ xsel_1_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_4 XI11_4/XI0/XI0_1/d__4_ xsel_1_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_3 XI11_4/XI0/XI0_1/d__3_ xsel_1_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_2 XI11_4/XI0/XI0_1/d__2_ xsel_1_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_1 XI11_4/XI0/XI0_1/d__1_ xsel_1_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_1/MN1_0 XI11_4/XI0/XI0_1/d__0_ xsel_1_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_15 XI11_4/net21_0_ xsel_0_ XI11_4/XI0/XI0_0/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_14 XI11_4/net21_1_ xsel_0_ XI11_4/XI0/XI0_0/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_13 XI11_4/net21_2_ xsel_0_ XI11_4/XI0/XI0_0/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_12 XI11_4/net21_3_ xsel_0_ XI11_4/XI0/XI0_0/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_11 XI11_4/net21_4_ xsel_0_ XI11_4/XI0/XI0_0/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_10 XI11_4/net21_5_ xsel_0_ XI11_4/XI0/XI0_0/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_9 XI11_4/net21_6_ xsel_0_ XI11_4/XI0/XI0_0/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_8 XI11_4/net21_7_ xsel_0_ XI11_4/XI0/XI0_0/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_7 XI11_4/net21_8_ xsel_0_ XI11_4/XI0/XI0_0/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_6 XI11_4/net21_9_ xsel_0_ XI11_4/XI0/XI0_0/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_5 XI11_4/net21_10_ xsel_0_ XI11_4/XI0/XI0_0/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_4 XI11_4/net21_11_ xsel_0_ XI11_4/XI0/XI0_0/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_3 XI11_4/net21_12_ xsel_0_ XI11_4/XI0/XI0_0/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_2 XI11_4/net21_13_ xsel_0_ XI11_4/XI0/XI0_0/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_1 XI11_4/net21_14_ xsel_0_ XI11_4/XI0/XI0_0/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN0_0 XI11_4/net21_15_ xsel_0_ XI11_4/XI0/XI0_0/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_15 XI11_4/XI0/XI0_0/d__15_ xsel_0_ XI11_4/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_14 XI11_4/XI0/XI0_0/d__14_ xsel_0_ XI11_4/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_13 XI11_4/XI0/XI0_0/d__13_ xsel_0_ XI11_4/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_12 XI11_4/XI0/XI0_0/d__12_ xsel_0_ XI11_4/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_11 XI11_4/XI0/XI0_0/d__11_ xsel_0_ XI11_4/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_10 XI11_4/XI0/XI0_0/d__10_ xsel_0_ XI11_4/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_9 XI11_4/XI0/XI0_0/d__9_ xsel_0_ XI11_4/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_8 XI11_4/XI0/XI0_0/d__8_ xsel_0_ XI11_4/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_7 XI11_4/XI0/XI0_0/d__7_ xsel_0_ XI11_4/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_6 XI11_4/XI0/XI0_0/d__6_ xsel_0_ XI11_4/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_5 XI11_4/XI0/XI0_0/d__5_ xsel_0_ XI11_4/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_4 XI11_4/XI0/XI0_0/d__4_ xsel_0_ XI11_4/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_3 XI11_4/XI0/XI0_0/d__3_ xsel_0_ XI11_4/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_2 XI11_4/XI0/XI0_0/d__2_ xsel_0_ XI11_4/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_1 XI11_4/XI0/XI0_0/d__1_ xsel_0_ XI11_4/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_4/XI0/XI0_0/MN1_0 XI11_4/XI0/XI0_0/d__0_ xsel_0_ XI11_4/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI2/MN0_15 XI11_3/net21_0_ ysel_15_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_14 XI11_3/net21_1_ ysel_14_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_13 XI11_3/net21_2_ ysel_13_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_12 XI11_3/net21_3_ ysel_12_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_11 XI11_3/net21_4_ ysel_11_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_10 XI11_3/net21_5_ ysel_10_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_9 XI11_3/net21_6_ ysel_9_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_8 XI11_3/net21_7_ ysel_8_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_7 XI11_3/net21_8_ ysel_7_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_6 XI11_3/net21_9_ ysel_6_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_5 XI11_3/net21_10_ ysel_5_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_4 XI11_3/net21_11_ ysel_4_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_3 XI11_3/net21_12_ ysel_3_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_2 XI11_3/net21_13_ ysel_2_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_1 XI11_3/net21_14_ ysel_1_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN0_0 XI11_3/net21_15_ ysel_0_ XI11_3/net9 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_15 XI11_3/net20_0_ ysel_15_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_14 XI11_3/net20_1_ ysel_14_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_13 XI11_3/net20_2_ ysel_13_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_12 XI11_3/net20_3_ ysel_12_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_11 XI11_3/net20_4_ ysel_11_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_10 XI11_3/net20_5_ ysel_10_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_9 XI11_3/net20_6_ ysel_9_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_8 XI11_3/net20_7_ ysel_8_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_7 XI11_3/net20_8_ ysel_7_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_6 XI11_3/net20_9_ ysel_6_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_5 XI11_3/net20_10_ ysel_5_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_4 XI11_3/net20_11_ ysel_4_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_3 XI11_3/net20_12_ ysel_3_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_2 XI11_3/net20_13_ ysel_2_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_1 XI11_3/net20_14_ ysel_1_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI2/MN1_0 XI11_3/net20_15_ ysel_0_ XI11_3/net12 gnd MN l=1.8e-07 w=1.5e-06 $[n18ll] 
XI11_3/XI4/MN8 vdd XI11_3/XI4/net8 XI11_3/net12 vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_3/XI4/MP0 XI11_3/net9 XI11_3/XI4/net23 vdd vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_3/XI4/MP4 XI11_3/net12 XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI4/MP1 XI11_3/net9 XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI4/MP5 XI11_3/net12 XI11_3/preck XI11_3/net9 vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI4/MN7 vdd XI11_3/XI4/net090 DOUT_3_ vdd MP l=1.8e-07 w=6e-06 $[p18ll] 
XI11_3/XI4/MP3 gnd XI11_3/XI4/net089 XI11_3/net12 gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_3/XI4/MN5 XI11_3/net9 XI11_3/XI4/net0103 gnd gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_3/XI4/MN4 XI11_3/XI4/data_out_ XI11_3/XI4/net32 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_3/XI4/MN0 XI11_3/XI4/data_out XI11_3/XI4/net52 gnd gnd MN l=1.8e-07 w=1e-06 $[n18ll] 
XI11_3/XI4/MN9 gnd XI11_3/XI4/net0112 DOUT_3_ gnd MN l=1.8e-07 w=2e-06 $[n18ll] 
XI11_3/XI1_15/MP2 XI11_3/net20_0_ XI11_3/preck XI11_3/net21_0_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_15/MP1 XI11_3/net20_0_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_15/MP0 XI11_3/net21_0_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_14/MP2 XI11_3/net20_1_ XI11_3/preck XI11_3/net21_1_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_14/MP1 XI11_3/net20_1_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_14/MP0 XI11_3/net21_1_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_13/MP2 XI11_3/net20_2_ XI11_3/preck XI11_3/net21_2_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_13/MP1 XI11_3/net20_2_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_13/MP0 XI11_3/net21_2_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_12/MP2 XI11_3/net20_3_ XI11_3/preck XI11_3/net21_3_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_12/MP1 XI11_3/net20_3_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_12/MP0 XI11_3/net21_3_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_11/MP2 XI11_3/net20_4_ XI11_3/preck XI11_3/net21_4_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_11/MP1 XI11_3/net20_4_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_11/MP0 XI11_3/net21_4_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_10/MP2 XI11_3/net20_5_ XI11_3/preck XI11_3/net21_5_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_10/MP1 XI11_3/net20_5_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_10/MP0 XI11_3/net21_5_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_9/MP2 XI11_3/net20_6_ XI11_3/preck XI11_3/net21_6_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_9/MP1 XI11_3/net20_6_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_9/MP0 XI11_3/net21_6_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_8/MP2 XI11_3/net20_7_ XI11_3/preck XI11_3/net21_7_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_8/MP1 XI11_3/net20_7_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_8/MP0 XI11_3/net21_7_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_7/MP2 XI11_3/net20_8_ XI11_3/preck XI11_3/net21_8_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_7/MP1 XI11_3/net20_8_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_7/MP0 XI11_3/net21_8_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_6/MP2 XI11_3/net20_9_ XI11_3/preck XI11_3/net21_9_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_6/MP1 XI11_3/net20_9_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_6/MP0 XI11_3/net21_9_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_5/MP2 XI11_3/net20_10_ XI11_3/preck XI11_3/net21_10_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_5/MP1 XI11_3/net20_10_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_5/MP0 XI11_3/net21_10_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_4/MP2 XI11_3/net20_11_ XI11_3/preck XI11_3/net21_11_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_4/MP1 XI11_3/net20_11_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_4/MP0 XI11_3/net21_11_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_3/MP2 XI11_3/net20_12_ XI11_3/preck XI11_3/net21_12_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_3/MP1 XI11_3/net20_12_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_3/MP0 XI11_3/net21_12_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_2/MP2 XI11_3/net20_13_ XI11_3/preck XI11_3/net21_13_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_2/MP1 XI11_3/net20_13_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_2/MP0 XI11_3/net21_13_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_1/MP2 XI11_3/net20_14_ XI11_3/preck XI11_3/net21_14_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_1/MP1 XI11_3/net20_14_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_1/MP0 XI11_3/net21_14_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_0/MP2 XI11_3/net20_15_ XI11_3/preck XI11_3/net21_15_ vdd MP l=1.8e-07 w=5e-07 $[p18ll] 
XI11_3/XI1_0/MP1 XI11_3/net20_15_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI1_0/MP0 XI11_3/net21_15_ XI11_3/preck vdd vdd MP l=1.8e-07 w=2e-06 $[p18ll] 
XI11_3/XI0/MN0_15 gnd gnd XI11_3/net21_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_14 gnd gnd XI11_3/net21_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_13 gnd gnd XI11_3/net21_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_12 gnd gnd XI11_3/net21_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_11 gnd gnd XI11_3/net21_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_10 gnd gnd XI11_3/net21_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_9 gnd gnd XI11_3/net21_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_8 gnd gnd XI11_3/net21_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_7 gnd gnd XI11_3/net21_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_6 gnd gnd XI11_3/net21_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_5 gnd gnd XI11_3/net21_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_4 gnd gnd XI11_3/net21_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_3 gnd gnd XI11_3/net21_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_2 gnd gnd XI11_3/net21_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_1 gnd gnd XI11_3/net21_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN0_0 gnd gnd XI11_3/net21_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_15 gnd gnd XI11_3/net20_0_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_14 gnd gnd XI11_3/net20_1_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_13 gnd gnd XI11_3/net20_2_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_12 gnd gnd XI11_3/net20_3_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_11 gnd gnd XI11_3/net20_4_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_10 gnd gnd XI11_3/net20_5_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_9 gnd gnd XI11_3/net20_6_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_8 gnd gnd XI11_3/net20_7_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_7 gnd gnd XI11_3/net20_8_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_6 gnd gnd XI11_3/net20_9_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_5 gnd gnd XI11_3/net20_10_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_4 gnd gnd XI11_3/net20_11_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_3 gnd gnd XI11_3/net20_12_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_2 gnd gnd XI11_3/net20_13_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_1 gnd gnd XI11_3/net20_14_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/MN1_0 gnd gnd XI11_3/net20_15_ gnd MN l=2.2e-07 w=4.8e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_15 XI11_3/net21_0_ xsel_63_ XI11_3/XI0/XI0_63/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_14 XI11_3/net21_1_ xsel_63_ XI11_3/XI0/XI0_63/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_13 XI11_3/net21_2_ xsel_63_ XI11_3/XI0/XI0_63/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_12 XI11_3/net21_3_ xsel_63_ XI11_3/XI0/XI0_63/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_11 XI11_3/net21_4_ xsel_63_ XI11_3/XI0/XI0_63/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_10 XI11_3/net21_5_ xsel_63_ XI11_3/XI0/XI0_63/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_9 XI11_3/net21_6_ xsel_63_ XI11_3/XI0/XI0_63/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_8 XI11_3/net21_7_ xsel_63_ XI11_3/XI0/XI0_63/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_7 XI11_3/net21_8_ xsel_63_ XI11_3/XI0/XI0_63/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_6 XI11_3/net21_9_ xsel_63_ XI11_3/XI0/XI0_63/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_5 XI11_3/net21_10_ xsel_63_ XI11_3/XI0/XI0_63/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_4 XI11_3/net21_11_ xsel_63_ XI11_3/XI0/XI0_63/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_3 XI11_3/net21_12_ xsel_63_ XI11_3/XI0/XI0_63/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_2 XI11_3/net21_13_ xsel_63_ XI11_3/XI0/XI0_63/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_1 XI11_3/net21_14_ xsel_63_ XI11_3/XI0/XI0_63/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN0_0 XI11_3/net21_15_ xsel_63_ XI11_3/XI0/XI0_63/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_15 XI11_3/XI0/XI0_63/d__15_ xsel_63_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_14 XI11_3/XI0/XI0_63/d__14_ xsel_63_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_13 XI11_3/XI0/XI0_63/d__13_ xsel_63_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_12 XI11_3/XI0/XI0_63/d__12_ xsel_63_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_11 XI11_3/XI0/XI0_63/d__11_ xsel_63_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_10 XI11_3/XI0/XI0_63/d__10_ xsel_63_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_9 XI11_3/XI0/XI0_63/d__9_ xsel_63_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_8 XI11_3/XI0/XI0_63/d__8_ xsel_63_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_7 XI11_3/XI0/XI0_63/d__7_ xsel_63_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_6 XI11_3/XI0/XI0_63/d__6_ xsel_63_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_5 XI11_3/XI0/XI0_63/d__5_ xsel_63_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_4 XI11_3/XI0/XI0_63/d__4_ xsel_63_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_3 XI11_3/XI0/XI0_63/d__3_ xsel_63_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_2 XI11_3/XI0/XI0_63/d__2_ xsel_63_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_1 XI11_3/XI0/XI0_63/d__1_ xsel_63_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_63/MN1_0 XI11_3/XI0/XI0_63/d__0_ xsel_63_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_15 XI11_3/net21_0_ xsel_62_ XI11_3/XI0/XI0_62/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_14 XI11_3/net21_1_ xsel_62_ XI11_3/XI0/XI0_62/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_13 XI11_3/net21_2_ xsel_62_ XI11_3/XI0/XI0_62/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_12 XI11_3/net21_3_ xsel_62_ XI11_3/XI0/XI0_62/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_11 XI11_3/net21_4_ xsel_62_ XI11_3/XI0/XI0_62/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_10 XI11_3/net21_5_ xsel_62_ XI11_3/XI0/XI0_62/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_9 XI11_3/net21_6_ xsel_62_ XI11_3/XI0/XI0_62/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_8 XI11_3/net21_7_ xsel_62_ XI11_3/XI0/XI0_62/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_7 XI11_3/net21_8_ xsel_62_ XI11_3/XI0/XI0_62/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_6 XI11_3/net21_9_ xsel_62_ XI11_3/XI0/XI0_62/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_5 XI11_3/net21_10_ xsel_62_ XI11_3/XI0/XI0_62/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_4 XI11_3/net21_11_ xsel_62_ XI11_3/XI0/XI0_62/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_3 XI11_3/net21_12_ xsel_62_ XI11_3/XI0/XI0_62/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_2 XI11_3/net21_13_ xsel_62_ XI11_3/XI0/XI0_62/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_1 XI11_3/net21_14_ xsel_62_ XI11_3/XI0/XI0_62/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN0_0 XI11_3/net21_15_ xsel_62_ XI11_3/XI0/XI0_62/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_15 XI11_3/XI0/XI0_62/d__15_ xsel_62_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_14 XI11_3/XI0/XI0_62/d__14_ xsel_62_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_13 XI11_3/XI0/XI0_62/d__13_ xsel_62_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_12 XI11_3/XI0/XI0_62/d__12_ xsel_62_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_11 XI11_3/XI0/XI0_62/d__11_ xsel_62_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_10 XI11_3/XI0/XI0_62/d__10_ xsel_62_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_9 XI11_3/XI0/XI0_62/d__9_ xsel_62_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_8 XI11_3/XI0/XI0_62/d__8_ xsel_62_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_7 XI11_3/XI0/XI0_62/d__7_ xsel_62_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_6 XI11_3/XI0/XI0_62/d__6_ xsel_62_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_5 XI11_3/XI0/XI0_62/d__5_ xsel_62_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_4 XI11_3/XI0/XI0_62/d__4_ xsel_62_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_3 XI11_3/XI0/XI0_62/d__3_ xsel_62_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_2 XI11_3/XI0/XI0_62/d__2_ xsel_62_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_1 XI11_3/XI0/XI0_62/d__1_ xsel_62_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_62/MN1_0 XI11_3/XI0/XI0_62/d__0_ xsel_62_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_15 XI11_3/net21_0_ xsel_61_ XI11_3/XI0/XI0_61/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_14 XI11_3/net21_1_ xsel_61_ XI11_3/XI0/XI0_61/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_13 XI11_3/net21_2_ xsel_61_ XI11_3/XI0/XI0_61/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_12 XI11_3/net21_3_ xsel_61_ XI11_3/XI0/XI0_61/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_11 XI11_3/net21_4_ xsel_61_ XI11_3/XI0/XI0_61/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_10 XI11_3/net21_5_ xsel_61_ XI11_3/XI0/XI0_61/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_9 XI11_3/net21_6_ xsel_61_ XI11_3/XI0/XI0_61/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_8 XI11_3/net21_7_ xsel_61_ XI11_3/XI0/XI0_61/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_7 XI11_3/net21_8_ xsel_61_ XI11_3/XI0/XI0_61/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_6 XI11_3/net21_9_ xsel_61_ XI11_3/XI0/XI0_61/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_5 XI11_3/net21_10_ xsel_61_ XI11_3/XI0/XI0_61/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_4 XI11_3/net21_11_ xsel_61_ XI11_3/XI0/XI0_61/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_3 XI11_3/net21_12_ xsel_61_ XI11_3/XI0/XI0_61/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_2 XI11_3/net21_13_ xsel_61_ XI11_3/XI0/XI0_61/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_1 XI11_3/net21_14_ xsel_61_ XI11_3/XI0/XI0_61/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN0_0 XI11_3/net21_15_ xsel_61_ XI11_3/XI0/XI0_61/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_15 XI11_3/XI0/XI0_61/d__15_ xsel_61_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_14 XI11_3/XI0/XI0_61/d__14_ xsel_61_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_13 XI11_3/XI0/XI0_61/d__13_ xsel_61_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_12 XI11_3/XI0/XI0_61/d__12_ xsel_61_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_11 XI11_3/XI0/XI0_61/d__11_ xsel_61_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_10 XI11_3/XI0/XI0_61/d__10_ xsel_61_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_9 XI11_3/XI0/XI0_61/d__9_ xsel_61_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_8 XI11_3/XI0/XI0_61/d__8_ xsel_61_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_7 XI11_3/XI0/XI0_61/d__7_ xsel_61_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_6 XI11_3/XI0/XI0_61/d__6_ xsel_61_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_5 XI11_3/XI0/XI0_61/d__5_ xsel_61_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_4 XI11_3/XI0/XI0_61/d__4_ xsel_61_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_3 XI11_3/XI0/XI0_61/d__3_ xsel_61_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_2 XI11_3/XI0/XI0_61/d__2_ xsel_61_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_1 XI11_3/XI0/XI0_61/d__1_ xsel_61_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_61/MN1_0 XI11_3/XI0/XI0_61/d__0_ xsel_61_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_15 XI11_3/net21_0_ xsel_60_ XI11_3/XI0/XI0_60/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_14 XI11_3/net21_1_ xsel_60_ XI11_3/XI0/XI0_60/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_13 XI11_3/net21_2_ xsel_60_ XI11_3/XI0/XI0_60/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_12 XI11_3/net21_3_ xsel_60_ XI11_3/XI0/XI0_60/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_11 XI11_3/net21_4_ xsel_60_ XI11_3/XI0/XI0_60/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_10 XI11_3/net21_5_ xsel_60_ XI11_3/XI0/XI0_60/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_9 XI11_3/net21_6_ xsel_60_ XI11_3/XI0/XI0_60/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_8 XI11_3/net21_7_ xsel_60_ XI11_3/XI0/XI0_60/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_7 XI11_3/net21_8_ xsel_60_ XI11_3/XI0/XI0_60/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_6 XI11_3/net21_9_ xsel_60_ XI11_3/XI0/XI0_60/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_5 XI11_3/net21_10_ xsel_60_ XI11_3/XI0/XI0_60/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_4 XI11_3/net21_11_ xsel_60_ XI11_3/XI0/XI0_60/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_3 XI11_3/net21_12_ xsel_60_ XI11_3/XI0/XI0_60/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_2 XI11_3/net21_13_ xsel_60_ XI11_3/XI0/XI0_60/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_1 XI11_3/net21_14_ xsel_60_ XI11_3/XI0/XI0_60/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN0_0 XI11_3/net21_15_ xsel_60_ XI11_3/XI0/XI0_60/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_15 XI11_3/XI0/XI0_60/d__15_ xsel_60_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_14 XI11_3/XI0/XI0_60/d__14_ xsel_60_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_13 XI11_3/XI0/XI0_60/d__13_ xsel_60_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_12 XI11_3/XI0/XI0_60/d__12_ xsel_60_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_11 XI11_3/XI0/XI0_60/d__11_ xsel_60_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_10 XI11_3/XI0/XI0_60/d__10_ xsel_60_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_9 XI11_3/XI0/XI0_60/d__9_ xsel_60_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_8 XI11_3/XI0/XI0_60/d__8_ xsel_60_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_7 XI11_3/XI0/XI0_60/d__7_ xsel_60_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_6 XI11_3/XI0/XI0_60/d__6_ xsel_60_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_5 XI11_3/XI0/XI0_60/d__5_ xsel_60_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_4 XI11_3/XI0/XI0_60/d__4_ xsel_60_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_3 XI11_3/XI0/XI0_60/d__3_ xsel_60_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_2 XI11_3/XI0/XI0_60/d__2_ xsel_60_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_1 XI11_3/XI0/XI0_60/d__1_ xsel_60_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_60/MN1_0 XI11_3/XI0/XI0_60/d__0_ xsel_60_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_15 XI11_3/net21_0_ xsel_59_ XI11_3/XI0/XI0_59/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_14 XI11_3/net21_1_ xsel_59_ XI11_3/XI0/XI0_59/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_13 XI11_3/net21_2_ xsel_59_ XI11_3/XI0/XI0_59/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_12 XI11_3/net21_3_ xsel_59_ XI11_3/XI0/XI0_59/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_11 XI11_3/net21_4_ xsel_59_ XI11_3/XI0/XI0_59/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_10 XI11_3/net21_5_ xsel_59_ XI11_3/XI0/XI0_59/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_9 XI11_3/net21_6_ xsel_59_ XI11_3/XI0/XI0_59/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_8 XI11_3/net21_7_ xsel_59_ XI11_3/XI0/XI0_59/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_7 XI11_3/net21_8_ xsel_59_ XI11_3/XI0/XI0_59/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_6 XI11_3/net21_9_ xsel_59_ XI11_3/XI0/XI0_59/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_5 XI11_3/net21_10_ xsel_59_ XI11_3/XI0/XI0_59/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_4 XI11_3/net21_11_ xsel_59_ XI11_3/XI0/XI0_59/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_3 XI11_3/net21_12_ xsel_59_ XI11_3/XI0/XI0_59/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_2 XI11_3/net21_13_ xsel_59_ XI11_3/XI0/XI0_59/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_1 XI11_3/net21_14_ xsel_59_ XI11_3/XI0/XI0_59/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN0_0 XI11_3/net21_15_ xsel_59_ XI11_3/XI0/XI0_59/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_15 XI11_3/XI0/XI0_59/d__15_ xsel_59_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_14 XI11_3/XI0/XI0_59/d__14_ xsel_59_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_13 XI11_3/XI0/XI0_59/d__13_ xsel_59_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_12 XI11_3/XI0/XI0_59/d__12_ xsel_59_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_11 XI11_3/XI0/XI0_59/d__11_ xsel_59_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_10 XI11_3/XI0/XI0_59/d__10_ xsel_59_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_9 XI11_3/XI0/XI0_59/d__9_ xsel_59_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_8 XI11_3/XI0/XI0_59/d__8_ xsel_59_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_7 XI11_3/XI0/XI0_59/d__7_ xsel_59_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_6 XI11_3/XI0/XI0_59/d__6_ xsel_59_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_5 XI11_3/XI0/XI0_59/d__5_ xsel_59_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_4 XI11_3/XI0/XI0_59/d__4_ xsel_59_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_3 XI11_3/XI0/XI0_59/d__3_ xsel_59_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_2 XI11_3/XI0/XI0_59/d__2_ xsel_59_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_1 XI11_3/XI0/XI0_59/d__1_ xsel_59_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_59/MN1_0 XI11_3/XI0/XI0_59/d__0_ xsel_59_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_15 XI11_3/net21_0_ xsel_58_ XI11_3/XI0/XI0_58/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_14 XI11_3/net21_1_ xsel_58_ XI11_3/XI0/XI0_58/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_13 XI11_3/net21_2_ xsel_58_ XI11_3/XI0/XI0_58/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_12 XI11_3/net21_3_ xsel_58_ XI11_3/XI0/XI0_58/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_11 XI11_3/net21_4_ xsel_58_ XI11_3/XI0/XI0_58/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_10 XI11_3/net21_5_ xsel_58_ XI11_3/XI0/XI0_58/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_9 XI11_3/net21_6_ xsel_58_ XI11_3/XI0/XI0_58/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_8 XI11_3/net21_7_ xsel_58_ XI11_3/XI0/XI0_58/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_7 XI11_3/net21_8_ xsel_58_ XI11_3/XI0/XI0_58/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_6 XI11_3/net21_9_ xsel_58_ XI11_3/XI0/XI0_58/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_5 XI11_3/net21_10_ xsel_58_ XI11_3/XI0/XI0_58/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_4 XI11_3/net21_11_ xsel_58_ XI11_3/XI0/XI0_58/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_3 XI11_3/net21_12_ xsel_58_ XI11_3/XI0/XI0_58/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_2 XI11_3/net21_13_ xsel_58_ XI11_3/XI0/XI0_58/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_1 XI11_3/net21_14_ xsel_58_ XI11_3/XI0/XI0_58/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN0_0 XI11_3/net21_15_ xsel_58_ XI11_3/XI0/XI0_58/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_15 XI11_3/XI0/XI0_58/d__15_ xsel_58_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_14 XI11_3/XI0/XI0_58/d__14_ xsel_58_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_13 XI11_3/XI0/XI0_58/d__13_ xsel_58_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_12 XI11_3/XI0/XI0_58/d__12_ xsel_58_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_11 XI11_3/XI0/XI0_58/d__11_ xsel_58_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_10 XI11_3/XI0/XI0_58/d__10_ xsel_58_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_9 XI11_3/XI0/XI0_58/d__9_ xsel_58_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_8 XI11_3/XI0/XI0_58/d__8_ xsel_58_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_7 XI11_3/XI0/XI0_58/d__7_ xsel_58_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_6 XI11_3/XI0/XI0_58/d__6_ xsel_58_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_5 XI11_3/XI0/XI0_58/d__5_ xsel_58_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_4 XI11_3/XI0/XI0_58/d__4_ xsel_58_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_3 XI11_3/XI0/XI0_58/d__3_ xsel_58_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_2 XI11_3/XI0/XI0_58/d__2_ xsel_58_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_1 XI11_3/XI0/XI0_58/d__1_ xsel_58_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_58/MN1_0 XI11_3/XI0/XI0_58/d__0_ xsel_58_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_15 XI11_3/net21_0_ xsel_57_ XI11_3/XI0/XI0_57/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_14 XI11_3/net21_1_ xsel_57_ XI11_3/XI0/XI0_57/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_13 XI11_3/net21_2_ xsel_57_ XI11_3/XI0/XI0_57/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_12 XI11_3/net21_3_ xsel_57_ XI11_3/XI0/XI0_57/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_11 XI11_3/net21_4_ xsel_57_ XI11_3/XI0/XI0_57/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_10 XI11_3/net21_5_ xsel_57_ XI11_3/XI0/XI0_57/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_9 XI11_3/net21_6_ xsel_57_ XI11_3/XI0/XI0_57/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_8 XI11_3/net21_7_ xsel_57_ XI11_3/XI0/XI0_57/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_7 XI11_3/net21_8_ xsel_57_ XI11_3/XI0/XI0_57/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_6 XI11_3/net21_9_ xsel_57_ XI11_3/XI0/XI0_57/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_5 XI11_3/net21_10_ xsel_57_ XI11_3/XI0/XI0_57/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_4 XI11_3/net21_11_ xsel_57_ XI11_3/XI0/XI0_57/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_3 XI11_3/net21_12_ xsel_57_ XI11_3/XI0/XI0_57/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_2 XI11_3/net21_13_ xsel_57_ XI11_3/XI0/XI0_57/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_1 XI11_3/net21_14_ xsel_57_ XI11_3/XI0/XI0_57/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN0_0 XI11_3/net21_15_ xsel_57_ XI11_3/XI0/XI0_57/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_15 XI11_3/XI0/XI0_57/d__15_ xsel_57_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_14 XI11_3/XI0/XI0_57/d__14_ xsel_57_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_13 XI11_3/XI0/XI0_57/d__13_ xsel_57_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_12 XI11_3/XI0/XI0_57/d__12_ xsel_57_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_11 XI11_3/XI0/XI0_57/d__11_ xsel_57_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_10 XI11_3/XI0/XI0_57/d__10_ xsel_57_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_9 XI11_3/XI0/XI0_57/d__9_ xsel_57_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_8 XI11_3/XI0/XI0_57/d__8_ xsel_57_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_7 XI11_3/XI0/XI0_57/d__7_ xsel_57_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_6 XI11_3/XI0/XI0_57/d__6_ xsel_57_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_5 XI11_3/XI0/XI0_57/d__5_ xsel_57_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_4 XI11_3/XI0/XI0_57/d__4_ xsel_57_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_3 XI11_3/XI0/XI0_57/d__3_ xsel_57_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_2 XI11_3/XI0/XI0_57/d__2_ xsel_57_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_1 XI11_3/XI0/XI0_57/d__1_ xsel_57_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_57/MN1_0 XI11_3/XI0/XI0_57/d__0_ xsel_57_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_15 XI11_3/net21_0_ xsel_56_ XI11_3/XI0/XI0_56/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_14 XI11_3/net21_1_ xsel_56_ XI11_3/XI0/XI0_56/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_13 XI11_3/net21_2_ xsel_56_ XI11_3/XI0/XI0_56/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_12 XI11_3/net21_3_ xsel_56_ XI11_3/XI0/XI0_56/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_11 XI11_3/net21_4_ xsel_56_ XI11_3/XI0/XI0_56/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_10 XI11_3/net21_5_ xsel_56_ XI11_3/XI0/XI0_56/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_9 XI11_3/net21_6_ xsel_56_ XI11_3/XI0/XI0_56/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_8 XI11_3/net21_7_ xsel_56_ XI11_3/XI0/XI0_56/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_7 XI11_3/net21_8_ xsel_56_ XI11_3/XI0/XI0_56/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_6 XI11_3/net21_9_ xsel_56_ XI11_3/XI0/XI0_56/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_5 XI11_3/net21_10_ xsel_56_ XI11_3/XI0/XI0_56/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_4 XI11_3/net21_11_ xsel_56_ XI11_3/XI0/XI0_56/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_3 XI11_3/net21_12_ xsel_56_ XI11_3/XI0/XI0_56/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_2 XI11_3/net21_13_ xsel_56_ XI11_3/XI0/XI0_56/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_1 XI11_3/net21_14_ xsel_56_ XI11_3/XI0/XI0_56/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN0_0 XI11_3/net21_15_ xsel_56_ XI11_3/XI0/XI0_56/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_15 XI11_3/XI0/XI0_56/d__15_ xsel_56_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_14 XI11_3/XI0/XI0_56/d__14_ xsel_56_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_13 XI11_3/XI0/XI0_56/d__13_ xsel_56_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_12 XI11_3/XI0/XI0_56/d__12_ xsel_56_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_11 XI11_3/XI0/XI0_56/d__11_ xsel_56_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_10 XI11_3/XI0/XI0_56/d__10_ xsel_56_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_9 XI11_3/XI0/XI0_56/d__9_ xsel_56_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_8 XI11_3/XI0/XI0_56/d__8_ xsel_56_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_7 XI11_3/XI0/XI0_56/d__7_ xsel_56_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_6 XI11_3/XI0/XI0_56/d__6_ xsel_56_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_5 XI11_3/XI0/XI0_56/d__5_ xsel_56_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_4 XI11_3/XI0/XI0_56/d__4_ xsel_56_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_3 XI11_3/XI0/XI0_56/d__3_ xsel_56_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_2 XI11_3/XI0/XI0_56/d__2_ xsel_56_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_1 XI11_3/XI0/XI0_56/d__1_ xsel_56_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_56/MN1_0 XI11_3/XI0/XI0_56/d__0_ xsel_56_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_15 XI11_3/net21_0_ xsel_55_ XI11_3/XI0/XI0_55/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_14 XI11_3/net21_1_ xsel_55_ XI11_3/XI0/XI0_55/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_13 XI11_3/net21_2_ xsel_55_ XI11_3/XI0/XI0_55/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_12 XI11_3/net21_3_ xsel_55_ XI11_3/XI0/XI0_55/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_11 XI11_3/net21_4_ xsel_55_ XI11_3/XI0/XI0_55/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_10 XI11_3/net21_5_ xsel_55_ XI11_3/XI0/XI0_55/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_9 XI11_3/net21_6_ xsel_55_ XI11_3/XI0/XI0_55/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_8 XI11_3/net21_7_ xsel_55_ XI11_3/XI0/XI0_55/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_7 XI11_3/net21_8_ xsel_55_ XI11_3/XI0/XI0_55/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_6 XI11_3/net21_9_ xsel_55_ XI11_3/XI0/XI0_55/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_5 XI11_3/net21_10_ xsel_55_ XI11_3/XI0/XI0_55/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_4 XI11_3/net21_11_ xsel_55_ XI11_3/XI0/XI0_55/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_3 XI11_3/net21_12_ xsel_55_ XI11_3/XI0/XI0_55/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_2 XI11_3/net21_13_ xsel_55_ XI11_3/XI0/XI0_55/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_1 XI11_3/net21_14_ xsel_55_ XI11_3/XI0/XI0_55/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN0_0 XI11_3/net21_15_ xsel_55_ XI11_3/XI0/XI0_55/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_15 XI11_3/XI0/XI0_55/d__15_ xsel_55_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_14 XI11_3/XI0/XI0_55/d__14_ xsel_55_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_13 XI11_3/XI0/XI0_55/d__13_ xsel_55_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_12 XI11_3/XI0/XI0_55/d__12_ xsel_55_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_11 XI11_3/XI0/XI0_55/d__11_ xsel_55_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_10 XI11_3/XI0/XI0_55/d__10_ xsel_55_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_9 XI11_3/XI0/XI0_55/d__9_ xsel_55_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_8 XI11_3/XI0/XI0_55/d__8_ xsel_55_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_7 XI11_3/XI0/XI0_55/d__7_ xsel_55_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_6 XI11_3/XI0/XI0_55/d__6_ xsel_55_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_5 XI11_3/XI0/XI0_55/d__5_ xsel_55_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_4 XI11_3/XI0/XI0_55/d__4_ xsel_55_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_3 XI11_3/XI0/XI0_55/d__3_ xsel_55_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_2 XI11_3/XI0/XI0_55/d__2_ xsel_55_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_1 XI11_3/XI0/XI0_55/d__1_ xsel_55_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_55/MN1_0 XI11_3/XI0/XI0_55/d__0_ xsel_55_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_15 XI11_3/net21_0_ xsel_54_ XI11_3/XI0/XI0_54/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_14 XI11_3/net21_1_ xsel_54_ XI11_3/XI0/XI0_54/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_13 XI11_3/net21_2_ xsel_54_ XI11_3/XI0/XI0_54/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_12 XI11_3/net21_3_ xsel_54_ XI11_3/XI0/XI0_54/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_11 XI11_3/net21_4_ xsel_54_ XI11_3/XI0/XI0_54/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_10 XI11_3/net21_5_ xsel_54_ XI11_3/XI0/XI0_54/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_9 XI11_3/net21_6_ xsel_54_ XI11_3/XI0/XI0_54/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_8 XI11_3/net21_7_ xsel_54_ XI11_3/XI0/XI0_54/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_7 XI11_3/net21_8_ xsel_54_ XI11_3/XI0/XI0_54/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_6 XI11_3/net21_9_ xsel_54_ XI11_3/XI0/XI0_54/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_5 XI11_3/net21_10_ xsel_54_ XI11_3/XI0/XI0_54/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_4 XI11_3/net21_11_ xsel_54_ XI11_3/XI0/XI0_54/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_3 XI11_3/net21_12_ xsel_54_ XI11_3/XI0/XI0_54/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_2 XI11_3/net21_13_ xsel_54_ XI11_3/XI0/XI0_54/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_1 XI11_3/net21_14_ xsel_54_ XI11_3/XI0/XI0_54/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN0_0 XI11_3/net21_15_ xsel_54_ XI11_3/XI0/XI0_54/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_15 XI11_3/XI0/XI0_54/d__15_ xsel_54_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_14 XI11_3/XI0/XI0_54/d__14_ xsel_54_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_13 XI11_3/XI0/XI0_54/d__13_ xsel_54_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_12 XI11_3/XI0/XI0_54/d__12_ xsel_54_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_11 XI11_3/XI0/XI0_54/d__11_ xsel_54_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_10 XI11_3/XI0/XI0_54/d__10_ xsel_54_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_9 XI11_3/XI0/XI0_54/d__9_ xsel_54_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_8 XI11_3/XI0/XI0_54/d__8_ xsel_54_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_7 XI11_3/XI0/XI0_54/d__7_ xsel_54_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_6 XI11_3/XI0/XI0_54/d__6_ xsel_54_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_5 XI11_3/XI0/XI0_54/d__5_ xsel_54_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_4 XI11_3/XI0/XI0_54/d__4_ xsel_54_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_3 XI11_3/XI0/XI0_54/d__3_ xsel_54_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_2 XI11_3/XI0/XI0_54/d__2_ xsel_54_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_1 XI11_3/XI0/XI0_54/d__1_ xsel_54_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_54/MN1_0 XI11_3/XI0/XI0_54/d__0_ xsel_54_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_15 XI11_3/net21_0_ xsel_53_ XI11_3/XI0/XI0_53/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_14 XI11_3/net21_1_ xsel_53_ XI11_3/XI0/XI0_53/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_13 XI11_3/net21_2_ xsel_53_ XI11_3/XI0/XI0_53/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_12 XI11_3/net21_3_ xsel_53_ XI11_3/XI0/XI0_53/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_11 XI11_3/net21_4_ xsel_53_ XI11_3/XI0/XI0_53/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_10 XI11_3/net21_5_ xsel_53_ XI11_3/XI0/XI0_53/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_9 XI11_3/net21_6_ xsel_53_ XI11_3/XI0/XI0_53/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_8 XI11_3/net21_7_ xsel_53_ XI11_3/XI0/XI0_53/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_7 XI11_3/net21_8_ xsel_53_ XI11_3/XI0/XI0_53/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_6 XI11_3/net21_9_ xsel_53_ XI11_3/XI0/XI0_53/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_5 XI11_3/net21_10_ xsel_53_ XI11_3/XI0/XI0_53/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_4 XI11_3/net21_11_ xsel_53_ XI11_3/XI0/XI0_53/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_3 XI11_3/net21_12_ xsel_53_ XI11_3/XI0/XI0_53/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_2 XI11_3/net21_13_ xsel_53_ XI11_3/XI0/XI0_53/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_1 XI11_3/net21_14_ xsel_53_ XI11_3/XI0/XI0_53/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN0_0 XI11_3/net21_15_ xsel_53_ XI11_3/XI0/XI0_53/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_15 XI11_3/XI0/XI0_53/d__15_ xsel_53_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_14 XI11_3/XI0/XI0_53/d__14_ xsel_53_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_13 XI11_3/XI0/XI0_53/d__13_ xsel_53_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_12 XI11_3/XI0/XI0_53/d__12_ xsel_53_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_11 XI11_3/XI0/XI0_53/d__11_ xsel_53_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_10 XI11_3/XI0/XI0_53/d__10_ xsel_53_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_9 XI11_3/XI0/XI0_53/d__9_ xsel_53_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_8 XI11_3/XI0/XI0_53/d__8_ xsel_53_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_7 XI11_3/XI0/XI0_53/d__7_ xsel_53_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_6 XI11_3/XI0/XI0_53/d__6_ xsel_53_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_5 XI11_3/XI0/XI0_53/d__5_ xsel_53_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_4 XI11_3/XI0/XI0_53/d__4_ xsel_53_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_3 XI11_3/XI0/XI0_53/d__3_ xsel_53_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_2 XI11_3/XI0/XI0_53/d__2_ xsel_53_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_1 XI11_3/XI0/XI0_53/d__1_ xsel_53_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_53/MN1_0 XI11_3/XI0/XI0_53/d__0_ xsel_53_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_15 XI11_3/net21_0_ xsel_52_ XI11_3/XI0/XI0_52/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_14 XI11_3/net21_1_ xsel_52_ XI11_3/XI0/XI0_52/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_13 XI11_3/net21_2_ xsel_52_ XI11_3/XI0/XI0_52/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_12 XI11_3/net21_3_ xsel_52_ XI11_3/XI0/XI0_52/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_11 XI11_3/net21_4_ xsel_52_ XI11_3/XI0/XI0_52/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_10 XI11_3/net21_5_ xsel_52_ XI11_3/XI0/XI0_52/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_9 XI11_3/net21_6_ xsel_52_ XI11_3/XI0/XI0_52/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_8 XI11_3/net21_7_ xsel_52_ XI11_3/XI0/XI0_52/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_7 XI11_3/net21_8_ xsel_52_ XI11_3/XI0/XI0_52/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_6 XI11_3/net21_9_ xsel_52_ XI11_3/XI0/XI0_52/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_5 XI11_3/net21_10_ xsel_52_ XI11_3/XI0/XI0_52/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_4 XI11_3/net21_11_ xsel_52_ XI11_3/XI0/XI0_52/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_3 XI11_3/net21_12_ xsel_52_ XI11_3/XI0/XI0_52/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_2 XI11_3/net21_13_ xsel_52_ XI11_3/XI0/XI0_52/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_1 XI11_3/net21_14_ xsel_52_ XI11_3/XI0/XI0_52/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN0_0 XI11_3/net21_15_ xsel_52_ XI11_3/XI0/XI0_52/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_15 XI11_3/XI0/XI0_52/d__15_ xsel_52_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_14 XI11_3/XI0/XI0_52/d__14_ xsel_52_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_13 XI11_3/XI0/XI0_52/d__13_ xsel_52_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_12 XI11_3/XI0/XI0_52/d__12_ xsel_52_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_11 XI11_3/XI0/XI0_52/d__11_ xsel_52_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_10 XI11_3/XI0/XI0_52/d__10_ xsel_52_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_9 XI11_3/XI0/XI0_52/d__9_ xsel_52_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_8 XI11_3/XI0/XI0_52/d__8_ xsel_52_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_7 XI11_3/XI0/XI0_52/d__7_ xsel_52_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_6 XI11_3/XI0/XI0_52/d__6_ xsel_52_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_5 XI11_3/XI0/XI0_52/d__5_ xsel_52_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_4 XI11_3/XI0/XI0_52/d__4_ xsel_52_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_3 XI11_3/XI0/XI0_52/d__3_ xsel_52_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_2 XI11_3/XI0/XI0_52/d__2_ xsel_52_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_1 XI11_3/XI0/XI0_52/d__1_ xsel_52_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_52/MN1_0 XI11_3/XI0/XI0_52/d__0_ xsel_52_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_15 XI11_3/net21_0_ xsel_51_ XI11_3/XI0/XI0_51/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_14 XI11_3/net21_1_ xsel_51_ XI11_3/XI0/XI0_51/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_13 XI11_3/net21_2_ xsel_51_ XI11_3/XI0/XI0_51/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_12 XI11_3/net21_3_ xsel_51_ XI11_3/XI0/XI0_51/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_11 XI11_3/net21_4_ xsel_51_ XI11_3/XI0/XI0_51/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_10 XI11_3/net21_5_ xsel_51_ XI11_3/XI0/XI0_51/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_9 XI11_3/net21_6_ xsel_51_ XI11_3/XI0/XI0_51/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_8 XI11_3/net21_7_ xsel_51_ XI11_3/XI0/XI0_51/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_7 XI11_3/net21_8_ xsel_51_ XI11_3/XI0/XI0_51/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_6 XI11_3/net21_9_ xsel_51_ XI11_3/XI0/XI0_51/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_5 XI11_3/net21_10_ xsel_51_ XI11_3/XI0/XI0_51/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_4 XI11_3/net21_11_ xsel_51_ XI11_3/XI0/XI0_51/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_3 XI11_3/net21_12_ xsel_51_ XI11_3/XI0/XI0_51/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_2 XI11_3/net21_13_ xsel_51_ XI11_3/XI0/XI0_51/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_1 XI11_3/net21_14_ xsel_51_ XI11_3/XI0/XI0_51/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN0_0 XI11_3/net21_15_ xsel_51_ XI11_3/XI0/XI0_51/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_15 XI11_3/XI0/XI0_51/d__15_ xsel_51_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_14 XI11_3/XI0/XI0_51/d__14_ xsel_51_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_13 XI11_3/XI0/XI0_51/d__13_ xsel_51_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_12 XI11_3/XI0/XI0_51/d__12_ xsel_51_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_11 XI11_3/XI0/XI0_51/d__11_ xsel_51_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_10 XI11_3/XI0/XI0_51/d__10_ xsel_51_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_9 XI11_3/XI0/XI0_51/d__9_ xsel_51_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_8 XI11_3/XI0/XI0_51/d__8_ xsel_51_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_7 XI11_3/XI0/XI0_51/d__7_ xsel_51_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_6 XI11_3/XI0/XI0_51/d__6_ xsel_51_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_5 XI11_3/XI0/XI0_51/d__5_ xsel_51_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_4 XI11_3/XI0/XI0_51/d__4_ xsel_51_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_3 XI11_3/XI0/XI0_51/d__3_ xsel_51_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_2 XI11_3/XI0/XI0_51/d__2_ xsel_51_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_1 XI11_3/XI0/XI0_51/d__1_ xsel_51_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_51/MN1_0 XI11_3/XI0/XI0_51/d__0_ xsel_51_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_15 XI11_3/net21_0_ xsel_50_ XI11_3/XI0/XI0_50/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_14 XI11_3/net21_1_ xsel_50_ XI11_3/XI0/XI0_50/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_13 XI11_3/net21_2_ xsel_50_ XI11_3/XI0/XI0_50/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_12 XI11_3/net21_3_ xsel_50_ XI11_3/XI0/XI0_50/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_11 XI11_3/net21_4_ xsel_50_ XI11_3/XI0/XI0_50/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_10 XI11_3/net21_5_ xsel_50_ XI11_3/XI0/XI0_50/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_9 XI11_3/net21_6_ xsel_50_ XI11_3/XI0/XI0_50/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_8 XI11_3/net21_7_ xsel_50_ XI11_3/XI0/XI0_50/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_7 XI11_3/net21_8_ xsel_50_ XI11_3/XI0/XI0_50/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_6 XI11_3/net21_9_ xsel_50_ XI11_3/XI0/XI0_50/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_5 XI11_3/net21_10_ xsel_50_ XI11_3/XI0/XI0_50/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_4 XI11_3/net21_11_ xsel_50_ XI11_3/XI0/XI0_50/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_3 XI11_3/net21_12_ xsel_50_ XI11_3/XI0/XI0_50/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_2 XI11_3/net21_13_ xsel_50_ XI11_3/XI0/XI0_50/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_1 XI11_3/net21_14_ xsel_50_ XI11_3/XI0/XI0_50/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN0_0 XI11_3/net21_15_ xsel_50_ XI11_3/XI0/XI0_50/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_15 XI11_3/XI0/XI0_50/d__15_ xsel_50_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_14 XI11_3/XI0/XI0_50/d__14_ xsel_50_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_13 XI11_3/XI0/XI0_50/d__13_ xsel_50_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_12 XI11_3/XI0/XI0_50/d__12_ xsel_50_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_11 XI11_3/XI0/XI0_50/d__11_ xsel_50_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_10 XI11_3/XI0/XI0_50/d__10_ xsel_50_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_9 XI11_3/XI0/XI0_50/d__9_ xsel_50_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_8 XI11_3/XI0/XI0_50/d__8_ xsel_50_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_7 XI11_3/XI0/XI0_50/d__7_ xsel_50_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_6 XI11_3/XI0/XI0_50/d__6_ xsel_50_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_5 XI11_3/XI0/XI0_50/d__5_ xsel_50_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_4 XI11_3/XI0/XI0_50/d__4_ xsel_50_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_3 XI11_3/XI0/XI0_50/d__3_ xsel_50_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_2 XI11_3/XI0/XI0_50/d__2_ xsel_50_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_1 XI11_3/XI0/XI0_50/d__1_ xsel_50_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_50/MN1_0 XI11_3/XI0/XI0_50/d__0_ xsel_50_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_15 XI11_3/net21_0_ xsel_49_ XI11_3/XI0/XI0_49/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_14 XI11_3/net21_1_ xsel_49_ XI11_3/XI0/XI0_49/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_13 XI11_3/net21_2_ xsel_49_ XI11_3/XI0/XI0_49/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_12 XI11_3/net21_3_ xsel_49_ XI11_3/XI0/XI0_49/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_11 XI11_3/net21_4_ xsel_49_ XI11_3/XI0/XI0_49/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_10 XI11_3/net21_5_ xsel_49_ XI11_3/XI0/XI0_49/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_9 XI11_3/net21_6_ xsel_49_ XI11_3/XI0/XI0_49/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_8 XI11_3/net21_7_ xsel_49_ XI11_3/XI0/XI0_49/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_7 XI11_3/net21_8_ xsel_49_ XI11_3/XI0/XI0_49/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_6 XI11_3/net21_9_ xsel_49_ XI11_3/XI0/XI0_49/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_5 XI11_3/net21_10_ xsel_49_ XI11_3/XI0/XI0_49/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_4 XI11_3/net21_11_ xsel_49_ XI11_3/XI0/XI0_49/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_3 XI11_3/net21_12_ xsel_49_ XI11_3/XI0/XI0_49/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_2 XI11_3/net21_13_ xsel_49_ XI11_3/XI0/XI0_49/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_1 XI11_3/net21_14_ xsel_49_ XI11_3/XI0/XI0_49/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN0_0 XI11_3/net21_15_ xsel_49_ XI11_3/XI0/XI0_49/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_15 XI11_3/XI0/XI0_49/d__15_ xsel_49_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_14 XI11_3/XI0/XI0_49/d__14_ xsel_49_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_13 XI11_3/XI0/XI0_49/d__13_ xsel_49_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_12 XI11_3/XI0/XI0_49/d__12_ xsel_49_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_11 XI11_3/XI0/XI0_49/d__11_ xsel_49_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_10 XI11_3/XI0/XI0_49/d__10_ xsel_49_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_9 XI11_3/XI0/XI0_49/d__9_ xsel_49_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_8 XI11_3/XI0/XI0_49/d__8_ xsel_49_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_7 XI11_3/XI0/XI0_49/d__7_ xsel_49_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_6 XI11_3/XI0/XI0_49/d__6_ xsel_49_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_5 XI11_3/XI0/XI0_49/d__5_ xsel_49_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_4 XI11_3/XI0/XI0_49/d__4_ xsel_49_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_3 XI11_3/XI0/XI0_49/d__3_ xsel_49_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_2 XI11_3/XI0/XI0_49/d__2_ xsel_49_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_1 XI11_3/XI0/XI0_49/d__1_ xsel_49_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_49/MN1_0 XI11_3/XI0/XI0_49/d__0_ xsel_49_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_15 XI11_3/net21_0_ xsel_48_ XI11_3/XI0/XI0_48/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_14 XI11_3/net21_1_ xsel_48_ XI11_3/XI0/XI0_48/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_13 XI11_3/net21_2_ xsel_48_ XI11_3/XI0/XI0_48/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_12 XI11_3/net21_3_ xsel_48_ XI11_3/XI0/XI0_48/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_11 XI11_3/net21_4_ xsel_48_ XI11_3/XI0/XI0_48/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_10 XI11_3/net21_5_ xsel_48_ XI11_3/XI0/XI0_48/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_9 XI11_3/net21_6_ xsel_48_ XI11_3/XI0/XI0_48/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_8 XI11_3/net21_7_ xsel_48_ XI11_3/XI0/XI0_48/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_7 XI11_3/net21_8_ xsel_48_ XI11_3/XI0/XI0_48/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_6 XI11_3/net21_9_ xsel_48_ XI11_3/XI0/XI0_48/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_5 XI11_3/net21_10_ xsel_48_ XI11_3/XI0/XI0_48/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_4 XI11_3/net21_11_ xsel_48_ XI11_3/XI0/XI0_48/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_3 XI11_3/net21_12_ xsel_48_ XI11_3/XI0/XI0_48/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_2 XI11_3/net21_13_ xsel_48_ XI11_3/XI0/XI0_48/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_1 XI11_3/net21_14_ xsel_48_ XI11_3/XI0/XI0_48/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN0_0 XI11_3/net21_15_ xsel_48_ XI11_3/XI0/XI0_48/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_15 XI11_3/XI0/XI0_48/d__15_ xsel_48_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_14 XI11_3/XI0/XI0_48/d__14_ xsel_48_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_13 XI11_3/XI0/XI0_48/d__13_ xsel_48_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_12 XI11_3/XI0/XI0_48/d__12_ xsel_48_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_11 XI11_3/XI0/XI0_48/d__11_ xsel_48_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_10 XI11_3/XI0/XI0_48/d__10_ xsel_48_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_9 XI11_3/XI0/XI0_48/d__9_ xsel_48_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_8 XI11_3/XI0/XI0_48/d__8_ xsel_48_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_7 XI11_3/XI0/XI0_48/d__7_ xsel_48_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_6 XI11_3/XI0/XI0_48/d__6_ xsel_48_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_5 XI11_3/XI0/XI0_48/d__5_ xsel_48_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_4 XI11_3/XI0/XI0_48/d__4_ xsel_48_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_3 XI11_3/XI0/XI0_48/d__3_ xsel_48_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_2 XI11_3/XI0/XI0_48/d__2_ xsel_48_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_1 XI11_3/XI0/XI0_48/d__1_ xsel_48_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_48/MN1_0 XI11_3/XI0/XI0_48/d__0_ xsel_48_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_15 XI11_3/net21_0_ xsel_47_ XI11_3/XI0/XI0_47/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_14 XI11_3/net21_1_ xsel_47_ XI11_3/XI0/XI0_47/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_13 XI11_3/net21_2_ xsel_47_ XI11_3/XI0/XI0_47/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_12 XI11_3/net21_3_ xsel_47_ XI11_3/XI0/XI0_47/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_11 XI11_3/net21_4_ xsel_47_ XI11_3/XI0/XI0_47/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_10 XI11_3/net21_5_ xsel_47_ XI11_3/XI0/XI0_47/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_9 XI11_3/net21_6_ xsel_47_ XI11_3/XI0/XI0_47/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_8 XI11_3/net21_7_ xsel_47_ XI11_3/XI0/XI0_47/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_7 XI11_3/net21_8_ xsel_47_ XI11_3/XI0/XI0_47/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_6 XI11_3/net21_9_ xsel_47_ XI11_3/XI0/XI0_47/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_5 XI11_3/net21_10_ xsel_47_ XI11_3/XI0/XI0_47/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_4 XI11_3/net21_11_ xsel_47_ XI11_3/XI0/XI0_47/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_3 XI11_3/net21_12_ xsel_47_ XI11_3/XI0/XI0_47/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_2 XI11_3/net21_13_ xsel_47_ XI11_3/XI0/XI0_47/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_1 XI11_3/net21_14_ xsel_47_ XI11_3/XI0/XI0_47/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN0_0 XI11_3/net21_15_ xsel_47_ XI11_3/XI0/XI0_47/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_15 XI11_3/XI0/XI0_47/d__15_ xsel_47_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_14 XI11_3/XI0/XI0_47/d__14_ xsel_47_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_13 XI11_3/XI0/XI0_47/d__13_ xsel_47_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_12 XI11_3/XI0/XI0_47/d__12_ xsel_47_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_11 XI11_3/XI0/XI0_47/d__11_ xsel_47_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_10 XI11_3/XI0/XI0_47/d__10_ xsel_47_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_9 XI11_3/XI0/XI0_47/d__9_ xsel_47_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_8 XI11_3/XI0/XI0_47/d__8_ xsel_47_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_7 XI11_3/XI0/XI0_47/d__7_ xsel_47_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_6 XI11_3/XI0/XI0_47/d__6_ xsel_47_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_5 XI11_3/XI0/XI0_47/d__5_ xsel_47_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_4 XI11_3/XI0/XI0_47/d__4_ xsel_47_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_3 XI11_3/XI0/XI0_47/d__3_ xsel_47_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_2 XI11_3/XI0/XI0_47/d__2_ xsel_47_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_1 XI11_3/XI0/XI0_47/d__1_ xsel_47_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_47/MN1_0 XI11_3/XI0/XI0_47/d__0_ xsel_47_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_15 XI11_3/net21_0_ xsel_46_ XI11_3/XI0/XI0_46/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_14 XI11_3/net21_1_ xsel_46_ XI11_3/XI0/XI0_46/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_13 XI11_3/net21_2_ xsel_46_ XI11_3/XI0/XI0_46/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_12 XI11_3/net21_3_ xsel_46_ XI11_3/XI0/XI0_46/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_11 XI11_3/net21_4_ xsel_46_ XI11_3/XI0/XI0_46/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_10 XI11_3/net21_5_ xsel_46_ XI11_3/XI0/XI0_46/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_9 XI11_3/net21_6_ xsel_46_ XI11_3/XI0/XI0_46/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_8 XI11_3/net21_7_ xsel_46_ XI11_3/XI0/XI0_46/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_7 XI11_3/net21_8_ xsel_46_ XI11_3/XI0/XI0_46/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_6 XI11_3/net21_9_ xsel_46_ XI11_3/XI0/XI0_46/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_5 XI11_3/net21_10_ xsel_46_ XI11_3/XI0/XI0_46/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_4 XI11_3/net21_11_ xsel_46_ XI11_3/XI0/XI0_46/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_3 XI11_3/net21_12_ xsel_46_ XI11_3/XI0/XI0_46/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_2 XI11_3/net21_13_ xsel_46_ XI11_3/XI0/XI0_46/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_1 XI11_3/net21_14_ xsel_46_ XI11_3/XI0/XI0_46/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN0_0 XI11_3/net21_15_ xsel_46_ XI11_3/XI0/XI0_46/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_15 XI11_3/XI0/XI0_46/d__15_ xsel_46_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_14 XI11_3/XI0/XI0_46/d__14_ xsel_46_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_13 XI11_3/XI0/XI0_46/d__13_ xsel_46_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_12 XI11_3/XI0/XI0_46/d__12_ xsel_46_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_11 XI11_3/XI0/XI0_46/d__11_ xsel_46_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_10 XI11_3/XI0/XI0_46/d__10_ xsel_46_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_9 XI11_3/XI0/XI0_46/d__9_ xsel_46_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_8 XI11_3/XI0/XI0_46/d__8_ xsel_46_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_7 XI11_3/XI0/XI0_46/d__7_ xsel_46_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_6 XI11_3/XI0/XI0_46/d__6_ xsel_46_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_5 XI11_3/XI0/XI0_46/d__5_ xsel_46_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_4 XI11_3/XI0/XI0_46/d__4_ xsel_46_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_3 XI11_3/XI0/XI0_46/d__3_ xsel_46_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_2 XI11_3/XI0/XI0_46/d__2_ xsel_46_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_1 XI11_3/XI0/XI0_46/d__1_ xsel_46_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_46/MN1_0 XI11_3/XI0/XI0_46/d__0_ xsel_46_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_15 XI11_3/net21_0_ xsel_45_ XI11_3/XI0/XI0_45/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_14 XI11_3/net21_1_ xsel_45_ XI11_3/XI0/XI0_45/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_13 XI11_3/net21_2_ xsel_45_ XI11_3/XI0/XI0_45/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_12 XI11_3/net21_3_ xsel_45_ XI11_3/XI0/XI0_45/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_11 XI11_3/net21_4_ xsel_45_ XI11_3/XI0/XI0_45/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_10 XI11_3/net21_5_ xsel_45_ XI11_3/XI0/XI0_45/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_9 XI11_3/net21_6_ xsel_45_ XI11_3/XI0/XI0_45/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_8 XI11_3/net21_7_ xsel_45_ XI11_3/XI0/XI0_45/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_7 XI11_3/net21_8_ xsel_45_ XI11_3/XI0/XI0_45/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_6 XI11_3/net21_9_ xsel_45_ XI11_3/XI0/XI0_45/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_5 XI11_3/net21_10_ xsel_45_ XI11_3/XI0/XI0_45/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_4 XI11_3/net21_11_ xsel_45_ XI11_3/XI0/XI0_45/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_3 XI11_3/net21_12_ xsel_45_ XI11_3/XI0/XI0_45/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_2 XI11_3/net21_13_ xsel_45_ XI11_3/XI0/XI0_45/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_1 XI11_3/net21_14_ xsel_45_ XI11_3/XI0/XI0_45/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN0_0 XI11_3/net21_15_ xsel_45_ XI11_3/XI0/XI0_45/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_15 XI11_3/XI0/XI0_45/d__15_ xsel_45_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_14 XI11_3/XI0/XI0_45/d__14_ xsel_45_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_13 XI11_3/XI0/XI0_45/d__13_ xsel_45_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_12 XI11_3/XI0/XI0_45/d__12_ xsel_45_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_11 XI11_3/XI0/XI0_45/d__11_ xsel_45_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_10 XI11_3/XI0/XI0_45/d__10_ xsel_45_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_9 XI11_3/XI0/XI0_45/d__9_ xsel_45_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_8 XI11_3/XI0/XI0_45/d__8_ xsel_45_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_7 XI11_3/XI0/XI0_45/d__7_ xsel_45_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_6 XI11_3/XI0/XI0_45/d__6_ xsel_45_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_5 XI11_3/XI0/XI0_45/d__5_ xsel_45_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_4 XI11_3/XI0/XI0_45/d__4_ xsel_45_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_3 XI11_3/XI0/XI0_45/d__3_ xsel_45_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_2 XI11_3/XI0/XI0_45/d__2_ xsel_45_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_1 XI11_3/XI0/XI0_45/d__1_ xsel_45_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_45/MN1_0 XI11_3/XI0/XI0_45/d__0_ xsel_45_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_15 XI11_3/net21_0_ xsel_44_ XI11_3/XI0/XI0_44/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_14 XI11_3/net21_1_ xsel_44_ XI11_3/XI0/XI0_44/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_13 XI11_3/net21_2_ xsel_44_ XI11_3/XI0/XI0_44/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_12 XI11_3/net21_3_ xsel_44_ XI11_3/XI0/XI0_44/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_11 XI11_3/net21_4_ xsel_44_ XI11_3/XI0/XI0_44/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_10 XI11_3/net21_5_ xsel_44_ XI11_3/XI0/XI0_44/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_9 XI11_3/net21_6_ xsel_44_ XI11_3/XI0/XI0_44/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_8 XI11_3/net21_7_ xsel_44_ XI11_3/XI0/XI0_44/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_7 XI11_3/net21_8_ xsel_44_ XI11_3/XI0/XI0_44/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_6 XI11_3/net21_9_ xsel_44_ XI11_3/XI0/XI0_44/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_5 XI11_3/net21_10_ xsel_44_ XI11_3/XI0/XI0_44/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_4 XI11_3/net21_11_ xsel_44_ XI11_3/XI0/XI0_44/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_3 XI11_3/net21_12_ xsel_44_ XI11_3/XI0/XI0_44/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_2 XI11_3/net21_13_ xsel_44_ XI11_3/XI0/XI0_44/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_1 XI11_3/net21_14_ xsel_44_ XI11_3/XI0/XI0_44/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN0_0 XI11_3/net21_15_ xsel_44_ XI11_3/XI0/XI0_44/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_15 XI11_3/XI0/XI0_44/d__15_ xsel_44_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_14 XI11_3/XI0/XI0_44/d__14_ xsel_44_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_13 XI11_3/XI0/XI0_44/d__13_ xsel_44_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_12 XI11_3/XI0/XI0_44/d__12_ xsel_44_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_11 XI11_3/XI0/XI0_44/d__11_ xsel_44_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_10 XI11_3/XI0/XI0_44/d__10_ xsel_44_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_9 XI11_3/XI0/XI0_44/d__9_ xsel_44_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_8 XI11_3/XI0/XI0_44/d__8_ xsel_44_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_7 XI11_3/XI0/XI0_44/d__7_ xsel_44_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_6 XI11_3/XI0/XI0_44/d__6_ xsel_44_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_5 XI11_3/XI0/XI0_44/d__5_ xsel_44_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_4 XI11_3/XI0/XI0_44/d__4_ xsel_44_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_3 XI11_3/XI0/XI0_44/d__3_ xsel_44_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_2 XI11_3/XI0/XI0_44/d__2_ xsel_44_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_1 XI11_3/XI0/XI0_44/d__1_ xsel_44_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_44/MN1_0 XI11_3/XI0/XI0_44/d__0_ xsel_44_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_15 XI11_3/net21_0_ xsel_43_ XI11_3/XI0/XI0_43/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_14 XI11_3/net21_1_ xsel_43_ XI11_3/XI0/XI0_43/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_13 XI11_3/net21_2_ xsel_43_ XI11_3/XI0/XI0_43/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_12 XI11_3/net21_3_ xsel_43_ XI11_3/XI0/XI0_43/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_11 XI11_3/net21_4_ xsel_43_ XI11_3/XI0/XI0_43/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_10 XI11_3/net21_5_ xsel_43_ XI11_3/XI0/XI0_43/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_9 XI11_3/net21_6_ xsel_43_ XI11_3/XI0/XI0_43/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_8 XI11_3/net21_7_ xsel_43_ XI11_3/XI0/XI0_43/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_7 XI11_3/net21_8_ xsel_43_ XI11_3/XI0/XI0_43/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_6 XI11_3/net21_9_ xsel_43_ XI11_3/XI0/XI0_43/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_5 XI11_3/net21_10_ xsel_43_ XI11_3/XI0/XI0_43/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_4 XI11_3/net21_11_ xsel_43_ XI11_3/XI0/XI0_43/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_3 XI11_3/net21_12_ xsel_43_ XI11_3/XI0/XI0_43/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_2 XI11_3/net21_13_ xsel_43_ XI11_3/XI0/XI0_43/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_1 XI11_3/net21_14_ xsel_43_ XI11_3/XI0/XI0_43/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN0_0 XI11_3/net21_15_ xsel_43_ XI11_3/XI0/XI0_43/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_15 XI11_3/XI0/XI0_43/d__15_ xsel_43_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_14 XI11_3/XI0/XI0_43/d__14_ xsel_43_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_13 XI11_3/XI0/XI0_43/d__13_ xsel_43_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_12 XI11_3/XI0/XI0_43/d__12_ xsel_43_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_11 XI11_3/XI0/XI0_43/d__11_ xsel_43_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_10 XI11_3/XI0/XI0_43/d__10_ xsel_43_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_9 XI11_3/XI0/XI0_43/d__9_ xsel_43_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_8 XI11_3/XI0/XI0_43/d__8_ xsel_43_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_7 XI11_3/XI0/XI0_43/d__7_ xsel_43_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_6 XI11_3/XI0/XI0_43/d__6_ xsel_43_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_5 XI11_3/XI0/XI0_43/d__5_ xsel_43_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_4 XI11_3/XI0/XI0_43/d__4_ xsel_43_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_3 XI11_3/XI0/XI0_43/d__3_ xsel_43_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_2 XI11_3/XI0/XI0_43/d__2_ xsel_43_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_1 XI11_3/XI0/XI0_43/d__1_ xsel_43_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_43/MN1_0 XI11_3/XI0/XI0_43/d__0_ xsel_43_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_15 XI11_3/net21_0_ xsel_42_ XI11_3/XI0/XI0_42/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_14 XI11_3/net21_1_ xsel_42_ XI11_3/XI0/XI0_42/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_13 XI11_3/net21_2_ xsel_42_ XI11_3/XI0/XI0_42/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_12 XI11_3/net21_3_ xsel_42_ XI11_3/XI0/XI0_42/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_11 XI11_3/net21_4_ xsel_42_ XI11_3/XI0/XI0_42/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_10 XI11_3/net21_5_ xsel_42_ XI11_3/XI0/XI0_42/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_9 XI11_3/net21_6_ xsel_42_ XI11_3/XI0/XI0_42/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_8 XI11_3/net21_7_ xsel_42_ XI11_3/XI0/XI0_42/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_7 XI11_3/net21_8_ xsel_42_ XI11_3/XI0/XI0_42/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_6 XI11_3/net21_9_ xsel_42_ XI11_3/XI0/XI0_42/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_5 XI11_3/net21_10_ xsel_42_ XI11_3/XI0/XI0_42/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_4 XI11_3/net21_11_ xsel_42_ XI11_3/XI0/XI0_42/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_3 XI11_3/net21_12_ xsel_42_ XI11_3/XI0/XI0_42/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_2 XI11_3/net21_13_ xsel_42_ XI11_3/XI0/XI0_42/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_1 XI11_3/net21_14_ xsel_42_ XI11_3/XI0/XI0_42/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN0_0 XI11_3/net21_15_ xsel_42_ XI11_3/XI0/XI0_42/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_15 XI11_3/XI0/XI0_42/d__15_ xsel_42_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_14 XI11_3/XI0/XI0_42/d__14_ xsel_42_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_13 XI11_3/XI0/XI0_42/d__13_ xsel_42_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_12 XI11_3/XI0/XI0_42/d__12_ xsel_42_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_11 XI11_3/XI0/XI0_42/d__11_ xsel_42_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_10 XI11_3/XI0/XI0_42/d__10_ xsel_42_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_9 XI11_3/XI0/XI0_42/d__9_ xsel_42_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_8 XI11_3/XI0/XI0_42/d__8_ xsel_42_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_7 XI11_3/XI0/XI0_42/d__7_ xsel_42_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_6 XI11_3/XI0/XI0_42/d__6_ xsel_42_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_5 XI11_3/XI0/XI0_42/d__5_ xsel_42_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_4 XI11_3/XI0/XI0_42/d__4_ xsel_42_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_3 XI11_3/XI0/XI0_42/d__3_ xsel_42_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_2 XI11_3/XI0/XI0_42/d__2_ xsel_42_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_1 XI11_3/XI0/XI0_42/d__1_ xsel_42_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_42/MN1_0 XI11_3/XI0/XI0_42/d__0_ xsel_42_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_15 XI11_3/net21_0_ xsel_41_ XI11_3/XI0/XI0_41/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_14 XI11_3/net21_1_ xsel_41_ XI11_3/XI0/XI0_41/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_13 XI11_3/net21_2_ xsel_41_ XI11_3/XI0/XI0_41/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_12 XI11_3/net21_3_ xsel_41_ XI11_3/XI0/XI0_41/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_11 XI11_3/net21_4_ xsel_41_ XI11_3/XI0/XI0_41/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_10 XI11_3/net21_5_ xsel_41_ XI11_3/XI0/XI0_41/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_9 XI11_3/net21_6_ xsel_41_ XI11_3/XI0/XI0_41/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_8 XI11_3/net21_7_ xsel_41_ XI11_3/XI0/XI0_41/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_7 XI11_3/net21_8_ xsel_41_ XI11_3/XI0/XI0_41/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_6 XI11_3/net21_9_ xsel_41_ XI11_3/XI0/XI0_41/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_5 XI11_3/net21_10_ xsel_41_ XI11_3/XI0/XI0_41/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_4 XI11_3/net21_11_ xsel_41_ XI11_3/XI0/XI0_41/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_3 XI11_3/net21_12_ xsel_41_ XI11_3/XI0/XI0_41/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_2 XI11_3/net21_13_ xsel_41_ XI11_3/XI0/XI0_41/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_1 XI11_3/net21_14_ xsel_41_ XI11_3/XI0/XI0_41/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN0_0 XI11_3/net21_15_ xsel_41_ XI11_3/XI0/XI0_41/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_15 XI11_3/XI0/XI0_41/d__15_ xsel_41_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_14 XI11_3/XI0/XI0_41/d__14_ xsel_41_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_13 XI11_3/XI0/XI0_41/d__13_ xsel_41_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_12 XI11_3/XI0/XI0_41/d__12_ xsel_41_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_11 XI11_3/XI0/XI0_41/d__11_ xsel_41_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_10 XI11_3/XI0/XI0_41/d__10_ xsel_41_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_9 XI11_3/XI0/XI0_41/d__9_ xsel_41_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_8 XI11_3/XI0/XI0_41/d__8_ xsel_41_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_7 XI11_3/XI0/XI0_41/d__7_ xsel_41_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_6 XI11_3/XI0/XI0_41/d__6_ xsel_41_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_5 XI11_3/XI0/XI0_41/d__5_ xsel_41_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_4 XI11_3/XI0/XI0_41/d__4_ xsel_41_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_3 XI11_3/XI0/XI0_41/d__3_ xsel_41_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_2 XI11_3/XI0/XI0_41/d__2_ xsel_41_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_1 XI11_3/XI0/XI0_41/d__1_ xsel_41_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_41/MN1_0 XI11_3/XI0/XI0_41/d__0_ xsel_41_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_15 XI11_3/net21_0_ xsel_40_ XI11_3/XI0/XI0_40/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_14 XI11_3/net21_1_ xsel_40_ XI11_3/XI0/XI0_40/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_13 XI11_3/net21_2_ xsel_40_ XI11_3/XI0/XI0_40/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_12 XI11_3/net21_3_ xsel_40_ XI11_3/XI0/XI0_40/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_11 XI11_3/net21_4_ xsel_40_ XI11_3/XI0/XI0_40/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_10 XI11_3/net21_5_ xsel_40_ XI11_3/XI0/XI0_40/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_9 XI11_3/net21_6_ xsel_40_ XI11_3/XI0/XI0_40/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_8 XI11_3/net21_7_ xsel_40_ XI11_3/XI0/XI0_40/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_7 XI11_3/net21_8_ xsel_40_ XI11_3/XI0/XI0_40/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_6 XI11_3/net21_9_ xsel_40_ XI11_3/XI0/XI0_40/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_5 XI11_3/net21_10_ xsel_40_ XI11_3/XI0/XI0_40/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_4 XI11_3/net21_11_ xsel_40_ XI11_3/XI0/XI0_40/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_3 XI11_3/net21_12_ xsel_40_ XI11_3/XI0/XI0_40/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_2 XI11_3/net21_13_ xsel_40_ XI11_3/XI0/XI0_40/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_1 XI11_3/net21_14_ xsel_40_ XI11_3/XI0/XI0_40/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN0_0 XI11_3/net21_15_ xsel_40_ XI11_3/XI0/XI0_40/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_15 XI11_3/XI0/XI0_40/d__15_ xsel_40_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_14 XI11_3/XI0/XI0_40/d__14_ xsel_40_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_13 XI11_3/XI0/XI0_40/d__13_ xsel_40_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_12 XI11_3/XI0/XI0_40/d__12_ xsel_40_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_11 XI11_3/XI0/XI0_40/d__11_ xsel_40_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_10 XI11_3/XI0/XI0_40/d__10_ xsel_40_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_9 XI11_3/XI0/XI0_40/d__9_ xsel_40_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_8 XI11_3/XI0/XI0_40/d__8_ xsel_40_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_7 XI11_3/XI0/XI0_40/d__7_ xsel_40_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_6 XI11_3/XI0/XI0_40/d__6_ xsel_40_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_5 XI11_3/XI0/XI0_40/d__5_ xsel_40_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_4 XI11_3/XI0/XI0_40/d__4_ xsel_40_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_3 XI11_3/XI0/XI0_40/d__3_ xsel_40_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_2 XI11_3/XI0/XI0_40/d__2_ xsel_40_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_1 XI11_3/XI0/XI0_40/d__1_ xsel_40_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_40/MN1_0 XI11_3/XI0/XI0_40/d__0_ xsel_40_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_15 XI11_3/net21_0_ xsel_39_ XI11_3/XI0/XI0_39/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_14 XI11_3/net21_1_ xsel_39_ XI11_3/XI0/XI0_39/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_13 XI11_3/net21_2_ xsel_39_ XI11_3/XI0/XI0_39/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_12 XI11_3/net21_3_ xsel_39_ XI11_3/XI0/XI0_39/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_11 XI11_3/net21_4_ xsel_39_ XI11_3/XI0/XI0_39/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_10 XI11_3/net21_5_ xsel_39_ XI11_3/XI0/XI0_39/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_9 XI11_3/net21_6_ xsel_39_ XI11_3/XI0/XI0_39/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_8 XI11_3/net21_7_ xsel_39_ XI11_3/XI0/XI0_39/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_7 XI11_3/net21_8_ xsel_39_ XI11_3/XI0/XI0_39/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_6 XI11_3/net21_9_ xsel_39_ XI11_3/XI0/XI0_39/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_5 XI11_3/net21_10_ xsel_39_ XI11_3/XI0/XI0_39/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_4 XI11_3/net21_11_ xsel_39_ XI11_3/XI0/XI0_39/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_3 XI11_3/net21_12_ xsel_39_ XI11_3/XI0/XI0_39/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_2 XI11_3/net21_13_ xsel_39_ XI11_3/XI0/XI0_39/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_1 XI11_3/net21_14_ xsel_39_ XI11_3/XI0/XI0_39/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN0_0 XI11_3/net21_15_ xsel_39_ XI11_3/XI0/XI0_39/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_15 XI11_3/XI0/XI0_39/d__15_ xsel_39_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_14 XI11_3/XI0/XI0_39/d__14_ xsel_39_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_13 XI11_3/XI0/XI0_39/d__13_ xsel_39_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_12 XI11_3/XI0/XI0_39/d__12_ xsel_39_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_11 XI11_3/XI0/XI0_39/d__11_ xsel_39_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_10 XI11_3/XI0/XI0_39/d__10_ xsel_39_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_9 XI11_3/XI0/XI0_39/d__9_ xsel_39_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_8 XI11_3/XI0/XI0_39/d__8_ xsel_39_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_7 XI11_3/XI0/XI0_39/d__7_ xsel_39_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_6 XI11_3/XI0/XI0_39/d__6_ xsel_39_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_5 XI11_3/XI0/XI0_39/d__5_ xsel_39_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_4 XI11_3/XI0/XI0_39/d__4_ xsel_39_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_3 XI11_3/XI0/XI0_39/d__3_ xsel_39_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_2 XI11_3/XI0/XI0_39/d__2_ xsel_39_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_1 XI11_3/XI0/XI0_39/d__1_ xsel_39_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_39/MN1_0 XI11_3/XI0/XI0_39/d__0_ xsel_39_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_15 XI11_3/net21_0_ xsel_38_ XI11_3/XI0/XI0_38/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_14 XI11_3/net21_1_ xsel_38_ XI11_3/XI0/XI0_38/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_13 XI11_3/net21_2_ xsel_38_ XI11_3/XI0/XI0_38/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_12 XI11_3/net21_3_ xsel_38_ XI11_3/XI0/XI0_38/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_11 XI11_3/net21_4_ xsel_38_ XI11_3/XI0/XI0_38/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_10 XI11_3/net21_5_ xsel_38_ XI11_3/XI0/XI0_38/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_9 XI11_3/net21_6_ xsel_38_ XI11_3/XI0/XI0_38/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_8 XI11_3/net21_7_ xsel_38_ XI11_3/XI0/XI0_38/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_7 XI11_3/net21_8_ xsel_38_ XI11_3/XI0/XI0_38/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_6 XI11_3/net21_9_ xsel_38_ XI11_3/XI0/XI0_38/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_5 XI11_3/net21_10_ xsel_38_ XI11_3/XI0/XI0_38/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_4 XI11_3/net21_11_ xsel_38_ XI11_3/XI0/XI0_38/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_3 XI11_3/net21_12_ xsel_38_ XI11_3/XI0/XI0_38/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_2 XI11_3/net21_13_ xsel_38_ XI11_3/XI0/XI0_38/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_1 XI11_3/net21_14_ xsel_38_ XI11_3/XI0/XI0_38/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN0_0 XI11_3/net21_15_ xsel_38_ XI11_3/XI0/XI0_38/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_15 XI11_3/XI0/XI0_38/d__15_ xsel_38_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_14 XI11_3/XI0/XI0_38/d__14_ xsel_38_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_13 XI11_3/XI0/XI0_38/d__13_ xsel_38_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_12 XI11_3/XI0/XI0_38/d__12_ xsel_38_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_11 XI11_3/XI0/XI0_38/d__11_ xsel_38_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_10 XI11_3/XI0/XI0_38/d__10_ xsel_38_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_9 XI11_3/XI0/XI0_38/d__9_ xsel_38_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_8 XI11_3/XI0/XI0_38/d__8_ xsel_38_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_7 XI11_3/XI0/XI0_38/d__7_ xsel_38_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_6 XI11_3/XI0/XI0_38/d__6_ xsel_38_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_5 XI11_3/XI0/XI0_38/d__5_ xsel_38_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_4 XI11_3/XI0/XI0_38/d__4_ xsel_38_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_3 XI11_3/XI0/XI0_38/d__3_ xsel_38_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_2 XI11_3/XI0/XI0_38/d__2_ xsel_38_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_1 XI11_3/XI0/XI0_38/d__1_ xsel_38_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_38/MN1_0 XI11_3/XI0/XI0_38/d__0_ xsel_38_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_15 XI11_3/net21_0_ xsel_37_ XI11_3/XI0/XI0_37/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_14 XI11_3/net21_1_ xsel_37_ XI11_3/XI0/XI0_37/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_13 XI11_3/net21_2_ xsel_37_ XI11_3/XI0/XI0_37/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_12 XI11_3/net21_3_ xsel_37_ XI11_3/XI0/XI0_37/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_11 XI11_3/net21_4_ xsel_37_ XI11_3/XI0/XI0_37/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_10 XI11_3/net21_5_ xsel_37_ XI11_3/XI0/XI0_37/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_9 XI11_3/net21_6_ xsel_37_ XI11_3/XI0/XI0_37/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_8 XI11_3/net21_7_ xsel_37_ XI11_3/XI0/XI0_37/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_7 XI11_3/net21_8_ xsel_37_ XI11_3/XI0/XI0_37/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_6 XI11_3/net21_9_ xsel_37_ XI11_3/XI0/XI0_37/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_5 XI11_3/net21_10_ xsel_37_ XI11_3/XI0/XI0_37/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_4 XI11_3/net21_11_ xsel_37_ XI11_3/XI0/XI0_37/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_3 XI11_3/net21_12_ xsel_37_ XI11_3/XI0/XI0_37/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_2 XI11_3/net21_13_ xsel_37_ XI11_3/XI0/XI0_37/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_1 XI11_3/net21_14_ xsel_37_ XI11_3/XI0/XI0_37/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN0_0 XI11_3/net21_15_ xsel_37_ XI11_3/XI0/XI0_37/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_15 XI11_3/XI0/XI0_37/d__15_ xsel_37_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_14 XI11_3/XI0/XI0_37/d__14_ xsel_37_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_13 XI11_3/XI0/XI0_37/d__13_ xsel_37_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_12 XI11_3/XI0/XI0_37/d__12_ xsel_37_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_11 XI11_3/XI0/XI0_37/d__11_ xsel_37_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_10 XI11_3/XI0/XI0_37/d__10_ xsel_37_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_9 XI11_3/XI0/XI0_37/d__9_ xsel_37_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_8 XI11_3/XI0/XI0_37/d__8_ xsel_37_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_7 XI11_3/XI0/XI0_37/d__7_ xsel_37_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_6 XI11_3/XI0/XI0_37/d__6_ xsel_37_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_5 XI11_3/XI0/XI0_37/d__5_ xsel_37_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_4 XI11_3/XI0/XI0_37/d__4_ xsel_37_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_3 XI11_3/XI0/XI0_37/d__3_ xsel_37_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_2 XI11_3/XI0/XI0_37/d__2_ xsel_37_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_1 XI11_3/XI0/XI0_37/d__1_ xsel_37_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_37/MN1_0 XI11_3/XI0/XI0_37/d__0_ xsel_37_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_15 XI11_3/net21_0_ xsel_36_ XI11_3/XI0/XI0_36/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_14 XI11_3/net21_1_ xsel_36_ XI11_3/XI0/XI0_36/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_13 XI11_3/net21_2_ xsel_36_ XI11_3/XI0/XI0_36/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_12 XI11_3/net21_3_ xsel_36_ XI11_3/XI0/XI0_36/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_11 XI11_3/net21_4_ xsel_36_ XI11_3/XI0/XI0_36/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_10 XI11_3/net21_5_ xsel_36_ XI11_3/XI0/XI0_36/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_9 XI11_3/net21_6_ xsel_36_ XI11_3/XI0/XI0_36/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_8 XI11_3/net21_7_ xsel_36_ XI11_3/XI0/XI0_36/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_7 XI11_3/net21_8_ xsel_36_ XI11_3/XI0/XI0_36/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_6 XI11_3/net21_9_ xsel_36_ XI11_3/XI0/XI0_36/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_5 XI11_3/net21_10_ xsel_36_ XI11_3/XI0/XI0_36/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_4 XI11_3/net21_11_ xsel_36_ XI11_3/XI0/XI0_36/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_3 XI11_3/net21_12_ xsel_36_ XI11_3/XI0/XI0_36/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_2 XI11_3/net21_13_ xsel_36_ XI11_3/XI0/XI0_36/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_1 XI11_3/net21_14_ xsel_36_ XI11_3/XI0/XI0_36/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN0_0 XI11_3/net21_15_ xsel_36_ XI11_3/XI0/XI0_36/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_15 XI11_3/XI0/XI0_36/d__15_ xsel_36_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_14 XI11_3/XI0/XI0_36/d__14_ xsel_36_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_13 XI11_3/XI0/XI0_36/d__13_ xsel_36_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_12 XI11_3/XI0/XI0_36/d__12_ xsel_36_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_11 XI11_3/XI0/XI0_36/d__11_ xsel_36_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_10 XI11_3/XI0/XI0_36/d__10_ xsel_36_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_9 XI11_3/XI0/XI0_36/d__9_ xsel_36_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_8 XI11_3/XI0/XI0_36/d__8_ xsel_36_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_7 XI11_3/XI0/XI0_36/d__7_ xsel_36_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_6 XI11_3/XI0/XI0_36/d__6_ xsel_36_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_5 XI11_3/XI0/XI0_36/d__5_ xsel_36_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_4 XI11_3/XI0/XI0_36/d__4_ xsel_36_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_3 XI11_3/XI0/XI0_36/d__3_ xsel_36_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_2 XI11_3/XI0/XI0_36/d__2_ xsel_36_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_1 XI11_3/XI0/XI0_36/d__1_ xsel_36_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_36/MN1_0 XI11_3/XI0/XI0_36/d__0_ xsel_36_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_15 XI11_3/net21_0_ xsel_35_ XI11_3/XI0/XI0_35/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_14 XI11_3/net21_1_ xsel_35_ XI11_3/XI0/XI0_35/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_13 XI11_3/net21_2_ xsel_35_ XI11_3/XI0/XI0_35/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_12 XI11_3/net21_3_ xsel_35_ XI11_3/XI0/XI0_35/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_11 XI11_3/net21_4_ xsel_35_ XI11_3/XI0/XI0_35/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_10 XI11_3/net21_5_ xsel_35_ XI11_3/XI0/XI0_35/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_9 XI11_3/net21_6_ xsel_35_ XI11_3/XI0/XI0_35/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_8 XI11_3/net21_7_ xsel_35_ XI11_3/XI0/XI0_35/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_7 XI11_3/net21_8_ xsel_35_ XI11_3/XI0/XI0_35/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_6 XI11_3/net21_9_ xsel_35_ XI11_3/XI0/XI0_35/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_5 XI11_3/net21_10_ xsel_35_ XI11_3/XI0/XI0_35/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_4 XI11_3/net21_11_ xsel_35_ XI11_3/XI0/XI0_35/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_3 XI11_3/net21_12_ xsel_35_ XI11_3/XI0/XI0_35/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_2 XI11_3/net21_13_ xsel_35_ XI11_3/XI0/XI0_35/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_1 XI11_3/net21_14_ xsel_35_ XI11_3/XI0/XI0_35/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN0_0 XI11_3/net21_15_ xsel_35_ XI11_3/XI0/XI0_35/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_15 XI11_3/XI0/XI0_35/d__15_ xsel_35_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_14 XI11_3/XI0/XI0_35/d__14_ xsel_35_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_13 XI11_3/XI0/XI0_35/d__13_ xsel_35_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_12 XI11_3/XI0/XI0_35/d__12_ xsel_35_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_11 XI11_3/XI0/XI0_35/d__11_ xsel_35_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_10 XI11_3/XI0/XI0_35/d__10_ xsel_35_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_9 XI11_3/XI0/XI0_35/d__9_ xsel_35_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_8 XI11_3/XI0/XI0_35/d__8_ xsel_35_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_7 XI11_3/XI0/XI0_35/d__7_ xsel_35_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_6 XI11_3/XI0/XI0_35/d__6_ xsel_35_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_5 XI11_3/XI0/XI0_35/d__5_ xsel_35_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_4 XI11_3/XI0/XI0_35/d__4_ xsel_35_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_3 XI11_3/XI0/XI0_35/d__3_ xsel_35_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_2 XI11_3/XI0/XI0_35/d__2_ xsel_35_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_1 XI11_3/XI0/XI0_35/d__1_ xsel_35_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_35/MN1_0 XI11_3/XI0/XI0_35/d__0_ xsel_35_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_15 XI11_3/net21_0_ xsel_34_ XI11_3/XI0/XI0_34/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_14 XI11_3/net21_1_ xsel_34_ XI11_3/XI0/XI0_34/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_13 XI11_3/net21_2_ xsel_34_ XI11_3/XI0/XI0_34/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_12 XI11_3/net21_3_ xsel_34_ XI11_3/XI0/XI0_34/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_11 XI11_3/net21_4_ xsel_34_ XI11_3/XI0/XI0_34/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_10 XI11_3/net21_5_ xsel_34_ XI11_3/XI0/XI0_34/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_9 XI11_3/net21_6_ xsel_34_ XI11_3/XI0/XI0_34/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_8 XI11_3/net21_7_ xsel_34_ XI11_3/XI0/XI0_34/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_7 XI11_3/net21_8_ xsel_34_ XI11_3/XI0/XI0_34/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_6 XI11_3/net21_9_ xsel_34_ XI11_3/XI0/XI0_34/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_5 XI11_3/net21_10_ xsel_34_ XI11_3/XI0/XI0_34/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_4 XI11_3/net21_11_ xsel_34_ XI11_3/XI0/XI0_34/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_3 XI11_3/net21_12_ xsel_34_ XI11_3/XI0/XI0_34/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_2 XI11_3/net21_13_ xsel_34_ XI11_3/XI0/XI0_34/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_1 XI11_3/net21_14_ xsel_34_ XI11_3/XI0/XI0_34/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN0_0 XI11_3/net21_15_ xsel_34_ XI11_3/XI0/XI0_34/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_15 XI11_3/XI0/XI0_34/d__15_ xsel_34_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_14 XI11_3/XI0/XI0_34/d__14_ xsel_34_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_13 XI11_3/XI0/XI0_34/d__13_ xsel_34_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_12 XI11_3/XI0/XI0_34/d__12_ xsel_34_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_11 XI11_3/XI0/XI0_34/d__11_ xsel_34_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_10 XI11_3/XI0/XI0_34/d__10_ xsel_34_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_9 XI11_3/XI0/XI0_34/d__9_ xsel_34_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_8 XI11_3/XI0/XI0_34/d__8_ xsel_34_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_7 XI11_3/XI0/XI0_34/d__7_ xsel_34_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_6 XI11_3/XI0/XI0_34/d__6_ xsel_34_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_5 XI11_3/XI0/XI0_34/d__5_ xsel_34_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_4 XI11_3/XI0/XI0_34/d__4_ xsel_34_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_3 XI11_3/XI0/XI0_34/d__3_ xsel_34_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_2 XI11_3/XI0/XI0_34/d__2_ xsel_34_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_1 XI11_3/XI0/XI0_34/d__1_ xsel_34_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_34/MN1_0 XI11_3/XI0/XI0_34/d__0_ xsel_34_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_15 XI11_3/net21_0_ xsel_33_ XI11_3/XI0/XI0_33/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_14 XI11_3/net21_1_ xsel_33_ XI11_3/XI0/XI0_33/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_13 XI11_3/net21_2_ xsel_33_ XI11_3/XI0/XI0_33/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_12 XI11_3/net21_3_ xsel_33_ XI11_3/XI0/XI0_33/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_11 XI11_3/net21_4_ xsel_33_ XI11_3/XI0/XI0_33/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_10 XI11_3/net21_5_ xsel_33_ XI11_3/XI0/XI0_33/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_9 XI11_3/net21_6_ xsel_33_ XI11_3/XI0/XI0_33/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_8 XI11_3/net21_7_ xsel_33_ XI11_3/XI0/XI0_33/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_7 XI11_3/net21_8_ xsel_33_ XI11_3/XI0/XI0_33/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_6 XI11_3/net21_9_ xsel_33_ XI11_3/XI0/XI0_33/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_5 XI11_3/net21_10_ xsel_33_ XI11_3/XI0/XI0_33/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_4 XI11_3/net21_11_ xsel_33_ XI11_3/XI0/XI0_33/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_3 XI11_3/net21_12_ xsel_33_ XI11_3/XI0/XI0_33/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_2 XI11_3/net21_13_ xsel_33_ XI11_3/XI0/XI0_33/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_1 XI11_3/net21_14_ xsel_33_ XI11_3/XI0/XI0_33/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN0_0 XI11_3/net21_15_ xsel_33_ XI11_3/XI0/XI0_33/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_15 XI11_3/XI0/XI0_33/d__15_ xsel_33_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_14 XI11_3/XI0/XI0_33/d__14_ xsel_33_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_13 XI11_3/XI0/XI0_33/d__13_ xsel_33_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_12 XI11_3/XI0/XI0_33/d__12_ xsel_33_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_11 XI11_3/XI0/XI0_33/d__11_ xsel_33_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_10 XI11_3/XI0/XI0_33/d__10_ xsel_33_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_9 XI11_3/XI0/XI0_33/d__9_ xsel_33_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_8 XI11_3/XI0/XI0_33/d__8_ xsel_33_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_7 XI11_3/XI0/XI0_33/d__7_ xsel_33_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_6 XI11_3/XI0/XI0_33/d__6_ xsel_33_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_5 XI11_3/XI0/XI0_33/d__5_ xsel_33_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_4 XI11_3/XI0/XI0_33/d__4_ xsel_33_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_3 XI11_3/XI0/XI0_33/d__3_ xsel_33_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_2 XI11_3/XI0/XI0_33/d__2_ xsel_33_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_1 XI11_3/XI0/XI0_33/d__1_ xsel_33_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_33/MN1_0 XI11_3/XI0/XI0_33/d__0_ xsel_33_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_15 XI11_3/net21_0_ xsel_32_ XI11_3/XI0/XI0_32/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_14 XI11_3/net21_1_ xsel_32_ XI11_3/XI0/XI0_32/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_13 XI11_3/net21_2_ xsel_32_ XI11_3/XI0/XI0_32/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_12 XI11_3/net21_3_ xsel_32_ XI11_3/XI0/XI0_32/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_11 XI11_3/net21_4_ xsel_32_ XI11_3/XI0/XI0_32/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_10 XI11_3/net21_5_ xsel_32_ XI11_3/XI0/XI0_32/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_9 XI11_3/net21_6_ xsel_32_ XI11_3/XI0/XI0_32/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_8 XI11_3/net21_7_ xsel_32_ XI11_3/XI0/XI0_32/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_7 XI11_3/net21_8_ xsel_32_ XI11_3/XI0/XI0_32/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_6 XI11_3/net21_9_ xsel_32_ XI11_3/XI0/XI0_32/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_5 XI11_3/net21_10_ xsel_32_ XI11_3/XI0/XI0_32/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_4 XI11_3/net21_11_ xsel_32_ XI11_3/XI0/XI0_32/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_3 XI11_3/net21_12_ xsel_32_ XI11_3/XI0/XI0_32/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_2 XI11_3/net21_13_ xsel_32_ XI11_3/XI0/XI0_32/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_1 XI11_3/net21_14_ xsel_32_ XI11_3/XI0/XI0_32/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN0_0 XI11_3/net21_15_ xsel_32_ XI11_3/XI0/XI0_32/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_15 XI11_3/XI0/XI0_32/d__15_ xsel_32_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_14 XI11_3/XI0/XI0_32/d__14_ xsel_32_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_13 XI11_3/XI0/XI0_32/d__13_ xsel_32_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_12 XI11_3/XI0/XI0_32/d__12_ xsel_32_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_11 XI11_3/XI0/XI0_32/d__11_ xsel_32_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_10 XI11_3/XI0/XI0_32/d__10_ xsel_32_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_9 XI11_3/XI0/XI0_32/d__9_ xsel_32_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_8 XI11_3/XI0/XI0_32/d__8_ xsel_32_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_7 XI11_3/XI0/XI0_32/d__7_ xsel_32_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_6 XI11_3/XI0/XI0_32/d__6_ xsel_32_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_5 XI11_3/XI0/XI0_32/d__5_ xsel_32_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_4 XI11_3/XI0/XI0_32/d__4_ xsel_32_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_3 XI11_3/XI0/XI0_32/d__3_ xsel_32_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_2 XI11_3/XI0/XI0_32/d__2_ xsel_32_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_1 XI11_3/XI0/XI0_32/d__1_ xsel_32_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_32/MN1_0 XI11_3/XI0/XI0_32/d__0_ xsel_32_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_15 XI11_3/net21_0_ xsel_31_ XI11_3/XI0/XI0_31/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_14 XI11_3/net21_1_ xsel_31_ XI11_3/XI0/XI0_31/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_13 XI11_3/net21_2_ xsel_31_ XI11_3/XI0/XI0_31/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_12 XI11_3/net21_3_ xsel_31_ XI11_3/XI0/XI0_31/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_11 XI11_3/net21_4_ xsel_31_ XI11_3/XI0/XI0_31/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_10 XI11_3/net21_5_ xsel_31_ XI11_3/XI0/XI0_31/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_9 XI11_3/net21_6_ xsel_31_ XI11_3/XI0/XI0_31/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_8 XI11_3/net21_7_ xsel_31_ XI11_3/XI0/XI0_31/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_7 XI11_3/net21_8_ xsel_31_ XI11_3/XI0/XI0_31/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_6 XI11_3/net21_9_ xsel_31_ XI11_3/XI0/XI0_31/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_5 XI11_3/net21_10_ xsel_31_ XI11_3/XI0/XI0_31/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_4 XI11_3/net21_11_ xsel_31_ XI11_3/XI0/XI0_31/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_3 XI11_3/net21_12_ xsel_31_ XI11_3/XI0/XI0_31/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_2 XI11_3/net21_13_ xsel_31_ XI11_3/XI0/XI0_31/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_1 XI11_3/net21_14_ xsel_31_ XI11_3/XI0/XI0_31/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN0_0 XI11_3/net21_15_ xsel_31_ XI11_3/XI0/XI0_31/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_15 XI11_3/XI0/XI0_31/d__15_ xsel_31_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_14 XI11_3/XI0/XI0_31/d__14_ xsel_31_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_13 XI11_3/XI0/XI0_31/d__13_ xsel_31_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_12 XI11_3/XI0/XI0_31/d__12_ xsel_31_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_11 XI11_3/XI0/XI0_31/d__11_ xsel_31_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_10 XI11_3/XI0/XI0_31/d__10_ xsel_31_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_9 XI11_3/XI0/XI0_31/d__9_ xsel_31_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_8 XI11_3/XI0/XI0_31/d__8_ xsel_31_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_7 XI11_3/XI0/XI0_31/d__7_ xsel_31_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_6 XI11_3/XI0/XI0_31/d__6_ xsel_31_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_5 XI11_3/XI0/XI0_31/d__5_ xsel_31_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_4 XI11_3/XI0/XI0_31/d__4_ xsel_31_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_3 XI11_3/XI0/XI0_31/d__3_ xsel_31_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_2 XI11_3/XI0/XI0_31/d__2_ xsel_31_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_1 XI11_3/XI0/XI0_31/d__1_ xsel_31_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_31/MN1_0 XI11_3/XI0/XI0_31/d__0_ xsel_31_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_15 XI11_3/net21_0_ xsel_30_ XI11_3/XI0/XI0_30/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_14 XI11_3/net21_1_ xsel_30_ XI11_3/XI0/XI0_30/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_13 XI11_3/net21_2_ xsel_30_ XI11_3/XI0/XI0_30/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_12 XI11_3/net21_3_ xsel_30_ XI11_3/XI0/XI0_30/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_11 XI11_3/net21_4_ xsel_30_ XI11_3/XI0/XI0_30/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_10 XI11_3/net21_5_ xsel_30_ XI11_3/XI0/XI0_30/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_9 XI11_3/net21_6_ xsel_30_ XI11_3/XI0/XI0_30/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_8 XI11_3/net21_7_ xsel_30_ XI11_3/XI0/XI0_30/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_7 XI11_3/net21_8_ xsel_30_ XI11_3/XI0/XI0_30/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_6 XI11_3/net21_9_ xsel_30_ XI11_3/XI0/XI0_30/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_5 XI11_3/net21_10_ xsel_30_ XI11_3/XI0/XI0_30/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_4 XI11_3/net21_11_ xsel_30_ XI11_3/XI0/XI0_30/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_3 XI11_3/net21_12_ xsel_30_ XI11_3/XI0/XI0_30/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_2 XI11_3/net21_13_ xsel_30_ XI11_3/XI0/XI0_30/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_1 XI11_3/net21_14_ xsel_30_ XI11_3/XI0/XI0_30/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN0_0 XI11_3/net21_15_ xsel_30_ XI11_3/XI0/XI0_30/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_15 XI11_3/XI0/XI0_30/d__15_ xsel_30_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_14 XI11_3/XI0/XI0_30/d__14_ xsel_30_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_13 XI11_3/XI0/XI0_30/d__13_ xsel_30_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_12 XI11_3/XI0/XI0_30/d__12_ xsel_30_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_11 XI11_3/XI0/XI0_30/d__11_ xsel_30_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_10 XI11_3/XI0/XI0_30/d__10_ xsel_30_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_9 XI11_3/XI0/XI0_30/d__9_ xsel_30_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_8 XI11_3/XI0/XI0_30/d__8_ xsel_30_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_7 XI11_3/XI0/XI0_30/d__7_ xsel_30_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_6 XI11_3/XI0/XI0_30/d__6_ xsel_30_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_5 XI11_3/XI0/XI0_30/d__5_ xsel_30_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_4 XI11_3/XI0/XI0_30/d__4_ xsel_30_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_3 XI11_3/XI0/XI0_30/d__3_ xsel_30_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_2 XI11_3/XI0/XI0_30/d__2_ xsel_30_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_1 XI11_3/XI0/XI0_30/d__1_ xsel_30_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_30/MN1_0 XI11_3/XI0/XI0_30/d__0_ xsel_30_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_15 XI11_3/net21_0_ xsel_29_ XI11_3/XI0/XI0_29/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_14 XI11_3/net21_1_ xsel_29_ XI11_3/XI0/XI0_29/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_13 XI11_3/net21_2_ xsel_29_ XI11_3/XI0/XI0_29/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_12 XI11_3/net21_3_ xsel_29_ XI11_3/XI0/XI0_29/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_11 XI11_3/net21_4_ xsel_29_ XI11_3/XI0/XI0_29/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_10 XI11_3/net21_5_ xsel_29_ XI11_3/XI0/XI0_29/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_9 XI11_3/net21_6_ xsel_29_ XI11_3/XI0/XI0_29/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_8 XI11_3/net21_7_ xsel_29_ XI11_3/XI0/XI0_29/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_7 XI11_3/net21_8_ xsel_29_ XI11_3/XI0/XI0_29/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_6 XI11_3/net21_9_ xsel_29_ XI11_3/XI0/XI0_29/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_5 XI11_3/net21_10_ xsel_29_ XI11_3/XI0/XI0_29/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_4 XI11_3/net21_11_ xsel_29_ XI11_3/XI0/XI0_29/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_3 XI11_3/net21_12_ xsel_29_ XI11_3/XI0/XI0_29/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_2 XI11_3/net21_13_ xsel_29_ XI11_3/XI0/XI0_29/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_1 XI11_3/net21_14_ xsel_29_ XI11_3/XI0/XI0_29/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN0_0 XI11_3/net21_15_ xsel_29_ XI11_3/XI0/XI0_29/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_15 XI11_3/XI0/XI0_29/d__15_ xsel_29_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_14 XI11_3/XI0/XI0_29/d__14_ xsel_29_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_13 XI11_3/XI0/XI0_29/d__13_ xsel_29_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_12 XI11_3/XI0/XI0_29/d__12_ xsel_29_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_11 XI11_3/XI0/XI0_29/d__11_ xsel_29_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_10 XI11_3/XI0/XI0_29/d__10_ xsel_29_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_9 XI11_3/XI0/XI0_29/d__9_ xsel_29_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_8 XI11_3/XI0/XI0_29/d__8_ xsel_29_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_7 XI11_3/XI0/XI0_29/d__7_ xsel_29_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_6 XI11_3/XI0/XI0_29/d__6_ xsel_29_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_5 XI11_3/XI0/XI0_29/d__5_ xsel_29_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_4 XI11_3/XI0/XI0_29/d__4_ xsel_29_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_3 XI11_3/XI0/XI0_29/d__3_ xsel_29_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_2 XI11_3/XI0/XI0_29/d__2_ xsel_29_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_1 XI11_3/XI0/XI0_29/d__1_ xsel_29_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_29/MN1_0 XI11_3/XI0/XI0_29/d__0_ xsel_29_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_15 XI11_3/net21_0_ xsel_28_ XI11_3/XI0/XI0_28/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_14 XI11_3/net21_1_ xsel_28_ XI11_3/XI0/XI0_28/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_13 XI11_3/net21_2_ xsel_28_ XI11_3/XI0/XI0_28/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_12 XI11_3/net21_3_ xsel_28_ XI11_3/XI0/XI0_28/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_11 XI11_3/net21_4_ xsel_28_ XI11_3/XI0/XI0_28/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_10 XI11_3/net21_5_ xsel_28_ XI11_3/XI0/XI0_28/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_9 XI11_3/net21_6_ xsel_28_ XI11_3/XI0/XI0_28/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_8 XI11_3/net21_7_ xsel_28_ XI11_3/XI0/XI0_28/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_7 XI11_3/net21_8_ xsel_28_ XI11_3/XI0/XI0_28/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_6 XI11_3/net21_9_ xsel_28_ XI11_3/XI0/XI0_28/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_5 XI11_3/net21_10_ xsel_28_ XI11_3/XI0/XI0_28/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_4 XI11_3/net21_11_ xsel_28_ XI11_3/XI0/XI0_28/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_3 XI11_3/net21_12_ xsel_28_ XI11_3/XI0/XI0_28/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_2 XI11_3/net21_13_ xsel_28_ XI11_3/XI0/XI0_28/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_1 XI11_3/net21_14_ xsel_28_ XI11_3/XI0/XI0_28/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN0_0 XI11_3/net21_15_ xsel_28_ XI11_3/XI0/XI0_28/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_15 XI11_3/XI0/XI0_28/d__15_ xsel_28_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_14 XI11_3/XI0/XI0_28/d__14_ xsel_28_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_13 XI11_3/XI0/XI0_28/d__13_ xsel_28_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_12 XI11_3/XI0/XI0_28/d__12_ xsel_28_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_11 XI11_3/XI0/XI0_28/d__11_ xsel_28_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_10 XI11_3/XI0/XI0_28/d__10_ xsel_28_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_9 XI11_3/XI0/XI0_28/d__9_ xsel_28_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_8 XI11_3/XI0/XI0_28/d__8_ xsel_28_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_7 XI11_3/XI0/XI0_28/d__7_ xsel_28_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_6 XI11_3/XI0/XI0_28/d__6_ xsel_28_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_5 XI11_3/XI0/XI0_28/d__5_ xsel_28_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_4 XI11_3/XI0/XI0_28/d__4_ xsel_28_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_3 XI11_3/XI0/XI0_28/d__3_ xsel_28_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_2 XI11_3/XI0/XI0_28/d__2_ xsel_28_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_1 XI11_3/XI0/XI0_28/d__1_ xsel_28_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_28/MN1_0 XI11_3/XI0/XI0_28/d__0_ xsel_28_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_15 XI11_3/net21_0_ xsel_27_ XI11_3/XI0/XI0_27/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_14 XI11_3/net21_1_ xsel_27_ XI11_3/XI0/XI0_27/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_13 XI11_3/net21_2_ xsel_27_ XI11_3/XI0/XI0_27/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_12 XI11_3/net21_3_ xsel_27_ XI11_3/XI0/XI0_27/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_11 XI11_3/net21_4_ xsel_27_ XI11_3/XI0/XI0_27/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_10 XI11_3/net21_5_ xsel_27_ XI11_3/XI0/XI0_27/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_9 XI11_3/net21_6_ xsel_27_ XI11_3/XI0/XI0_27/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_8 XI11_3/net21_7_ xsel_27_ XI11_3/XI0/XI0_27/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_7 XI11_3/net21_8_ xsel_27_ XI11_3/XI0/XI0_27/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_6 XI11_3/net21_9_ xsel_27_ XI11_3/XI0/XI0_27/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_5 XI11_3/net21_10_ xsel_27_ XI11_3/XI0/XI0_27/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_4 XI11_3/net21_11_ xsel_27_ XI11_3/XI0/XI0_27/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_3 XI11_3/net21_12_ xsel_27_ XI11_3/XI0/XI0_27/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_2 XI11_3/net21_13_ xsel_27_ XI11_3/XI0/XI0_27/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_1 XI11_3/net21_14_ xsel_27_ XI11_3/XI0/XI0_27/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN0_0 XI11_3/net21_15_ xsel_27_ XI11_3/XI0/XI0_27/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_15 XI11_3/XI0/XI0_27/d__15_ xsel_27_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_14 XI11_3/XI0/XI0_27/d__14_ xsel_27_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_13 XI11_3/XI0/XI0_27/d__13_ xsel_27_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_12 XI11_3/XI0/XI0_27/d__12_ xsel_27_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_11 XI11_3/XI0/XI0_27/d__11_ xsel_27_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_10 XI11_3/XI0/XI0_27/d__10_ xsel_27_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_9 XI11_3/XI0/XI0_27/d__9_ xsel_27_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_8 XI11_3/XI0/XI0_27/d__8_ xsel_27_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_7 XI11_3/XI0/XI0_27/d__7_ xsel_27_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_6 XI11_3/XI0/XI0_27/d__6_ xsel_27_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_5 XI11_3/XI0/XI0_27/d__5_ xsel_27_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_4 XI11_3/XI0/XI0_27/d__4_ xsel_27_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_3 XI11_3/XI0/XI0_27/d__3_ xsel_27_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_2 XI11_3/XI0/XI0_27/d__2_ xsel_27_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_1 XI11_3/XI0/XI0_27/d__1_ xsel_27_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_27/MN1_0 XI11_3/XI0/XI0_27/d__0_ xsel_27_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_15 XI11_3/net21_0_ xsel_26_ XI11_3/XI0/XI0_26/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_14 XI11_3/net21_1_ xsel_26_ XI11_3/XI0/XI0_26/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_13 XI11_3/net21_2_ xsel_26_ XI11_3/XI0/XI0_26/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_12 XI11_3/net21_3_ xsel_26_ XI11_3/XI0/XI0_26/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_11 XI11_3/net21_4_ xsel_26_ XI11_3/XI0/XI0_26/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_10 XI11_3/net21_5_ xsel_26_ XI11_3/XI0/XI0_26/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_9 XI11_3/net21_6_ xsel_26_ XI11_3/XI0/XI0_26/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_8 XI11_3/net21_7_ xsel_26_ XI11_3/XI0/XI0_26/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_7 XI11_3/net21_8_ xsel_26_ XI11_3/XI0/XI0_26/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_6 XI11_3/net21_9_ xsel_26_ XI11_3/XI0/XI0_26/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_5 XI11_3/net21_10_ xsel_26_ XI11_3/XI0/XI0_26/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_4 XI11_3/net21_11_ xsel_26_ XI11_3/XI0/XI0_26/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_3 XI11_3/net21_12_ xsel_26_ XI11_3/XI0/XI0_26/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_2 XI11_3/net21_13_ xsel_26_ XI11_3/XI0/XI0_26/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_1 XI11_3/net21_14_ xsel_26_ XI11_3/XI0/XI0_26/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN0_0 XI11_3/net21_15_ xsel_26_ XI11_3/XI0/XI0_26/d_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_15 XI11_3/XI0/XI0_26/d__15_ xsel_26_ XI11_3/net20_0_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_14 XI11_3/XI0/XI0_26/d__14_ xsel_26_ XI11_3/net20_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_13 XI11_3/XI0/XI0_26/d__13_ xsel_26_ XI11_3/net20_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_12 XI11_3/XI0/XI0_26/d__12_ xsel_26_ XI11_3/net20_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_11 XI11_3/XI0/XI0_26/d__11_ xsel_26_ XI11_3/net20_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_10 XI11_3/XI0/XI0_26/d__10_ xsel_26_ XI11_3/net20_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_9 XI11_3/XI0/XI0_26/d__9_ xsel_26_ XI11_3/net20_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_8 XI11_3/XI0/XI0_26/d__8_ xsel_26_ XI11_3/net20_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_7 XI11_3/XI0/XI0_26/d__7_ xsel_26_ XI11_3/net20_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_6 XI11_3/XI0/XI0_26/d__6_ xsel_26_ XI11_3/net20_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_5 XI11_3/XI0/XI0_26/d__5_ xsel_26_ XI11_3/net20_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_4 XI11_3/XI0/XI0_26/d__4_ xsel_26_ XI11_3/net20_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_3 XI11_3/XI0/XI0_26/d__3_ xsel_26_ XI11_3/net20_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_2 XI11_3/XI0/XI0_26/d__2_ xsel_26_ XI11_3/net20_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_1 XI11_3/XI0/XI0_26/d__1_ xsel_26_ XI11_3/net20_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_26/MN1_0 XI11_3/XI0/XI0_26/d__0_ xsel_26_ XI11_3/net20_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_15 XI11_3/net21_0_ xsel_25_ XI11_3/XI0/XI0_25/d_15_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_14 XI11_3/net21_1_ xsel_25_ XI11_3/XI0/XI0_25/d_14_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_13 XI11_3/net21_2_ xsel_25_ XI11_3/XI0/XI0_25/d_13_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_12 XI11_3/net21_3_ xsel_25_ XI11_3/XI0/XI0_25/d_12_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_11 XI11_3/net21_4_ xsel_25_ XI11_3/XI0/XI0_25/d_11_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_10 XI11_3/net21_5_ xsel_25_ XI11_3/XI0/XI0_25/d_10_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_9 XI11_3/net21_6_ xsel_25_ XI11_3/XI0/XI0_25/d_9_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_8 XI11_3/net21_7_ xsel_25_ XI11_3/XI0/XI0_25/d_8_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_7 XI11_3/net21_8_ xsel_25_ XI11_3/XI0/XI0_25/d_7_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_6 XI11_3/net21_9_ xsel_25_ XI11_3/XI0/XI0_25/d_6_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_5 XI11_3/net21_10_ xsel_25_ XI11_3/XI0/XI0_25/d_5_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_4 XI11_3/net21_11_ xsel_25_ XI11_3/XI0/XI0_25/d_4_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_3 XI11_3/net21_12_ xsel_25_ XI11_3/XI0/XI0_25/d_3_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_2 XI11_3/net21_13_ xsel_25_ XI11_3/XI0/XI0_25/d_2_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll] 
XI11_3/XI0/XI0_25/MN0_1 XI11_3/net21_14_ xsel_25_ XI11_3/XI0/XI0_25/d_1_ gnd MN l=2.2e-07 w=2.4e-07 $[n18ll]
.ENDS
